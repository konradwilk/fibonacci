VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_fibonacci
  CLASS BLOCK ;
  FOREIGN wrapper_fibonacci ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 296.000 25.670 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.720 300.000 1.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.400 300.000 87.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.560 300.000 95.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.200 300.000 110.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.680 300.000 118.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.320 300.000 133.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.480 300.000 142.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.960 300.000 149.560 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.120 300.000 157.720 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.600 300.000 165.200 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.760 300.000 173.360 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.240 300.000 180.840 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.400 300.000 189.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.880 300.000 196.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.520 300.000 212.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.680 300.000 220.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.160 300.000 227.760 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.320 300.000 235.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.800 300.000 243.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.960 300.000 251.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.080 300.000 274.680 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.240 300.000 282.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.720 300.000 290.320 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.000 300.000 32.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.480 300.000 40.080 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.120 300.000 55.720 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 63.280 300.000 63.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.760 300.000 71.360 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.680 300.000 84.280 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.840 300.000 92.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.480 300.000 108.080 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.960 300.000 115.560 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.120 300.000 123.720 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.400 300.000 155.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.880 300.000 162.480 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.040 300.000 170.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.520 300.000 178.120 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.680 300.000 186.280 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.800 300.000 209.400 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.960 300.000 217.560 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.600 300.000 233.200 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.120 300.000 21.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.720 300.000 256.320 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.880 300.000 264.480 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.360 300.000 271.960 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.520 300.000 280.120 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.160 300.000 295.760 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.280 300.000 29.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.760 300.000 37.360 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.400 300.000 53.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.560 300.000 61.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.040 300.000 68.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.200 300.000 76.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.760 300.000 3.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.960 300.000 81.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.120 300.000 89.720 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.600 300.000 97.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.760 300.000 105.360 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.240 300.000 112.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.400 300.000 121.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.520 300.000 144.120 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.680 300.000 152.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.160 300.000 159.760 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.320 300.000 167.920 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.800 300.000 175.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.960 300.000 183.560 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.440 300.000 191.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.600 300.000 199.200 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 206.080 300.000 206.680 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.240 300.000 214.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.880 300.000 230.480 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.400 300.000 19.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.360 300.000 237.960 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.520 300.000 246.120 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.800 300.000 277.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.280 300.000 284.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.440 300.000 293.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.560 300.000 27.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.680 300.000 50.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.840 300.000 58.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.320 300.000 65.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 296.000 297.990 300.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.880 300.000 298.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.960 4.000 251.560 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END la_oenb[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 296.000 2.210 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 296.000 21.530 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 296.000 45.450 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 296.000 85.010 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 296.000 88.690 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 296.000 92.830 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 296.000 96.510 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 296.000 100.650 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 296.000 104.790 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 296.000 108.470 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 296.000 112.610 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 296.000 116.290 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 296.000 120.430 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 296.000 49.130 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 296.000 124.110 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 296.000 128.250 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 296.000 132.390 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 296.000 136.070 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 296.000 140.210 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 296.000 143.890 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 296.000 148.030 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 296.000 152.170 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 296.000 155.850 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 296.000 159.990 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 296.000 53.270 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 296.000 163.670 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 296.000 167.810 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 296.000 57.410 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 296.000 61.090 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 296.000 65.230 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 296.000 68.910 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 296.000 73.050 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 296.000 77.190 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 296.000 80.870 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 296.000 13.710 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 296.000 171.490 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 296.000 211.050 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 296.000 215.190 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 296.000 218.870 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 296.000 223.010 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 296.000 227.150 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 296.000 230.830 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 296.000 234.970 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 296.000 238.650 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 296.000 242.790 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 296.000 246.470 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 296.000 175.630 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 296.000 250.610 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 296.000 254.750 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 296.000 258.430 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 296.000 262.570 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 296.000 266.250 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 296.000 270.390 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 296.000 274.070 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 296.000 278.210 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 296.000 282.350 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 296.000 286.030 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 296.000 179.770 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 296.000 290.170 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 296.000 293.850 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 296.000 183.450 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 296.000 187.590 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 296.000 191.270 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 296.000 195.410 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 296.000 199.090 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 296.000 203.230 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 296.000 207.370 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 4.000 135.960 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 296.000 29.810 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 296.000 33.490 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 296.000 37.630 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 296.000 41.310 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 296.000 10.030 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 296.000 17.850 300.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 288.320 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 288.320 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 288.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 288.320 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 288.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 288.320 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 288.320 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 288.320 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 288.320 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 288.320 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 1.910 0.720 298.010 289.640 ;
      LAYER met2 ;
        RECT 2.490 295.720 5.330 298.365 ;
        RECT 6.170 295.720 9.470 298.365 ;
        RECT 10.310 295.720 13.150 298.365 ;
        RECT 13.990 295.720 17.290 298.365 ;
        RECT 18.130 295.720 20.970 298.365 ;
        RECT 21.810 295.720 25.110 298.365 ;
        RECT 25.950 295.720 29.250 298.365 ;
        RECT 30.090 295.720 32.930 298.365 ;
        RECT 33.770 295.720 37.070 298.365 ;
        RECT 37.910 295.720 40.750 298.365 ;
        RECT 41.590 295.720 44.890 298.365 ;
        RECT 45.730 295.720 48.570 298.365 ;
        RECT 49.410 295.720 52.710 298.365 ;
        RECT 53.550 295.720 56.850 298.365 ;
        RECT 57.690 295.720 60.530 298.365 ;
        RECT 61.370 295.720 64.670 298.365 ;
        RECT 65.510 295.720 68.350 298.365 ;
        RECT 69.190 295.720 72.490 298.365 ;
        RECT 73.330 295.720 76.630 298.365 ;
        RECT 77.470 295.720 80.310 298.365 ;
        RECT 81.150 295.720 84.450 298.365 ;
        RECT 85.290 295.720 88.130 298.365 ;
        RECT 88.970 295.720 92.270 298.365 ;
        RECT 93.110 295.720 95.950 298.365 ;
        RECT 96.790 295.720 100.090 298.365 ;
        RECT 100.930 295.720 104.230 298.365 ;
        RECT 105.070 295.720 107.910 298.365 ;
        RECT 108.750 295.720 112.050 298.365 ;
        RECT 112.890 295.720 115.730 298.365 ;
        RECT 116.570 295.720 119.870 298.365 ;
        RECT 120.710 295.720 123.550 298.365 ;
        RECT 124.390 295.720 127.690 298.365 ;
        RECT 128.530 295.720 131.830 298.365 ;
        RECT 132.670 295.720 135.510 298.365 ;
        RECT 136.350 295.720 139.650 298.365 ;
        RECT 140.490 295.720 143.330 298.365 ;
        RECT 144.170 295.720 147.470 298.365 ;
        RECT 148.310 295.720 151.610 298.365 ;
        RECT 152.450 295.720 155.290 298.365 ;
        RECT 156.130 295.720 159.430 298.365 ;
        RECT 160.270 295.720 163.110 298.365 ;
        RECT 163.950 295.720 167.250 298.365 ;
        RECT 168.090 295.720 170.930 298.365 ;
        RECT 171.770 295.720 175.070 298.365 ;
        RECT 175.910 295.720 179.210 298.365 ;
        RECT 180.050 295.720 182.890 298.365 ;
        RECT 183.730 295.720 187.030 298.365 ;
        RECT 187.870 295.720 190.710 298.365 ;
        RECT 191.550 295.720 194.850 298.365 ;
        RECT 195.690 295.720 198.530 298.365 ;
        RECT 199.370 295.720 202.670 298.365 ;
        RECT 203.510 295.720 206.810 298.365 ;
        RECT 207.650 295.720 210.490 298.365 ;
        RECT 211.330 295.720 214.630 298.365 ;
        RECT 215.470 295.720 218.310 298.365 ;
        RECT 219.150 295.720 222.450 298.365 ;
        RECT 223.290 295.720 226.590 298.365 ;
        RECT 227.430 295.720 230.270 298.365 ;
        RECT 231.110 295.720 234.410 298.365 ;
        RECT 235.250 295.720 238.090 298.365 ;
        RECT 238.930 295.720 242.230 298.365 ;
        RECT 243.070 295.720 245.910 298.365 ;
        RECT 246.750 295.720 250.050 298.365 ;
        RECT 250.890 295.720 254.190 298.365 ;
        RECT 255.030 295.720 257.870 298.365 ;
        RECT 258.710 295.720 262.010 298.365 ;
        RECT 262.850 295.720 265.690 298.365 ;
        RECT 266.530 295.720 269.830 298.365 ;
        RECT 270.670 295.720 273.510 298.365 ;
        RECT 274.350 295.720 277.650 298.365 ;
        RECT 278.490 295.720 281.790 298.365 ;
        RECT 282.630 295.720 285.470 298.365 ;
        RECT 286.310 295.720 289.610 298.365 ;
        RECT 290.450 295.720 293.290 298.365 ;
        RECT 294.130 295.720 297.430 298.365 ;
        RECT 1.940 4.280 297.980 295.720 ;
        RECT 1.940 0.690 2.110 4.280 ;
        RECT 2.950 0.690 6.710 4.280 ;
        RECT 7.550 0.690 11.310 4.280 ;
        RECT 12.150 0.690 15.910 4.280 ;
        RECT 16.750 0.690 20.510 4.280 ;
        RECT 21.350 0.690 25.110 4.280 ;
        RECT 25.950 0.690 30.170 4.280 ;
        RECT 31.010 0.690 34.770 4.280 ;
        RECT 35.610 0.690 39.370 4.280 ;
        RECT 40.210 0.690 43.970 4.280 ;
        RECT 44.810 0.690 48.570 4.280 ;
        RECT 49.410 0.690 53.630 4.280 ;
        RECT 54.470 0.690 58.230 4.280 ;
        RECT 59.070 0.690 62.830 4.280 ;
        RECT 63.670 0.690 67.430 4.280 ;
        RECT 68.270 0.690 72.030 4.280 ;
        RECT 72.870 0.690 77.090 4.280 ;
        RECT 77.930 0.690 81.690 4.280 ;
        RECT 82.530 0.690 86.290 4.280 ;
        RECT 87.130 0.690 90.890 4.280 ;
        RECT 91.730 0.690 95.490 4.280 ;
        RECT 96.330 0.690 100.090 4.280 ;
        RECT 100.930 0.690 105.150 4.280 ;
        RECT 105.990 0.690 109.750 4.280 ;
        RECT 110.590 0.690 114.350 4.280 ;
        RECT 115.190 0.690 118.950 4.280 ;
        RECT 119.790 0.690 123.550 4.280 ;
        RECT 124.390 0.690 128.610 4.280 ;
        RECT 129.450 0.690 133.210 4.280 ;
        RECT 134.050 0.690 137.810 4.280 ;
        RECT 138.650 0.690 142.410 4.280 ;
        RECT 143.250 0.690 147.010 4.280 ;
        RECT 147.850 0.690 152.070 4.280 ;
        RECT 152.910 0.690 156.670 4.280 ;
        RECT 157.510 0.690 161.270 4.280 ;
        RECT 162.110 0.690 165.870 4.280 ;
        RECT 166.710 0.690 170.470 4.280 ;
        RECT 171.310 0.690 175.070 4.280 ;
        RECT 175.910 0.690 180.130 4.280 ;
        RECT 180.970 0.690 184.730 4.280 ;
        RECT 185.570 0.690 189.330 4.280 ;
        RECT 190.170 0.690 193.930 4.280 ;
        RECT 194.770 0.690 198.530 4.280 ;
        RECT 199.370 0.690 203.590 4.280 ;
        RECT 204.430 0.690 208.190 4.280 ;
        RECT 209.030 0.690 212.790 4.280 ;
        RECT 213.630 0.690 217.390 4.280 ;
        RECT 218.230 0.690 221.990 4.280 ;
        RECT 222.830 0.690 227.050 4.280 ;
        RECT 227.890 0.690 231.650 4.280 ;
        RECT 232.490 0.690 236.250 4.280 ;
        RECT 237.090 0.690 240.850 4.280 ;
        RECT 241.690 0.690 245.450 4.280 ;
        RECT 246.290 0.690 250.050 4.280 ;
        RECT 250.890 0.690 255.110 4.280 ;
        RECT 255.950 0.690 259.710 4.280 ;
        RECT 260.550 0.690 264.310 4.280 ;
        RECT 265.150 0.690 268.910 4.280 ;
        RECT 269.750 0.690 273.510 4.280 ;
        RECT 274.350 0.690 278.570 4.280 ;
        RECT 279.410 0.690 283.170 4.280 ;
        RECT 284.010 0.690 287.770 4.280 ;
        RECT 288.610 0.690 292.370 4.280 ;
        RECT 293.210 0.690 296.970 4.280 ;
        RECT 297.810 0.690 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.000 298.200 295.600 298.345 ;
        RECT 4.400 297.480 295.600 298.200 ;
        RECT 4.400 296.800 296.000 297.480 ;
        RECT 4.000 296.160 296.000 296.800 ;
        RECT 4.000 294.760 295.600 296.160 ;
        RECT 4.000 293.440 296.000 294.760 ;
        RECT 4.400 292.040 295.600 293.440 ;
        RECT 4.000 290.720 296.000 292.040 ;
        RECT 4.000 289.320 295.600 290.720 ;
        RECT 4.000 288.680 296.000 289.320 ;
        RECT 4.400 288.000 296.000 288.680 ;
        RECT 4.400 287.280 295.600 288.000 ;
        RECT 4.000 286.600 295.600 287.280 ;
        RECT 4.000 285.280 296.000 286.600 ;
        RECT 4.000 283.920 295.600 285.280 ;
        RECT 4.400 283.880 295.600 283.920 ;
        RECT 4.400 283.240 296.000 283.880 ;
        RECT 4.400 282.520 295.600 283.240 ;
        RECT 4.000 281.840 295.600 282.520 ;
        RECT 4.000 280.520 296.000 281.840 ;
        RECT 4.000 279.840 295.600 280.520 ;
        RECT 4.400 279.120 295.600 279.840 ;
        RECT 4.400 278.440 296.000 279.120 ;
        RECT 4.000 277.800 296.000 278.440 ;
        RECT 4.000 276.400 295.600 277.800 ;
        RECT 4.000 275.080 296.000 276.400 ;
        RECT 4.400 273.680 295.600 275.080 ;
        RECT 4.000 272.360 296.000 273.680 ;
        RECT 4.000 270.960 295.600 272.360 ;
        RECT 4.000 270.320 296.000 270.960 ;
        RECT 4.400 269.640 296.000 270.320 ;
        RECT 4.400 268.920 295.600 269.640 ;
        RECT 4.000 268.240 295.600 268.920 ;
        RECT 4.000 267.600 296.000 268.240 ;
        RECT 4.000 266.200 295.600 267.600 ;
        RECT 4.000 265.560 296.000 266.200 ;
        RECT 4.400 264.880 296.000 265.560 ;
        RECT 4.400 264.160 295.600 264.880 ;
        RECT 4.000 263.480 295.600 264.160 ;
        RECT 4.000 262.160 296.000 263.480 ;
        RECT 4.000 260.800 295.600 262.160 ;
        RECT 4.400 260.760 295.600 260.800 ;
        RECT 4.400 259.440 296.000 260.760 ;
        RECT 4.400 259.400 295.600 259.440 ;
        RECT 4.000 258.040 295.600 259.400 ;
        RECT 4.000 256.720 296.000 258.040 ;
        RECT 4.400 255.320 295.600 256.720 ;
        RECT 4.000 254.000 296.000 255.320 ;
        RECT 4.000 252.600 295.600 254.000 ;
        RECT 4.000 251.960 296.000 252.600 ;
        RECT 4.400 250.560 295.600 251.960 ;
        RECT 4.000 249.240 296.000 250.560 ;
        RECT 4.000 247.840 295.600 249.240 ;
        RECT 4.000 247.200 296.000 247.840 ;
        RECT 4.400 246.520 296.000 247.200 ;
        RECT 4.400 245.800 295.600 246.520 ;
        RECT 4.000 245.120 295.600 245.800 ;
        RECT 4.000 243.800 296.000 245.120 ;
        RECT 4.000 242.440 295.600 243.800 ;
        RECT 4.400 242.400 295.600 242.440 ;
        RECT 4.400 241.080 296.000 242.400 ;
        RECT 4.400 241.040 295.600 241.080 ;
        RECT 4.000 239.680 295.600 241.040 ;
        RECT 4.000 238.360 296.000 239.680 ;
        RECT 4.400 236.960 295.600 238.360 ;
        RECT 4.000 236.320 296.000 236.960 ;
        RECT 4.000 234.920 295.600 236.320 ;
        RECT 4.000 233.600 296.000 234.920 ;
        RECT 4.400 232.200 295.600 233.600 ;
        RECT 4.000 230.880 296.000 232.200 ;
        RECT 4.000 229.480 295.600 230.880 ;
        RECT 4.000 228.840 296.000 229.480 ;
        RECT 4.400 228.160 296.000 228.840 ;
        RECT 4.400 227.440 295.600 228.160 ;
        RECT 4.000 226.760 295.600 227.440 ;
        RECT 4.000 225.440 296.000 226.760 ;
        RECT 4.000 224.080 295.600 225.440 ;
        RECT 4.400 224.040 295.600 224.080 ;
        RECT 4.400 222.720 296.000 224.040 ;
        RECT 4.400 222.680 295.600 222.720 ;
        RECT 4.000 221.320 295.600 222.680 ;
        RECT 4.000 220.680 296.000 221.320 ;
        RECT 4.000 219.320 295.600 220.680 ;
        RECT 4.400 219.280 295.600 219.320 ;
        RECT 4.400 217.960 296.000 219.280 ;
        RECT 4.400 217.920 295.600 217.960 ;
        RECT 4.000 216.560 295.600 217.920 ;
        RECT 4.000 215.240 296.000 216.560 ;
        RECT 4.400 213.840 295.600 215.240 ;
        RECT 4.000 212.520 296.000 213.840 ;
        RECT 4.000 211.120 295.600 212.520 ;
        RECT 4.000 210.480 296.000 211.120 ;
        RECT 4.400 209.800 296.000 210.480 ;
        RECT 4.400 209.080 295.600 209.800 ;
        RECT 4.000 208.400 295.600 209.080 ;
        RECT 4.000 207.080 296.000 208.400 ;
        RECT 4.000 205.720 295.600 207.080 ;
        RECT 4.400 205.680 295.600 205.720 ;
        RECT 4.400 205.040 296.000 205.680 ;
        RECT 4.400 204.320 295.600 205.040 ;
        RECT 4.000 203.640 295.600 204.320 ;
        RECT 4.000 202.320 296.000 203.640 ;
        RECT 4.000 200.960 295.600 202.320 ;
        RECT 4.400 200.920 295.600 200.960 ;
        RECT 4.400 199.600 296.000 200.920 ;
        RECT 4.400 199.560 295.600 199.600 ;
        RECT 4.000 198.200 295.600 199.560 ;
        RECT 4.000 196.880 296.000 198.200 ;
        RECT 4.000 196.200 295.600 196.880 ;
        RECT 4.400 195.480 295.600 196.200 ;
        RECT 4.400 194.800 296.000 195.480 ;
        RECT 4.000 194.160 296.000 194.800 ;
        RECT 4.000 192.760 295.600 194.160 ;
        RECT 4.000 192.120 296.000 192.760 ;
        RECT 4.400 191.440 296.000 192.120 ;
        RECT 4.400 190.720 295.600 191.440 ;
        RECT 4.000 190.040 295.600 190.720 ;
        RECT 4.000 189.400 296.000 190.040 ;
        RECT 4.000 188.000 295.600 189.400 ;
        RECT 4.000 187.360 296.000 188.000 ;
        RECT 4.400 186.680 296.000 187.360 ;
        RECT 4.400 185.960 295.600 186.680 ;
        RECT 4.000 185.280 295.600 185.960 ;
        RECT 4.000 183.960 296.000 185.280 ;
        RECT 4.000 182.600 295.600 183.960 ;
        RECT 4.400 182.560 295.600 182.600 ;
        RECT 4.400 181.240 296.000 182.560 ;
        RECT 4.400 181.200 295.600 181.240 ;
        RECT 4.000 179.840 295.600 181.200 ;
        RECT 4.000 178.520 296.000 179.840 ;
        RECT 4.000 177.840 295.600 178.520 ;
        RECT 4.400 177.120 295.600 177.840 ;
        RECT 4.400 176.440 296.000 177.120 ;
        RECT 4.000 175.800 296.000 176.440 ;
        RECT 4.000 174.400 295.600 175.800 ;
        RECT 4.000 173.760 296.000 174.400 ;
        RECT 4.400 172.360 295.600 173.760 ;
        RECT 4.000 171.040 296.000 172.360 ;
        RECT 4.000 169.640 295.600 171.040 ;
        RECT 4.000 169.000 296.000 169.640 ;
        RECT 4.400 168.320 296.000 169.000 ;
        RECT 4.400 167.600 295.600 168.320 ;
        RECT 4.000 166.920 295.600 167.600 ;
        RECT 4.000 165.600 296.000 166.920 ;
        RECT 4.000 164.240 295.600 165.600 ;
        RECT 4.400 164.200 295.600 164.240 ;
        RECT 4.400 162.880 296.000 164.200 ;
        RECT 4.400 162.840 295.600 162.880 ;
        RECT 4.000 161.480 295.600 162.840 ;
        RECT 4.000 160.160 296.000 161.480 ;
        RECT 4.000 159.480 295.600 160.160 ;
        RECT 4.400 158.760 295.600 159.480 ;
        RECT 4.400 158.120 296.000 158.760 ;
        RECT 4.400 158.080 295.600 158.120 ;
        RECT 4.000 156.720 295.600 158.080 ;
        RECT 4.000 155.400 296.000 156.720 ;
        RECT 4.000 154.720 295.600 155.400 ;
        RECT 4.400 154.000 295.600 154.720 ;
        RECT 4.400 153.320 296.000 154.000 ;
        RECT 4.000 152.680 296.000 153.320 ;
        RECT 4.000 151.280 295.600 152.680 ;
        RECT 4.000 150.640 296.000 151.280 ;
        RECT 4.400 149.960 296.000 150.640 ;
        RECT 4.400 149.240 295.600 149.960 ;
        RECT 4.000 148.560 295.600 149.240 ;
        RECT 4.000 147.240 296.000 148.560 ;
        RECT 4.000 145.880 295.600 147.240 ;
        RECT 4.400 145.840 295.600 145.880 ;
        RECT 4.400 144.520 296.000 145.840 ;
        RECT 4.400 144.480 295.600 144.520 ;
        RECT 4.000 143.120 295.600 144.480 ;
        RECT 4.000 142.480 296.000 143.120 ;
        RECT 4.000 141.120 295.600 142.480 ;
        RECT 4.400 141.080 295.600 141.120 ;
        RECT 4.400 139.760 296.000 141.080 ;
        RECT 4.400 139.720 295.600 139.760 ;
        RECT 4.000 138.360 295.600 139.720 ;
        RECT 4.000 137.040 296.000 138.360 ;
        RECT 4.000 136.360 295.600 137.040 ;
        RECT 4.400 135.640 295.600 136.360 ;
        RECT 4.400 134.960 296.000 135.640 ;
        RECT 4.000 134.320 296.000 134.960 ;
        RECT 4.000 132.920 295.600 134.320 ;
        RECT 4.000 131.600 296.000 132.920 ;
        RECT 4.400 130.200 295.600 131.600 ;
        RECT 4.000 128.880 296.000 130.200 ;
        RECT 4.000 127.520 295.600 128.880 ;
        RECT 4.400 127.480 295.600 127.520 ;
        RECT 4.400 126.840 296.000 127.480 ;
        RECT 4.400 126.120 295.600 126.840 ;
        RECT 4.000 125.440 295.600 126.120 ;
        RECT 4.000 124.120 296.000 125.440 ;
        RECT 4.000 122.760 295.600 124.120 ;
        RECT 4.400 122.720 295.600 122.760 ;
        RECT 4.400 121.400 296.000 122.720 ;
        RECT 4.400 121.360 295.600 121.400 ;
        RECT 4.000 120.000 295.600 121.360 ;
        RECT 4.000 118.680 296.000 120.000 ;
        RECT 4.000 118.000 295.600 118.680 ;
        RECT 4.400 117.280 295.600 118.000 ;
        RECT 4.400 116.600 296.000 117.280 ;
        RECT 4.000 115.960 296.000 116.600 ;
        RECT 4.000 114.560 295.600 115.960 ;
        RECT 4.000 113.240 296.000 114.560 ;
        RECT 4.400 111.840 295.600 113.240 ;
        RECT 4.000 111.200 296.000 111.840 ;
        RECT 4.000 109.800 295.600 111.200 ;
        RECT 4.000 109.160 296.000 109.800 ;
        RECT 4.400 108.480 296.000 109.160 ;
        RECT 4.400 107.760 295.600 108.480 ;
        RECT 4.000 107.080 295.600 107.760 ;
        RECT 4.000 105.760 296.000 107.080 ;
        RECT 4.000 104.400 295.600 105.760 ;
        RECT 4.400 104.360 295.600 104.400 ;
        RECT 4.400 103.040 296.000 104.360 ;
        RECT 4.400 103.000 295.600 103.040 ;
        RECT 4.000 101.640 295.600 103.000 ;
        RECT 4.000 100.320 296.000 101.640 ;
        RECT 4.000 99.640 295.600 100.320 ;
        RECT 4.400 98.920 295.600 99.640 ;
        RECT 4.400 98.240 296.000 98.920 ;
        RECT 4.000 97.600 296.000 98.240 ;
        RECT 4.000 96.200 295.600 97.600 ;
        RECT 4.000 95.560 296.000 96.200 ;
        RECT 4.000 94.880 295.600 95.560 ;
        RECT 4.400 94.160 295.600 94.880 ;
        RECT 4.400 93.480 296.000 94.160 ;
        RECT 4.000 92.840 296.000 93.480 ;
        RECT 4.000 91.440 295.600 92.840 ;
        RECT 4.000 90.120 296.000 91.440 ;
        RECT 4.400 88.720 295.600 90.120 ;
        RECT 4.000 87.400 296.000 88.720 ;
        RECT 4.000 86.040 295.600 87.400 ;
        RECT 4.400 86.000 295.600 86.040 ;
        RECT 4.400 84.680 296.000 86.000 ;
        RECT 4.400 84.640 295.600 84.680 ;
        RECT 4.000 83.280 295.600 84.640 ;
        RECT 4.000 81.960 296.000 83.280 ;
        RECT 4.000 81.280 295.600 81.960 ;
        RECT 4.400 80.560 295.600 81.280 ;
        RECT 4.400 79.920 296.000 80.560 ;
        RECT 4.400 79.880 295.600 79.920 ;
        RECT 4.000 78.520 295.600 79.880 ;
        RECT 4.000 77.200 296.000 78.520 ;
        RECT 4.000 76.520 295.600 77.200 ;
        RECT 4.400 75.800 295.600 76.520 ;
        RECT 4.400 75.120 296.000 75.800 ;
        RECT 4.000 74.480 296.000 75.120 ;
        RECT 4.000 73.080 295.600 74.480 ;
        RECT 4.000 71.760 296.000 73.080 ;
        RECT 4.400 70.360 295.600 71.760 ;
        RECT 4.000 69.040 296.000 70.360 ;
        RECT 4.000 67.640 295.600 69.040 ;
        RECT 4.000 67.000 296.000 67.640 ;
        RECT 4.400 66.320 296.000 67.000 ;
        RECT 4.400 65.600 295.600 66.320 ;
        RECT 4.000 64.920 295.600 65.600 ;
        RECT 4.000 64.280 296.000 64.920 ;
        RECT 4.000 62.920 295.600 64.280 ;
        RECT 4.400 62.880 295.600 62.920 ;
        RECT 4.400 61.560 296.000 62.880 ;
        RECT 4.400 61.520 295.600 61.560 ;
        RECT 4.000 60.160 295.600 61.520 ;
        RECT 4.000 58.840 296.000 60.160 ;
        RECT 4.000 58.160 295.600 58.840 ;
        RECT 4.400 57.440 295.600 58.160 ;
        RECT 4.400 56.760 296.000 57.440 ;
        RECT 4.000 56.120 296.000 56.760 ;
        RECT 4.000 54.720 295.600 56.120 ;
        RECT 4.000 53.400 296.000 54.720 ;
        RECT 4.400 52.000 295.600 53.400 ;
        RECT 4.000 50.680 296.000 52.000 ;
        RECT 4.000 49.280 295.600 50.680 ;
        RECT 4.000 48.640 296.000 49.280 ;
        RECT 4.400 47.240 295.600 48.640 ;
        RECT 4.000 45.920 296.000 47.240 ;
        RECT 4.000 44.560 295.600 45.920 ;
        RECT 4.400 44.520 295.600 44.560 ;
        RECT 4.400 43.200 296.000 44.520 ;
        RECT 4.400 43.160 295.600 43.200 ;
        RECT 4.000 41.800 295.600 43.160 ;
        RECT 4.000 40.480 296.000 41.800 ;
        RECT 4.000 39.800 295.600 40.480 ;
        RECT 4.400 39.080 295.600 39.800 ;
        RECT 4.400 38.400 296.000 39.080 ;
        RECT 4.000 37.760 296.000 38.400 ;
        RECT 4.000 36.360 295.600 37.760 ;
        RECT 4.000 35.040 296.000 36.360 ;
        RECT 4.400 33.640 295.600 35.040 ;
        RECT 4.000 33.000 296.000 33.640 ;
        RECT 4.000 31.600 295.600 33.000 ;
        RECT 4.000 30.280 296.000 31.600 ;
        RECT 4.400 28.880 295.600 30.280 ;
        RECT 4.000 27.560 296.000 28.880 ;
        RECT 4.000 26.160 295.600 27.560 ;
        RECT 4.000 25.520 296.000 26.160 ;
        RECT 4.400 24.840 296.000 25.520 ;
        RECT 4.400 24.120 295.600 24.840 ;
        RECT 4.000 23.440 295.600 24.120 ;
        RECT 4.000 22.120 296.000 23.440 ;
        RECT 4.000 21.440 295.600 22.120 ;
        RECT 4.400 20.720 295.600 21.440 ;
        RECT 4.400 20.040 296.000 20.720 ;
        RECT 4.000 19.400 296.000 20.040 ;
        RECT 4.000 18.000 295.600 19.400 ;
        RECT 4.000 17.360 296.000 18.000 ;
        RECT 4.000 16.680 295.600 17.360 ;
        RECT 4.400 15.960 295.600 16.680 ;
        RECT 4.400 15.280 296.000 15.960 ;
        RECT 4.000 14.640 296.000 15.280 ;
        RECT 4.000 13.240 295.600 14.640 ;
        RECT 4.000 11.920 296.000 13.240 ;
        RECT 4.400 10.520 295.600 11.920 ;
        RECT 4.000 9.200 296.000 10.520 ;
        RECT 4.000 7.800 295.600 9.200 ;
        RECT 4.000 7.160 296.000 7.800 ;
        RECT 4.400 6.480 296.000 7.160 ;
        RECT 4.400 5.760 295.600 6.480 ;
        RECT 4.000 5.080 295.600 5.760 ;
        RECT 4.000 3.760 296.000 5.080 ;
        RECT 4.000 3.080 295.600 3.760 ;
        RECT 4.400 2.360 295.600 3.080 ;
        RECT 4.400 1.720 296.000 2.360 ;
        RECT 4.400 1.680 295.600 1.720 ;
        RECT 4.000 0.855 295.600 1.680 ;
      LAYER met4 ;
        RECT 221.095 95.375 251.040 269.785 ;
        RECT 253.440 95.375 254.340 269.785 ;
        RECT 256.740 95.375 257.640 269.785 ;
        RECT 260.040 95.375 260.940 269.785 ;
        RECT 263.340 95.375 288.585 269.785 ;
  END
END wrapper_fibonacci
END LIBRARY

