VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_fibonacci
  CLASS BLOCK ;
  FOREIGN wrapper_fibonacci ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 346.000 29.490 350.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1.100 350.000 2.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 92.220 350.000 93.420 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 101.060 350.000 102.260 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 110.580 350.000 111.780 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 119.420 350.000 120.620 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 128.940 350.000 130.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 137.780 350.000 138.980 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 146.620 350.000 147.820 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 156.140 350.000 157.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 164.980 350.000 166.180 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 174.500 350.000 175.700 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 9.940 350.000 11.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 183.340 350.000 184.540 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 192.860 350.000 194.060 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 201.700 350.000 202.900 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 211.220 350.000 212.420 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 220.060 350.000 221.260 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 228.900 350.000 230.100 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 238.420 350.000 239.620 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 247.260 350.000 248.460 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 256.780 350.000 257.980 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.620 350.000 266.820 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 18.780 350.000 19.980 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 275.140 350.000 276.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 283.980 350.000 285.180 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 292.820 350.000 294.020 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 302.340 350.000 303.540 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.180 350.000 312.380 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 320.700 350.000 321.900 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.540 350.000 330.740 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 339.060 350.000 340.260 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 28.300 350.000 29.500 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 37.140 350.000 38.340 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 46.660 350.000 47.860 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 55.500 350.000 56.700 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 65.020 350.000 66.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 73.860 350.000 75.060 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 82.700 350.000 83.900 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 6.540 350.000 7.740 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 98.340 350.000 99.540 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 107.180 350.000 108.380 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 116.700 350.000 117.900 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 125.540 350.000 126.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 135.060 350.000 136.260 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 143.900 350.000 145.100 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 152.740 350.000 153.940 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 162.260 350.000 163.460 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 171.100 350.000 172.300 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 180.620 350.000 181.820 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 16.060 350.000 17.260 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 189.460 350.000 190.660 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 198.980 350.000 200.180 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 207.820 350.000 209.020 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.660 350.000 217.860 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 226.180 350.000 227.380 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 235.020 350.000 236.220 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 244.540 350.000 245.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 253.380 350.000 254.580 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 262.900 350.000 264.100 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 271.740 350.000 272.940 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 24.900 350.000 26.100 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 281.260 350.000 282.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 290.100 350.000 291.300 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 298.940 350.000 300.140 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 308.460 350.000 309.660 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.300 350.000 318.500 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 326.820 350.000 328.020 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.660 350.000 336.860 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 345.180 350.000 346.380 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.420 350.000 35.620 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 43.260 350.000 44.460 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 52.780 350.000 53.980 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 61.620 350.000 62.820 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 71.140 350.000 72.340 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 79.980 350.000 81.180 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 88.820 350.000 90.020 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 3.820 350.000 5.020 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 94.940 350.000 96.140 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 104.460 350.000 105.660 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 113.300 350.000 114.500 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 122.820 350.000 124.020 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 131.660 350.000 132.860 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 141.180 350.000 142.380 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 150.020 350.000 151.220 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 158.860 350.000 160.060 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 168.380 350.000 169.580 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 177.220 350.000 178.420 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 12.660 350.000 13.860 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 186.740 350.000 187.940 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 195.580 350.000 196.780 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 205.100 350.000 206.300 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 213.940 350.000 215.140 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 222.780 350.000 223.980 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 232.300 350.000 233.500 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 241.140 350.000 242.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 250.660 350.000 251.860 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 259.500 350.000 260.700 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 269.020 350.000 270.220 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 22.180 350.000 23.380 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 277.860 350.000 279.060 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 286.700 350.000 287.900 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 296.220 350.000 297.420 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 305.060 350.000 306.260 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.580 350.000 315.780 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.420 350.000 324.620 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 332.940 350.000 334.140 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 341.780 350.000 342.980 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 31.020 350.000 32.220 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.540 350.000 41.740 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 49.380 350.000 50.580 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 58.900 350.000 60.100 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 67.740 350.000 68.940 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 76.580 350.000 77.780 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 86.100 350.000 87.300 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 0.000 347.350 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 346.000 347.810 350.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 347.900 350.000 349.100 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 0.000 2.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 0.000 56.630 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 0.000 61.690 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.650 0.000 67.210 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.170 0.000 72.730 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.230 0.000 77.790 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 0.000 83.310 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.270 0.000 88.830 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.790 0.000 94.350 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 0.000 99.410 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 0.000 104.930 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.310 0.000 7.870 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 0.000 110.450 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 0.000 115.510 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 0.000 121.030 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 0.000 126.550 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.050 0.000 131.610 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.570 0.000 137.130 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.090 0.000 142.650 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.610 0.000 148.170 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.670 0.000 153.230 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.190 0.000 158.750 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.710 0.000 164.270 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.770 0.000 169.330 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.410 0.000 23.970 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.930 0.000 29.490 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.450 0.000 35.010 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 0.000 40.070 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.030 0.000 45.590 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 0.000 51.110 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.290 0.000 174.850 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 0.000 228.670 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.630 0.000 234.190 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 0.000 239.710 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.210 0.000 244.770 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.730 0.000 250.290 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 0.000 255.810 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.310 0.000 260.870 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.830 0.000 266.390 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.350 0.000 271.910 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.870 0.000 277.430 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 0.000 180.370 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.930 0.000 282.490 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.450 0.000 288.010 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.970 0.000 293.530 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 0.000 298.590 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.550 0.000 304.110 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 0.000 309.630 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.590 0.000 315.150 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 0.000 320.210 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.170 0.000 325.730 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.690 0.000 331.250 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.330 0.000 185.890 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 0.000 336.310 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 0.000 341.830 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.390 0.000 190.950 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.910 0.000 196.470 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 0.000 201.990 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.490 0.000 207.050 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.010 0.000 212.570 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.530 0.000 218.090 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.050 0.000 223.610 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.220 4.000 178.420 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.620 4.000 232.820 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.740 4.000 238.940 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.180 4.000 244.380 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.620 4.000 249.820 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.060 4.000 255.260 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.500 4.000 260.700 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.940 4.000 266.140 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.380 4.000 271.580 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.820 4.000 277.020 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.260 4.000 282.460 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.660 4.000 183.860 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.700 4.000 287.900 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.140 4.000 293.340 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.580 4.000 298.780 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.020 4.000 304.220 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.460 4.000 309.660 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.900 4.000 315.100 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.340 4.000 320.540 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.780 4.000 325.980 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.220 4.000 331.420 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.660 4.000 336.860 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.100 4.000 189.300 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.100 4.000 342.300 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.540 4.000 347.740 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.540 4.000 194.740 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.980 4.000 200.180 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.420 4.000 205.620 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.860 4.000 211.060 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.300 4.000 216.500 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.180 4.000 227.380 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.530 346.000 34.090 350.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 346.000 2.350 350.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.930 346.000 6.490 350.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.330 346.000 24.890 350.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.070 346.000 56.630 350.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.610 346.000 102.170 350.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.210 346.000 106.770 350.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.810 346.000 111.370 350.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 346.000 115.970 350.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.550 346.000 120.110 350.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.150 346.000 124.710 350.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 346.000 129.310 350.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 346.000 133.910 350.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.950 346.000 138.510 350.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 346.000 143.110 350.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.670 346.000 61.230 350.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.150 346.000 147.710 350.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.750 346.000 152.310 350.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 346.000 156.910 350.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.490 346.000 161.050 350.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.090 346.000 165.650 350.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.690 346.000 170.250 350.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.290 346.000 174.850 350.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.890 346.000 179.450 350.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.490 346.000 184.050 350.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.090 346.000 188.650 350.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.270 346.000 65.830 350.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 346.000 193.250 350.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.830 346.000 197.390 350.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.870 346.000 70.430 350.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.470 346.000 75.030 350.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 346.000 79.630 350.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.210 346.000 83.770 350.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.810 346.000 88.370 350.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.410 346.000 92.970 350.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 346.000 97.570 350.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.130 346.000 15.690 350.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.430 346.000 201.990 350.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.970 346.000 247.530 350.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.570 346.000 252.130 350.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.170 346.000 256.730 350.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.770 346.000 261.330 350.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.370 346.000 265.930 350.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 346.000 270.530 350.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.110 346.000 274.670 350.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.710 346.000 279.270 350.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 346.000 283.870 350.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.910 346.000 288.470 350.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 346.000 206.590 350.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.510 346.000 293.070 350.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 346.000 297.670 350.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.710 346.000 302.270 350.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.310 346.000 306.870 350.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.910 346.000 311.470 350.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.050 346.000 315.610 350.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 346.000 320.210 350.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.250 346.000 324.810 350.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.850 346.000 329.410 350.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 346.000 334.010 350.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.630 346.000 211.190 350.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.050 346.000 338.610 350.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.650 346.000 343.210 350.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 346.000 215.790 350.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 346.000 220.390 350.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.430 346.000 224.990 350.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.030 346.000 229.590 350.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.630 346.000 234.190 350.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.770 346.000 238.330 350.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 346.000 242.930 350.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.460 4.000 3.660 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.860 4.000 58.060 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.300 4.000 63.500 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.180 4.000 74.380 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.620 4.000 79.820 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.060 4.000 85.260 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.500 4.000 90.700 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.380 4.000 101.580 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.820 4.000 107.020 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.900 4.000 9.100 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.260 4.000 112.460 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.820 4.000 124.020 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.260 4.000 129.460 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.700 4.000 134.900 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.140 4.000 140.340 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.580 4.000 145.780 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.020 4.000 151.220 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.460 4.000 156.660 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.900 4.000 162.100 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.340 4.000 167.540 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.780 4.000 172.980 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.780 4.000 19.980 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.220 4.000 25.420 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.660 4.000 30.860 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.100 4.000 36.300 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.980 4.000 47.180 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.420 4.000 52.620 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 346.000 38.690 350.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.270 346.000 42.830 350.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 346.000 47.430 350.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 346.000 52.030 350.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.530 346.000 11.090 350.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.730 346.000 20.290 350.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 349.915 343.655 ;
      LAYER met1 ;
        RECT 0.070 10.640 349.975 345.740 ;
      LAYER met2 ;
        RECT 0.100 345.720 1.510 348.685 ;
        RECT 2.630 345.720 5.650 348.685 ;
        RECT 6.770 345.720 10.250 348.685 ;
        RECT 11.370 345.720 14.850 348.685 ;
        RECT 15.970 345.720 19.450 348.685 ;
        RECT 20.570 345.720 24.050 348.685 ;
        RECT 25.170 345.720 28.650 348.685 ;
        RECT 29.770 345.720 33.250 348.685 ;
        RECT 34.370 345.720 37.850 348.685 ;
        RECT 38.970 345.720 41.990 348.685 ;
        RECT 43.110 345.720 46.590 348.685 ;
        RECT 47.710 345.720 51.190 348.685 ;
        RECT 52.310 345.720 55.790 348.685 ;
        RECT 56.910 345.720 60.390 348.685 ;
        RECT 61.510 345.720 64.990 348.685 ;
        RECT 66.110 345.720 69.590 348.685 ;
        RECT 70.710 345.720 74.190 348.685 ;
        RECT 75.310 345.720 78.790 348.685 ;
        RECT 79.910 345.720 82.930 348.685 ;
        RECT 84.050 345.720 87.530 348.685 ;
        RECT 88.650 345.720 92.130 348.685 ;
        RECT 93.250 345.720 96.730 348.685 ;
        RECT 97.850 345.720 101.330 348.685 ;
        RECT 102.450 345.720 105.930 348.685 ;
        RECT 107.050 345.720 110.530 348.685 ;
        RECT 111.650 345.720 115.130 348.685 ;
        RECT 116.250 345.720 119.270 348.685 ;
        RECT 120.390 345.720 123.870 348.685 ;
        RECT 124.990 345.720 128.470 348.685 ;
        RECT 129.590 345.720 133.070 348.685 ;
        RECT 134.190 345.720 137.670 348.685 ;
        RECT 138.790 345.720 142.270 348.685 ;
        RECT 143.390 345.720 146.870 348.685 ;
        RECT 147.990 345.720 151.470 348.685 ;
        RECT 152.590 345.720 156.070 348.685 ;
        RECT 157.190 345.720 160.210 348.685 ;
        RECT 161.330 345.720 164.810 348.685 ;
        RECT 165.930 345.720 169.410 348.685 ;
        RECT 170.530 345.720 174.010 348.685 ;
        RECT 175.130 345.720 178.610 348.685 ;
        RECT 179.730 345.720 183.210 348.685 ;
        RECT 184.330 345.720 187.810 348.685 ;
        RECT 188.930 345.720 192.410 348.685 ;
        RECT 193.530 345.720 196.550 348.685 ;
        RECT 197.670 345.720 201.150 348.685 ;
        RECT 202.270 345.720 205.750 348.685 ;
        RECT 206.870 345.720 210.350 348.685 ;
        RECT 211.470 345.720 214.950 348.685 ;
        RECT 216.070 345.720 219.550 348.685 ;
        RECT 220.670 345.720 224.150 348.685 ;
        RECT 225.270 345.720 228.750 348.685 ;
        RECT 229.870 345.720 233.350 348.685 ;
        RECT 234.470 345.720 237.490 348.685 ;
        RECT 238.610 345.720 242.090 348.685 ;
        RECT 243.210 345.720 246.690 348.685 ;
        RECT 247.810 345.720 251.290 348.685 ;
        RECT 252.410 345.720 255.890 348.685 ;
        RECT 257.010 345.720 260.490 348.685 ;
        RECT 261.610 345.720 265.090 348.685 ;
        RECT 266.210 345.720 269.690 348.685 ;
        RECT 270.810 345.720 273.830 348.685 ;
        RECT 274.950 345.720 278.430 348.685 ;
        RECT 279.550 345.720 283.030 348.685 ;
        RECT 284.150 345.720 287.630 348.685 ;
        RECT 288.750 345.720 292.230 348.685 ;
        RECT 293.350 345.720 296.830 348.685 ;
        RECT 297.950 345.720 301.430 348.685 ;
        RECT 302.550 345.720 306.030 348.685 ;
        RECT 307.150 345.720 310.630 348.685 ;
        RECT 311.750 345.720 314.770 348.685 ;
        RECT 315.890 345.720 319.370 348.685 ;
        RECT 320.490 345.720 323.970 348.685 ;
        RECT 325.090 345.720 328.570 348.685 ;
        RECT 329.690 345.720 333.170 348.685 ;
        RECT 334.290 345.720 337.770 348.685 ;
        RECT 338.890 345.720 342.370 348.685 ;
        RECT 343.490 345.720 346.970 348.685 ;
        RECT 348.090 345.720 348.590 348.685 ;
        RECT 0.100 4.280 348.590 345.720 ;
        RECT 0.100 2.875 1.970 4.280 ;
        RECT 3.090 2.875 7.030 4.280 ;
        RECT 8.150 2.875 12.550 4.280 ;
        RECT 13.670 2.875 18.070 4.280 ;
        RECT 19.190 2.875 23.130 4.280 ;
        RECT 24.250 2.875 28.650 4.280 ;
        RECT 29.770 2.875 34.170 4.280 ;
        RECT 35.290 2.875 39.230 4.280 ;
        RECT 40.350 2.875 44.750 4.280 ;
        RECT 45.870 2.875 50.270 4.280 ;
        RECT 51.390 2.875 55.790 4.280 ;
        RECT 56.910 2.875 60.850 4.280 ;
        RECT 61.970 2.875 66.370 4.280 ;
        RECT 67.490 2.875 71.890 4.280 ;
        RECT 73.010 2.875 76.950 4.280 ;
        RECT 78.070 2.875 82.470 4.280 ;
        RECT 83.590 2.875 87.990 4.280 ;
        RECT 89.110 2.875 93.510 4.280 ;
        RECT 94.630 2.875 98.570 4.280 ;
        RECT 99.690 2.875 104.090 4.280 ;
        RECT 105.210 2.875 109.610 4.280 ;
        RECT 110.730 2.875 114.670 4.280 ;
        RECT 115.790 2.875 120.190 4.280 ;
        RECT 121.310 2.875 125.710 4.280 ;
        RECT 126.830 2.875 130.770 4.280 ;
        RECT 131.890 2.875 136.290 4.280 ;
        RECT 137.410 2.875 141.810 4.280 ;
        RECT 142.930 2.875 147.330 4.280 ;
        RECT 148.450 2.875 152.390 4.280 ;
        RECT 153.510 2.875 157.910 4.280 ;
        RECT 159.030 2.875 163.430 4.280 ;
        RECT 164.550 2.875 168.490 4.280 ;
        RECT 169.610 2.875 174.010 4.280 ;
        RECT 175.130 2.875 179.530 4.280 ;
        RECT 180.650 2.875 185.050 4.280 ;
        RECT 186.170 2.875 190.110 4.280 ;
        RECT 191.230 2.875 195.630 4.280 ;
        RECT 196.750 2.875 201.150 4.280 ;
        RECT 202.270 2.875 206.210 4.280 ;
        RECT 207.330 2.875 211.730 4.280 ;
        RECT 212.850 2.875 217.250 4.280 ;
        RECT 218.370 2.875 222.770 4.280 ;
        RECT 223.890 2.875 227.830 4.280 ;
        RECT 228.950 2.875 233.350 4.280 ;
        RECT 234.470 2.875 238.870 4.280 ;
        RECT 239.990 2.875 243.930 4.280 ;
        RECT 245.050 2.875 249.450 4.280 ;
        RECT 250.570 2.875 254.970 4.280 ;
        RECT 256.090 2.875 260.030 4.280 ;
        RECT 261.150 2.875 265.550 4.280 ;
        RECT 266.670 2.875 271.070 4.280 ;
        RECT 272.190 2.875 276.590 4.280 ;
        RECT 277.710 2.875 281.650 4.280 ;
        RECT 282.770 2.875 287.170 4.280 ;
        RECT 288.290 2.875 292.690 4.280 ;
        RECT 293.810 2.875 297.750 4.280 ;
        RECT 298.870 2.875 303.270 4.280 ;
        RECT 304.390 2.875 308.790 4.280 ;
        RECT 309.910 2.875 314.310 4.280 ;
        RECT 315.430 2.875 319.370 4.280 ;
        RECT 320.490 2.875 324.890 4.280 ;
        RECT 326.010 2.875 330.410 4.280 ;
        RECT 331.530 2.875 335.470 4.280 ;
        RECT 336.590 2.875 340.990 4.280 ;
        RECT 342.110 2.875 346.510 4.280 ;
        RECT 347.630 2.875 348.590 4.280 ;
      LAYER met3 ;
        RECT 4.000 348.140 345.600 348.665 ;
        RECT 4.400 347.500 345.600 348.140 ;
        RECT 4.400 346.780 348.615 347.500 ;
        RECT 4.400 346.140 345.600 346.780 ;
        RECT 4.000 344.780 345.600 346.140 ;
        RECT 4.000 343.380 348.615 344.780 ;
        RECT 4.000 342.700 345.600 343.380 ;
        RECT 4.400 341.380 345.600 342.700 ;
        RECT 4.400 340.700 348.615 341.380 ;
        RECT 4.000 340.660 348.615 340.700 ;
        RECT 4.000 338.660 345.600 340.660 ;
        RECT 4.000 337.260 348.615 338.660 ;
        RECT 4.400 335.260 345.600 337.260 ;
        RECT 4.000 334.540 348.615 335.260 ;
        RECT 4.000 332.540 345.600 334.540 ;
        RECT 4.000 331.820 348.615 332.540 ;
        RECT 4.400 331.140 348.615 331.820 ;
        RECT 4.400 329.820 345.600 331.140 ;
        RECT 4.000 329.140 345.600 329.820 ;
        RECT 4.000 328.420 348.615 329.140 ;
        RECT 4.000 326.420 345.600 328.420 ;
        RECT 4.000 326.380 348.615 326.420 ;
        RECT 4.400 325.020 348.615 326.380 ;
        RECT 4.400 324.380 345.600 325.020 ;
        RECT 4.000 323.020 345.600 324.380 ;
        RECT 4.000 322.300 348.615 323.020 ;
        RECT 4.000 320.940 345.600 322.300 ;
        RECT 4.400 320.300 345.600 320.940 ;
        RECT 4.400 318.940 348.615 320.300 ;
        RECT 4.000 318.900 348.615 318.940 ;
        RECT 4.000 316.900 345.600 318.900 ;
        RECT 4.000 316.180 348.615 316.900 ;
        RECT 4.000 315.500 345.600 316.180 ;
        RECT 4.400 314.180 345.600 315.500 ;
        RECT 4.400 313.500 348.615 314.180 ;
        RECT 4.000 312.780 348.615 313.500 ;
        RECT 4.000 310.780 345.600 312.780 ;
        RECT 4.000 310.060 348.615 310.780 ;
        RECT 4.400 308.060 345.600 310.060 ;
        RECT 4.000 306.660 348.615 308.060 ;
        RECT 4.000 304.660 345.600 306.660 ;
        RECT 4.000 304.620 348.615 304.660 ;
        RECT 4.400 303.940 348.615 304.620 ;
        RECT 4.400 302.620 345.600 303.940 ;
        RECT 4.000 301.940 345.600 302.620 ;
        RECT 4.000 300.540 348.615 301.940 ;
        RECT 4.000 299.180 345.600 300.540 ;
        RECT 4.400 298.540 345.600 299.180 ;
        RECT 4.400 297.820 348.615 298.540 ;
        RECT 4.400 297.180 345.600 297.820 ;
        RECT 4.000 295.820 345.600 297.180 ;
        RECT 4.000 294.420 348.615 295.820 ;
        RECT 4.000 293.740 345.600 294.420 ;
        RECT 4.400 292.420 345.600 293.740 ;
        RECT 4.400 291.740 348.615 292.420 ;
        RECT 4.000 291.700 348.615 291.740 ;
        RECT 4.000 289.700 345.600 291.700 ;
        RECT 4.000 288.300 348.615 289.700 ;
        RECT 4.400 286.300 345.600 288.300 ;
        RECT 4.000 285.580 348.615 286.300 ;
        RECT 4.000 283.580 345.600 285.580 ;
        RECT 4.000 282.860 348.615 283.580 ;
        RECT 4.400 280.860 345.600 282.860 ;
        RECT 4.000 279.460 348.615 280.860 ;
        RECT 4.000 277.460 345.600 279.460 ;
        RECT 4.000 277.420 348.615 277.460 ;
        RECT 4.400 276.740 348.615 277.420 ;
        RECT 4.400 275.420 345.600 276.740 ;
        RECT 4.000 274.740 345.600 275.420 ;
        RECT 4.000 273.340 348.615 274.740 ;
        RECT 4.000 271.980 345.600 273.340 ;
        RECT 4.400 271.340 345.600 271.980 ;
        RECT 4.400 270.620 348.615 271.340 ;
        RECT 4.400 269.980 345.600 270.620 ;
        RECT 4.000 268.620 345.600 269.980 ;
        RECT 4.000 267.220 348.615 268.620 ;
        RECT 4.000 266.540 345.600 267.220 ;
        RECT 4.400 265.220 345.600 266.540 ;
        RECT 4.400 264.540 348.615 265.220 ;
        RECT 4.000 264.500 348.615 264.540 ;
        RECT 4.000 262.500 345.600 264.500 ;
        RECT 4.000 261.100 348.615 262.500 ;
        RECT 4.400 259.100 345.600 261.100 ;
        RECT 4.000 258.380 348.615 259.100 ;
        RECT 4.000 256.380 345.600 258.380 ;
        RECT 4.000 255.660 348.615 256.380 ;
        RECT 4.400 254.980 348.615 255.660 ;
        RECT 4.400 253.660 345.600 254.980 ;
        RECT 4.000 252.980 345.600 253.660 ;
        RECT 4.000 252.260 348.615 252.980 ;
        RECT 4.000 250.260 345.600 252.260 ;
        RECT 4.000 250.220 348.615 250.260 ;
        RECT 4.400 248.860 348.615 250.220 ;
        RECT 4.400 248.220 345.600 248.860 ;
        RECT 4.000 246.860 345.600 248.220 ;
        RECT 4.000 246.140 348.615 246.860 ;
        RECT 4.000 244.780 345.600 246.140 ;
        RECT 4.400 244.140 345.600 244.780 ;
        RECT 4.400 242.780 348.615 244.140 ;
        RECT 4.000 242.740 348.615 242.780 ;
        RECT 4.000 240.740 345.600 242.740 ;
        RECT 4.000 240.020 348.615 240.740 ;
        RECT 4.000 239.340 345.600 240.020 ;
        RECT 4.400 238.020 345.600 239.340 ;
        RECT 4.400 237.340 348.615 238.020 ;
        RECT 4.000 236.620 348.615 237.340 ;
        RECT 4.000 234.620 345.600 236.620 ;
        RECT 4.000 233.900 348.615 234.620 ;
        RECT 4.000 233.220 345.600 233.900 ;
        RECT 4.400 231.900 345.600 233.220 ;
        RECT 4.400 231.220 348.615 231.900 ;
        RECT 4.000 230.500 348.615 231.220 ;
        RECT 4.000 228.500 345.600 230.500 ;
        RECT 4.000 227.780 348.615 228.500 ;
        RECT 4.400 225.780 345.600 227.780 ;
        RECT 4.000 224.380 348.615 225.780 ;
        RECT 4.000 222.380 345.600 224.380 ;
        RECT 4.000 222.340 348.615 222.380 ;
        RECT 4.400 221.660 348.615 222.340 ;
        RECT 4.400 220.340 345.600 221.660 ;
        RECT 4.000 219.660 345.600 220.340 ;
        RECT 4.000 218.260 348.615 219.660 ;
        RECT 4.000 216.900 345.600 218.260 ;
        RECT 4.400 216.260 345.600 216.900 ;
        RECT 4.400 215.540 348.615 216.260 ;
        RECT 4.400 214.900 345.600 215.540 ;
        RECT 4.000 213.540 345.600 214.900 ;
        RECT 4.000 212.820 348.615 213.540 ;
        RECT 4.000 211.460 345.600 212.820 ;
        RECT 4.400 210.820 345.600 211.460 ;
        RECT 4.400 209.460 348.615 210.820 ;
        RECT 4.000 209.420 348.615 209.460 ;
        RECT 4.000 207.420 345.600 209.420 ;
        RECT 4.000 206.700 348.615 207.420 ;
        RECT 4.000 206.020 345.600 206.700 ;
        RECT 4.400 204.700 345.600 206.020 ;
        RECT 4.400 204.020 348.615 204.700 ;
        RECT 4.000 203.300 348.615 204.020 ;
        RECT 4.000 201.300 345.600 203.300 ;
        RECT 4.000 200.580 348.615 201.300 ;
        RECT 4.400 198.580 345.600 200.580 ;
        RECT 4.000 197.180 348.615 198.580 ;
        RECT 4.000 195.180 345.600 197.180 ;
        RECT 4.000 195.140 348.615 195.180 ;
        RECT 4.400 194.460 348.615 195.140 ;
        RECT 4.400 193.140 345.600 194.460 ;
        RECT 4.000 192.460 345.600 193.140 ;
        RECT 4.000 191.060 348.615 192.460 ;
        RECT 4.000 189.700 345.600 191.060 ;
        RECT 4.400 189.060 345.600 189.700 ;
        RECT 4.400 188.340 348.615 189.060 ;
        RECT 4.400 187.700 345.600 188.340 ;
        RECT 4.000 186.340 345.600 187.700 ;
        RECT 4.000 184.940 348.615 186.340 ;
        RECT 4.000 184.260 345.600 184.940 ;
        RECT 4.400 182.940 345.600 184.260 ;
        RECT 4.400 182.260 348.615 182.940 ;
        RECT 4.000 182.220 348.615 182.260 ;
        RECT 4.000 180.220 345.600 182.220 ;
        RECT 4.000 178.820 348.615 180.220 ;
        RECT 4.400 176.820 345.600 178.820 ;
        RECT 4.000 176.100 348.615 176.820 ;
        RECT 4.000 174.100 345.600 176.100 ;
        RECT 4.000 173.380 348.615 174.100 ;
        RECT 4.400 172.700 348.615 173.380 ;
        RECT 4.400 171.380 345.600 172.700 ;
        RECT 4.000 170.700 345.600 171.380 ;
        RECT 4.000 169.980 348.615 170.700 ;
        RECT 4.000 167.980 345.600 169.980 ;
        RECT 4.000 167.940 348.615 167.980 ;
        RECT 4.400 166.580 348.615 167.940 ;
        RECT 4.400 165.940 345.600 166.580 ;
        RECT 4.000 164.580 345.600 165.940 ;
        RECT 4.000 163.860 348.615 164.580 ;
        RECT 4.000 162.500 345.600 163.860 ;
        RECT 4.400 161.860 345.600 162.500 ;
        RECT 4.400 160.500 348.615 161.860 ;
        RECT 4.000 160.460 348.615 160.500 ;
        RECT 4.000 158.460 345.600 160.460 ;
        RECT 4.000 157.740 348.615 158.460 ;
        RECT 4.000 157.060 345.600 157.740 ;
        RECT 4.400 155.740 345.600 157.060 ;
        RECT 4.400 155.060 348.615 155.740 ;
        RECT 4.000 154.340 348.615 155.060 ;
        RECT 4.000 152.340 345.600 154.340 ;
        RECT 4.000 151.620 348.615 152.340 ;
        RECT 4.400 149.620 345.600 151.620 ;
        RECT 4.000 148.220 348.615 149.620 ;
        RECT 4.000 146.220 345.600 148.220 ;
        RECT 4.000 146.180 348.615 146.220 ;
        RECT 4.400 145.500 348.615 146.180 ;
        RECT 4.400 144.180 345.600 145.500 ;
        RECT 4.000 143.500 345.600 144.180 ;
        RECT 4.000 142.780 348.615 143.500 ;
        RECT 4.000 140.780 345.600 142.780 ;
        RECT 4.000 140.740 348.615 140.780 ;
        RECT 4.400 139.380 348.615 140.740 ;
        RECT 4.400 138.740 345.600 139.380 ;
        RECT 4.000 137.380 345.600 138.740 ;
        RECT 4.000 136.660 348.615 137.380 ;
        RECT 4.000 135.300 345.600 136.660 ;
        RECT 4.400 134.660 345.600 135.300 ;
        RECT 4.400 133.300 348.615 134.660 ;
        RECT 4.000 133.260 348.615 133.300 ;
        RECT 4.000 131.260 345.600 133.260 ;
        RECT 4.000 130.540 348.615 131.260 ;
        RECT 4.000 129.860 345.600 130.540 ;
        RECT 4.400 128.540 345.600 129.860 ;
        RECT 4.400 127.860 348.615 128.540 ;
        RECT 4.000 127.140 348.615 127.860 ;
        RECT 4.000 125.140 345.600 127.140 ;
        RECT 4.000 124.420 348.615 125.140 ;
        RECT 4.400 122.420 345.600 124.420 ;
        RECT 4.000 121.020 348.615 122.420 ;
        RECT 4.000 119.020 345.600 121.020 ;
        RECT 4.000 118.300 348.615 119.020 ;
        RECT 4.400 116.300 345.600 118.300 ;
        RECT 4.000 114.900 348.615 116.300 ;
        RECT 4.000 112.900 345.600 114.900 ;
        RECT 4.000 112.860 348.615 112.900 ;
        RECT 4.400 112.180 348.615 112.860 ;
        RECT 4.400 110.860 345.600 112.180 ;
        RECT 4.000 110.180 345.600 110.860 ;
        RECT 4.000 108.780 348.615 110.180 ;
        RECT 4.000 107.420 345.600 108.780 ;
        RECT 4.400 106.780 345.600 107.420 ;
        RECT 4.400 106.060 348.615 106.780 ;
        RECT 4.400 105.420 345.600 106.060 ;
        RECT 4.000 104.060 345.600 105.420 ;
        RECT 4.000 102.660 348.615 104.060 ;
        RECT 4.000 101.980 345.600 102.660 ;
        RECT 4.400 100.660 345.600 101.980 ;
        RECT 4.400 99.980 348.615 100.660 ;
        RECT 4.000 99.940 348.615 99.980 ;
        RECT 4.000 97.940 345.600 99.940 ;
        RECT 4.000 96.540 348.615 97.940 ;
        RECT 4.400 94.540 345.600 96.540 ;
        RECT 4.000 93.820 348.615 94.540 ;
        RECT 4.000 91.820 345.600 93.820 ;
        RECT 4.000 91.100 348.615 91.820 ;
        RECT 4.400 90.420 348.615 91.100 ;
        RECT 4.400 89.100 345.600 90.420 ;
        RECT 4.000 88.420 345.600 89.100 ;
        RECT 4.000 87.700 348.615 88.420 ;
        RECT 4.000 85.700 345.600 87.700 ;
        RECT 4.000 85.660 348.615 85.700 ;
        RECT 4.400 84.300 348.615 85.660 ;
        RECT 4.400 83.660 345.600 84.300 ;
        RECT 4.000 82.300 345.600 83.660 ;
        RECT 4.000 81.580 348.615 82.300 ;
        RECT 4.000 80.220 345.600 81.580 ;
        RECT 4.400 79.580 345.600 80.220 ;
        RECT 4.400 78.220 348.615 79.580 ;
        RECT 4.000 78.180 348.615 78.220 ;
        RECT 4.000 76.180 345.600 78.180 ;
        RECT 4.000 75.460 348.615 76.180 ;
        RECT 4.000 74.780 345.600 75.460 ;
        RECT 4.400 73.460 345.600 74.780 ;
        RECT 4.400 72.780 348.615 73.460 ;
        RECT 4.000 72.740 348.615 72.780 ;
        RECT 4.000 70.740 345.600 72.740 ;
        RECT 4.000 69.340 348.615 70.740 ;
        RECT 4.400 67.340 345.600 69.340 ;
        RECT 4.000 66.620 348.615 67.340 ;
        RECT 4.000 64.620 345.600 66.620 ;
        RECT 4.000 63.900 348.615 64.620 ;
        RECT 4.400 63.220 348.615 63.900 ;
        RECT 4.400 61.900 345.600 63.220 ;
        RECT 4.000 61.220 345.600 61.900 ;
        RECT 4.000 60.500 348.615 61.220 ;
        RECT 4.000 58.500 345.600 60.500 ;
        RECT 4.000 58.460 348.615 58.500 ;
        RECT 4.400 57.100 348.615 58.460 ;
        RECT 4.400 56.460 345.600 57.100 ;
        RECT 4.000 55.100 345.600 56.460 ;
        RECT 4.000 54.380 348.615 55.100 ;
        RECT 4.000 53.020 345.600 54.380 ;
        RECT 4.400 52.380 345.600 53.020 ;
        RECT 4.400 51.020 348.615 52.380 ;
        RECT 4.000 50.980 348.615 51.020 ;
        RECT 4.000 48.980 345.600 50.980 ;
        RECT 4.000 48.260 348.615 48.980 ;
        RECT 4.000 47.580 345.600 48.260 ;
        RECT 4.400 46.260 345.600 47.580 ;
        RECT 4.400 45.580 348.615 46.260 ;
        RECT 4.000 44.860 348.615 45.580 ;
        RECT 4.000 42.860 345.600 44.860 ;
        RECT 4.000 42.140 348.615 42.860 ;
        RECT 4.400 40.140 345.600 42.140 ;
        RECT 4.000 38.740 348.615 40.140 ;
        RECT 4.000 36.740 345.600 38.740 ;
        RECT 4.000 36.700 348.615 36.740 ;
        RECT 4.400 36.020 348.615 36.700 ;
        RECT 4.400 34.700 345.600 36.020 ;
        RECT 4.000 34.020 345.600 34.700 ;
        RECT 4.000 32.620 348.615 34.020 ;
        RECT 4.000 31.260 345.600 32.620 ;
        RECT 4.400 30.620 345.600 31.260 ;
        RECT 4.400 29.900 348.615 30.620 ;
        RECT 4.400 29.260 345.600 29.900 ;
        RECT 4.000 27.900 345.600 29.260 ;
        RECT 4.000 26.500 348.615 27.900 ;
        RECT 4.000 25.820 345.600 26.500 ;
        RECT 4.400 24.500 345.600 25.820 ;
        RECT 4.400 23.820 348.615 24.500 ;
        RECT 4.000 23.780 348.615 23.820 ;
        RECT 4.000 21.780 345.600 23.780 ;
        RECT 4.000 20.380 348.615 21.780 ;
        RECT 4.400 18.380 345.600 20.380 ;
        RECT 4.000 17.660 348.615 18.380 ;
        RECT 4.000 15.660 345.600 17.660 ;
        RECT 4.000 14.940 348.615 15.660 ;
        RECT 4.400 14.260 348.615 14.940 ;
        RECT 4.400 12.940 345.600 14.260 ;
        RECT 4.000 12.260 345.600 12.940 ;
        RECT 4.000 11.540 348.615 12.260 ;
        RECT 4.000 9.540 345.600 11.540 ;
        RECT 4.000 9.500 348.615 9.540 ;
        RECT 4.400 8.140 348.615 9.500 ;
        RECT 4.400 7.500 345.600 8.140 ;
        RECT 4.000 6.140 345.600 7.500 ;
        RECT 4.000 5.420 348.615 6.140 ;
        RECT 4.000 4.060 345.600 5.420 ;
        RECT 4.400 3.420 345.600 4.060 ;
        RECT 4.400 2.895 348.615 3.420 ;
      LAYER met4 ;
        RECT 53.655 337.920 337.345 340.505 ;
        RECT 53.655 95.375 97.440 337.920 ;
        RECT 99.840 95.375 174.240 337.920 ;
        RECT 176.640 95.375 251.040 337.920 ;
        RECT 253.440 95.375 327.840 337.920 ;
        RECT 330.240 95.375 337.345 337.920 ;
  END
END wrapper_fibonacci
END LIBRARY

