VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapper_fibonacci
  CLASS BLOCK ;
  FOREIGN wrapper_fibonacci ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 296.000 25.210 300.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 0.720 300.000 1.320 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 78.920 300.000 79.520 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 86.400 300.000 87.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 94.560 300.000 95.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 102.040 300.000 102.640 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 110.200 300.000 110.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 117.680 300.000 118.280 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 125.840 300.000 126.440 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 133.320 300.000 133.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 141.480 300.000 142.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 148.960 300.000 149.560 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 8.200 300.000 8.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 157.120 300.000 157.720 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 164.600 300.000 165.200 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 172.760 300.000 173.360 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 180.240 300.000 180.840 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 188.400 300.000 189.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 195.880 300.000 196.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 204.040 300.000 204.640 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 211.520 300.000 212.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 219.680 300.000 220.280 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 227.160 300.000 227.760 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 16.360 300.000 16.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 235.320 300.000 235.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 242.800 300.000 243.400 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 250.960 300.000 251.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 258.440 300.000 259.040 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 266.600 300.000 267.200 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 274.080 300.000 274.680 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 282.240 300.000 282.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 289.720 300.000 290.320 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 32.000 300.000 32.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 39.480 300.000 40.080 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 55.120 300.000 55.720 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 63.280 300.000 63.880 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 70.760 300.000 71.360 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 5.480 300.000 6.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 83.680 300.000 84.280 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 91.840 300.000 92.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 99.320 300.000 99.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 107.480 300.000 108.080 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 114.960 300.000 115.560 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 123.120 300.000 123.720 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 130.600 300.000 131.200 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 138.760 300.000 139.360 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 146.240 300.000 146.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 154.400 300.000 155.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 161.880 300.000 162.480 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 170.040 300.000 170.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 177.520 300.000 178.120 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 185.680 300.000 186.280 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 193.160 300.000 193.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 201.320 300.000 201.920 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 208.800 300.000 209.400 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 216.960 300.000 217.560 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 224.440 300.000 225.040 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 232.600 300.000 233.200 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 21.120 300.000 21.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 240.080 300.000 240.680 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 248.240 300.000 248.840 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 255.720 300.000 256.320 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 263.880 300.000 264.480 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 271.360 300.000 271.960 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 279.520 300.000 280.120 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 287.000 300.000 287.600 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 295.160 300.000 295.760 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 29.280 300.000 29.880 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 36.760 300.000 37.360 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 44.920 300.000 45.520 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 52.400 300.000 53.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 60.560 300.000 61.160 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 68.040 300.000 68.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 76.200 300.000 76.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 2.760 300.000 3.360 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 80.960 300.000 81.560 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 89.120 300.000 89.720 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 96.600 300.000 97.200 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 104.760 300.000 105.360 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.240 300.000 112.840 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 120.400 300.000 121.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 127.880 300.000 128.480 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 143.520 300.000 144.120 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 151.680 300.000 152.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.920 300.000 11.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 159.160 300.000 159.760 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 167.320 300.000 167.920 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 174.800 300.000 175.400 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 182.960 300.000 183.560 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 190.440 300.000 191.040 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 198.600 300.000 199.200 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 206.080 300.000 206.680 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 214.240 300.000 214.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 221.720 300.000 222.320 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 229.880 300.000 230.480 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 18.400 300.000 19.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 237.360 300.000 237.960 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 245.520 300.000 246.120 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 253.000 300.000 253.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 261.160 300.000 261.760 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 268.640 300.000 269.240 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 276.800 300.000 277.400 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 284.280 300.000 284.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 292.440 300.000 293.040 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 26.560 300.000 27.160 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 42.200 300.000 42.800 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 49.680 300.000 50.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.840 300.000 58.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 65.320 300.000 65.920 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 73.480 300.000 74.080 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 296.000 294.310 300.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 297.880 300.000 298.480 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 296.000 297.990 300.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.680 4.000 288.280 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 296.000 28.890 300.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 296.000 2.210 300.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 296.000 5.890 300.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 296.000 21.070 300.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 296.000 48.210 300.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 296.000 86.390 300.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 296.000 90.530 300.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 296.000 94.210 300.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 296.000 97.890 300.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 296.000 102.030 300.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 296.000 105.710 300.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 296.000 109.850 300.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 296.000 113.530 300.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 296.000 117.210 300.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 296.000 121.350 300.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 296.000 51.890 300.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 296.000 125.030 300.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 296.000 128.710 300.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 296.000 132.850 300.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 296.000 136.530 300.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 296.000 140.210 300.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 296.000 144.350 300.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 296.000 148.030 300.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 296.000 152.170 300.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 296.000 155.850 300.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 296.000 159.530 300.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 296.000 56.030 300.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 296.000 163.670 300.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 296.000 167.350 300.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 296.000 59.710 300.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 296.000 63.390 300.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 296.000 67.530 300.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 296.000 71.210 300.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 296.000 74.890 300.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 296.000 79.030 300.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 296.000 82.710 300.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 296.000 13.710 300.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 296.000 171.030 300.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 296.000 209.670 300.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 296.000 213.350 300.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 296.000 217.490 300.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 296.000 221.170 300.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 296.000 224.850 300.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 296.000 228.990 300.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 296.000 232.670 300.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 296.000 236.350 300.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 296.000 240.490 300.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 296.000 244.170 300.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 296.000 175.170 300.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 296.000 247.850 300.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 296.000 251.990 300.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 296.000 255.670 300.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 296.000 259.810 300.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 296.000 263.490 300.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 296.000 267.170 300.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 296.000 271.310 300.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 296.000 274.990 300.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 296.000 278.670 300.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 296.000 282.810 300.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 296.000 178.850 300.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 296.000 286.490 300.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 296.000 290.170 300.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 296.000 182.530 300.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 296.000 186.670 300.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 296.000 190.350 300.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 296.000 194.030 300.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 296.000 198.170 300.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 296.000 201.850 300.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 296.000 205.990 300.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 296.000 32.570 300.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 296.000 36.710 300.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 296.000 40.390 300.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 296.000 44.070 300.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 296.000 9.570 300.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 296.000 17.390 300.000 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 288.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 288.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 288.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 288.560 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 288.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 288.320 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 288.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 288.320 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 288.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 288.320 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 288.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 288.320 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 288.320 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 288.320 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 288.320 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 288.320 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 294.400 288.405 ;
      LAYER met1 ;
        RECT 1.910 1.400 298.010 290.320 ;
      LAYER met2 ;
        RECT 2.490 295.720 5.330 298.365 ;
        RECT 6.170 295.720 9.010 298.365 ;
        RECT 9.850 295.720 13.150 298.365 ;
        RECT 13.990 295.720 16.830 298.365 ;
        RECT 17.670 295.720 20.510 298.365 ;
        RECT 21.350 295.720 24.650 298.365 ;
        RECT 25.490 295.720 28.330 298.365 ;
        RECT 29.170 295.720 32.010 298.365 ;
        RECT 32.850 295.720 36.150 298.365 ;
        RECT 36.990 295.720 39.830 298.365 ;
        RECT 40.670 295.720 43.510 298.365 ;
        RECT 44.350 295.720 47.650 298.365 ;
        RECT 48.490 295.720 51.330 298.365 ;
        RECT 52.170 295.720 55.470 298.365 ;
        RECT 56.310 295.720 59.150 298.365 ;
        RECT 59.990 295.720 62.830 298.365 ;
        RECT 63.670 295.720 66.970 298.365 ;
        RECT 67.810 295.720 70.650 298.365 ;
        RECT 71.490 295.720 74.330 298.365 ;
        RECT 75.170 295.720 78.470 298.365 ;
        RECT 79.310 295.720 82.150 298.365 ;
        RECT 82.990 295.720 85.830 298.365 ;
        RECT 86.670 295.720 89.970 298.365 ;
        RECT 90.810 295.720 93.650 298.365 ;
        RECT 94.490 295.720 97.330 298.365 ;
        RECT 98.170 295.720 101.470 298.365 ;
        RECT 102.310 295.720 105.150 298.365 ;
        RECT 105.990 295.720 109.290 298.365 ;
        RECT 110.130 295.720 112.970 298.365 ;
        RECT 113.810 295.720 116.650 298.365 ;
        RECT 117.490 295.720 120.790 298.365 ;
        RECT 121.630 295.720 124.470 298.365 ;
        RECT 125.310 295.720 128.150 298.365 ;
        RECT 128.990 295.720 132.290 298.365 ;
        RECT 133.130 295.720 135.970 298.365 ;
        RECT 136.810 295.720 139.650 298.365 ;
        RECT 140.490 295.720 143.790 298.365 ;
        RECT 144.630 295.720 147.470 298.365 ;
        RECT 148.310 295.720 151.610 298.365 ;
        RECT 152.450 295.720 155.290 298.365 ;
        RECT 156.130 295.720 158.970 298.365 ;
        RECT 159.810 295.720 163.110 298.365 ;
        RECT 163.950 295.720 166.790 298.365 ;
        RECT 167.630 295.720 170.470 298.365 ;
        RECT 171.310 295.720 174.610 298.365 ;
        RECT 175.450 295.720 178.290 298.365 ;
        RECT 179.130 295.720 181.970 298.365 ;
        RECT 182.810 295.720 186.110 298.365 ;
        RECT 186.950 295.720 189.790 298.365 ;
        RECT 190.630 295.720 193.470 298.365 ;
        RECT 194.310 295.720 197.610 298.365 ;
        RECT 198.450 295.720 201.290 298.365 ;
        RECT 202.130 295.720 205.430 298.365 ;
        RECT 206.270 295.720 209.110 298.365 ;
        RECT 209.950 295.720 212.790 298.365 ;
        RECT 213.630 295.720 216.930 298.365 ;
        RECT 217.770 295.720 220.610 298.365 ;
        RECT 221.450 295.720 224.290 298.365 ;
        RECT 225.130 295.720 228.430 298.365 ;
        RECT 229.270 295.720 232.110 298.365 ;
        RECT 232.950 295.720 235.790 298.365 ;
        RECT 236.630 295.720 239.930 298.365 ;
        RECT 240.770 295.720 243.610 298.365 ;
        RECT 244.450 295.720 247.290 298.365 ;
        RECT 248.130 295.720 251.430 298.365 ;
        RECT 252.270 295.720 255.110 298.365 ;
        RECT 255.950 295.720 259.250 298.365 ;
        RECT 260.090 295.720 262.930 298.365 ;
        RECT 263.770 295.720 266.610 298.365 ;
        RECT 267.450 295.720 270.750 298.365 ;
        RECT 271.590 295.720 274.430 298.365 ;
        RECT 275.270 295.720 278.110 298.365 ;
        RECT 278.950 295.720 282.250 298.365 ;
        RECT 283.090 295.720 285.930 298.365 ;
        RECT 286.770 295.720 289.610 298.365 ;
        RECT 290.450 295.720 293.750 298.365 ;
        RECT 294.590 295.720 297.430 298.365 ;
        RECT 1.940 4.280 297.980 295.720 ;
        RECT 1.940 0.835 2.110 4.280 ;
        RECT 2.950 0.835 6.710 4.280 ;
        RECT 7.550 0.835 11.310 4.280 ;
        RECT 12.150 0.835 15.910 4.280 ;
        RECT 16.750 0.835 20.510 4.280 ;
        RECT 21.350 0.835 25.110 4.280 ;
        RECT 25.950 0.835 30.170 4.280 ;
        RECT 31.010 0.835 34.770 4.280 ;
        RECT 35.610 0.835 39.370 4.280 ;
        RECT 40.210 0.835 43.970 4.280 ;
        RECT 44.810 0.835 48.570 4.280 ;
        RECT 49.410 0.835 53.630 4.280 ;
        RECT 54.470 0.835 58.230 4.280 ;
        RECT 59.070 0.835 62.830 4.280 ;
        RECT 63.670 0.835 67.430 4.280 ;
        RECT 68.270 0.835 72.030 4.280 ;
        RECT 72.870 0.835 77.090 4.280 ;
        RECT 77.930 0.835 81.690 4.280 ;
        RECT 82.530 0.835 86.290 4.280 ;
        RECT 87.130 0.835 90.890 4.280 ;
        RECT 91.730 0.835 95.490 4.280 ;
        RECT 96.330 0.835 100.090 4.280 ;
        RECT 100.930 0.835 105.150 4.280 ;
        RECT 105.990 0.835 109.750 4.280 ;
        RECT 110.590 0.835 114.350 4.280 ;
        RECT 115.190 0.835 118.950 4.280 ;
        RECT 119.790 0.835 123.550 4.280 ;
        RECT 124.390 0.835 128.610 4.280 ;
        RECT 129.450 0.835 133.210 4.280 ;
        RECT 134.050 0.835 137.810 4.280 ;
        RECT 138.650 0.835 142.410 4.280 ;
        RECT 143.250 0.835 147.010 4.280 ;
        RECT 147.850 0.835 152.070 4.280 ;
        RECT 152.910 0.835 156.670 4.280 ;
        RECT 157.510 0.835 161.270 4.280 ;
        RECT 162.110 0.835 165.870 4.280 ;
        RECT 166.710 0.835 170.470 4.280 ;
        RECT 171.310 0.835 175.070 4.280 ;
        RECT 175.910 0.835 180.130 4.280 ;
        RECT 180.970 0.835 184.730 4.280 ;
        RECT 185.570 0.835 189.330 4.280 ;
        RECT 190.170 0.835 193.930 4.280 ;
        RECT 194.770 0.835 198.530 4.280 ;
        RECT 199.370 0.835 203.590 4.280 ;
        RECT 204.430 0.835 208.190 4.280 ;
        RECT 209.030 0.835 212.790 4.280 ;
        RECT 213.630 0.835 217.390 4.280 ;
        RECT 218.230 0.835 221.990 4.280 ;
        RECT 222.830 0.835 227.050 4.280 ;
        RECT 227.890 0.835 231.650 4.280 ;
        RECT 232.490 0.835 236.250 4.280 ;
        RECT 237.090 0.835 240.850 4.280 ;
        RECT 241.690 0.835 245.450 4.280 ;
        RECT 246.290 0.835 250.050 4.280 ;
        RECT 250.890 0.835 255.110 4.280 ;
        RECT 255.950 0.835 259.710 4.280 ;
        RECT 260.550 0.835 264.310 4.280 ;
        RECT 265.150 0.835 268.910 4.280 ;
        RECT 269.750 0.835 273.510 4.280 ;
        RECT 274.350 0.835 278.570 4.280 ;
        RECT 279.410 0.835 283.170 4.280 ;
        RECT 284.010 0.835 287.770 4.280 ;
        RECT 288.610 0.835 292.370 4.280 ;
        RECT 293.210 0.835 296.970 4.280 ;
        RECT 297.810 0.835 297.980 4.280 ;
      LAYER met3 ;
        RECT 4.000 298.200 295.600 298.345 ;
        RECT 4.400 297.480 295.600 298.200 ;
        RECT 4.400 296.800 296.000 297.480 ;
        RECT 4.000 296.160 296.000 296.800 ;
        RECT 4.000 294.760 295.600 296.160 ;
        RECT 4.000 293.440 296.000 294.760 ;
        RECT 4.400 292.040 295.600 293.440 ;
        RECT 4.000 290.720 296.000 292.040 ;
        RECT 4.000 289.320 295.600 290.720 ;
        RECT 4.000 288.680 296.000 289.320 ;
        RECT 4.400 288.000 296.000 288.680 ;
        RECT 4.400 287.280 295.600 288.000 ;
        RECT 4.000 286.600 295.600 287.280 ;
        RECT 4.000 285.280 296.000 286.600 ;
        RECT 4.000 283.920 295.600 285.280 ;
        RECT 4.400 283.880 295.600 283.920 ;
        RECT 4.400 283.240 296.000 283.880 ;
        RECT 4.400 282.520 295.600 283.240 ;
        RECT 4.000 281.840 295.600 282.520 ;
        RECT 4.000 280.520 296.000 281.840 ;
        RECT 4.000 279.160 295.600 280.520 ;
        RECT 4.400 279.120 295.600 279.160 ;
        RECT 4.400 277.800 296.000 279.120 ;
        RECT 4.400 277.760 295.600 277.800 ;
        RECT 4.000 276.400 295.600 277.760 ;
        RECT 4.000 275.080 296.000 276.400 ;
        RECT 4.000 274.400 295.600 275.080 ;
        RECT 4.400 273.680 295.600 274.400 ;
        RECT 4.400 273.000 296.000 273.680 ;
        RECT 4.000 272.360 296.000 273.000 ;
        RECT 4.000 270.960 295.600 272.360 ;
        RECT 4.000 269.640 296.000 270.960 ;
        RECT 4.400 268.240 295.600 269.640 ;
        RECT 4.000 267.600 296.000 268.240 ;
        RECT 4.000 266.200 295.600 267.600 ;
        RECT 4.000 264.880 296.000 266.200 ;
        RECT 4.400 263.480 295.600 264.880 ;
        RECT 4.000 262.160 296.000 263.480 ;
        RECT 4.000 260.760 295.600 262.160 ;
        RECT 4.000 260.120 296.000 260.760 ;
        RECT 4.400 259.440 296.000 260.120 ;
        RECT 4.400 258.720 295.600 259.440 ;
        RECT 4.000 258.040 295.600 258.720 ;
        RECT 4.000 256.720 296.000 258.040 ;
        RECT 4.000 256.040 295.600 256.720 ;
        RECT 4.400 255.320 295.600 256.040 ;
        RECT 4.400 254.640 296.000 255.320 ;
        RECT 4.000 254.000 296.000 254.640 ;
        RECT 4.000 252.600 295.600 254.000 ;
        RECT 4.000 251.960 296.000 252.600 ;
        RECT 4.000 251.280 295.600 251.960 ;
        RECT 4.400 250.560 295.600 251.280 ;
        RECT 4.400 249.880 296.000 250.560 ;
        RECT 4.000 249.240 296.000 249.880 ;
        RECT 4.000 247.840 295.600 249.240 ;
        RECT 4.000 246.520 296.000 247.840 ;
        RECT 4.400 245.120 295.600 246.520 ;
        RECT 4.000 243.800 296.000 245.120 ;
        RECT 4.000 242.400 295.600 243.800 ;
        RECT 4.000 241.760 296.000 242.400 ;
        RECT 4.400 241.080 296.000 241.760 ;
        RECT 4.400 240.360 295.600 241.080 ;
        RECT 4.000 239.680 295.600 240.360 ;
        RECT 4.000 238.360 296.000 239.680 ;
        RECT 4.000 237.000 295.600 238.360 ;
        RECT 4.400 236.960 295.600 237.000 ;
        RECT 4.400 236.320 296.000 236.960 ;
        RECT 4.400 235.600 295.600 236.320 ;
        RECT 4.000 234.920 295.600 235.600 ;
        RECT 4.000 233.600 296.000 234.920 ;
        RECT 4.000 232.240 295.600 233.600 ;
        RECT 4.400 232.200 295.600 232.240 ;
        RECT 4.400 230.880 296.000 232.200 ;
        RECT 4.400 230.840 295.600 230.880 ;
        RECT 4.000 229.480 295.600 230.840 ;
        RECT 4.000 228.160 296.000 229.480 ;
        RECT 4.000 227.480 295.600 228.160 ;
        RECT 4.400 226.760 295.600 227.480 ;
        RECT 4.400 226.080 296.000 226.760 ;
        RECT 4.000 225.440 296.000 226.080 ;
        RECT 4.000 224.040 295.600 225.440 ;
        RECT 4.000 222.720 296.000 224.040 ;
        RECT 4.400 221.320 295.600 222.720 ;
        RECT 4.000 220.680 296.000 221.320 ;
        RECT 4.000 219.280 295.600 220.680 ;
        RECT 4.000 217.960 296.000 219.280 ;
        RECT 4.400 216.560 295.600 217.960 ;
        RECT 4.000 215.240 296.000 216.560 ;
        RECT 4.000 213.880 295.600 215.240 ;
        RECT 4.400 213.840 295.600 213.880 ;
        RECT 4.400 212.520 296.000 213.840 ;
        RECT 4.400 212.480 295.600 212.520 ;
        RECT 4.000 211.120 295.600 212.480 ;
        RECT 4.000 209.800 296.000 211.120 ;
        RECT 4.000 209.120 295.600 209.800 ;
        RECT 4.400 208.400 295.600 209.120 ;
        RECT 4.400 207.720 296.000 208.400 ;
        RECT 4.000 207.080 296.000 207.720 ;
        RECT 4.000 205.680 295.600 207.080 ;
        RECT 4.000 205.040 296.000 205.680 ;
        RECT 4.000 204.360 295.600 205.040 ;
        RECT 4.400 203.640 295.600 204.360 ;
        RECT 4.400 202.960 296.000 203.640 ;
        RECT 4.000 202.320 296.000 202.960 ;
        RECT 4.000 200.920 295.600 202.320 ;
        RECT 4.000 199.600 296.000 200.920 ;
        RECT 4.400 198.200 295.600 199.600 ;
        RECT 4.000 196.880 296.000 198.200 ;
        RECT 4.000 195.480 295.600 196.880 ;
        RECT 4.000 194.840 296.000 195.480 ;
        RECT 4.400 194.160 296.000 194.840 ;
        RECT 4.400 193.440 295.600 194.160 ;
        RECT 4.000 192.760 295.600 193.440 ;
        RECT 4.000 191.440 296.000 192.760 ;
        RECT 4.000 190.080 295.600 191.440 ;
        RECT 4.400 190.040 295.600 190.080 ;
        RECT 4.400 189.400 296.000 190.040 ;
        RECT 4.400 188.680 295.600 189.400 ;
        RECT 4.000 188.000 295.600 188.680 ;
        RECT 4.000 186.680 296.000 188.000 ;
        RECT 4.000 185.320 295.600 186.680 ;
        RECT 4.400 185.280 295.600 185.320 ;
        RECT 4.400 183.960 296.000 185.280 ;
        RECT 4.400 183.920 295.600 183.960 ;
        RECT 4.000 182.560 295.600 183.920 ;
        RECT 4.000 181.240 296.000 182.560 ;
        RECT 4.000 180.560 295.600 181.240 ;
        RECT 4.400 179.840 295.600 180.560 ;
        RECT 4.400 179.160 296.000 179.840 ;
        RECT 4.000 178.520 296.000 179.160 ;
        RECT 4.000 177.120 295.600 178.520 ;
        RECT 4.000 175.800 296.000 177.120 ;
        RECT 4.400 174.400 295.600 175.800 ;
        RECT 4.000 173.760 296.000 174.400 ;
        RECT 4.000 172.360 295.600 173.760 ;
        RECT 4.000 171.720 296.000 172.360 ;
        RECT 4.400 171.040 296.000 171.720 ;
        RECT 4.400 170.320 295.600 171.040 ;
        RECT 4.000 169.640 295.600 170.320 ;
        RECT 4.000 168.320 296.000 169.640 ;
        RECT 4.000 166.960 295.600 168.320 ;
        RECT 4.400 166.920 295.600 166.960 ;
        RECT 4.400 165.600 296.000 166.920 ;
        RECT 4.400 165.560 295.600 165.600 ;
        RECT 4.000 164.200 295.600 165.560 ;
        RECT 4.000 162.880 296.000 164.200 ;
        RECT 4.000 162.200 295.600 162.880 ;
        RECT 4.400 161.480 295.600 162.200 ;
        RECT 4.400 160.800 296.000 161.480 ;
        RECT 4.000 160.160 296.000 160.800 ;
        RECT 4.000 158.760 295.600 160.160 ;
        RECT 4.000 158.120 296.000 158.760 ;
        RECT 4.000 157.440 295.600 158.120 ;
        RECT 4.400 156.720 295.600 157.440 ;
        RECT 4.400 156.040 296.000 156.720 ;
        RECT 4.000 155.400 296.000 156.040 ;
        RECT 4.000 154.000 295.600 155.400 ;
        RECT 4.000 152.680 296.000 154.000 ;
        RECT 4.400 151.280 295.600 152.680 ;
        RECT 4.000 149.960 296.000 151.280 ;
        RECT 4.000 148.560 295.600 149.960 ;
        RECT 4.000 147.920 296.000 148.560 ;
        RECT 4.400 147.240 296.000 147.920 ;
        RECT 4.400 146.520 295.600 147.240 ;
        RECT 4.000 145.840 295.600 146.520 ;
        RECT 4.000 144.520 296.000 145.840 ;
        RECT 4.000 143.160 295.600 144.520 ;
        RECT 4.400 143.120 295.600 143.160 ;
        RECT 4.400 142.480 296.000 143.120 ;
        RECT 4.400 141.760 295.600 142.480 ;
        RECT 4.000 141.080 295.600 141.760 ;
        RECT 4.000 139.760 296.000 141.080 ;
        RECT 4.000 138.400 295.600 139.760 ;
        RECT 4.400 138.360 295.600 138.400 ;
        RECT 4.400 137.040 296.000 138.360 ;
        RECT 4.400 137.000 295.600 137.040 ;
        RECT 4.000 135.640 295.600 137.000 ;
        RECT 4.000 134.320 296.000 135.640 ;
        RECT 4.000 133.640 295.600 134.320 ;
        RECT 4.400 132.920 295.600 133.640 ;
        RECT 4.400 132.240 296.000 132.920 ;
        RECT 4.000 131.600 296.000 132.240 ;
        RECT 4.000 130.200 295.600 131.600 ;
        RECT 4.000 129.560 296.000 130.200 ;
        RECT 4.400 128.880 296.000 129.560 ;
        RECT 4.400 128.160 295.600 128.880 ;
        RECT 4.000 127.480 295.600 128.160 ;
        RECT 4.000 126.840 296.000 127.480 ;
        RECT 4.000 125.440 295.600 126.840 ;
        RECT 4.000 124.800 296.000 125.440 ;
        RECT 4.400 124.120 296.000 124.800 ;
        RECT 4.400 123.400 295.600 124.120 ;
        RECT 4.000 122.720 295.600 123.400 ;
        RECT 4.000 121.400 296.000 122.720 ;
        RECT 4.000 120.040 295.600 121.400 ;
        RECT 4.400 120.000 295.600 120.040 ;
        RECT 4.400 118.680 296.000 120.000 ;
        RECT 4.400 118.640 295.600 118.680 ;
        RECT 4.000 117.280 295.600 118.640 ;
        RECT 4.000 115.960 296.000 117.280 ;
        RECT 4.000 115.280 295.600 115.960 ;
        RECT 4.400 114.560 295.600 115.280 ;
        RECT 4.400 113.880 296.000 114.560 ;
        RECT 4.000 113.240 296.000 113.880 ;
        RECT 4.000 111.840 295.600 113.240 ;
        RECT 4.000 111.200 296.000 111.840 ;
        RECT 4.000 110.520 295.600 111.200 ;
        RECT 4.400 109.800 295.600 110.520 ;
        RECT 4.400 109.120 296.000 109.800 ;
        RECT 4.000 108.480 296.000 109.120 ;
        RECT 4.000 107.080 295.600 108.480 ;
        RECT 4.000 105.760 296.000 107.080 ;
        RECT 4.400 104.360 295.600 105.760 ;
        RECT 4.000 103.040 296.000 104.360 ;
        RECT 4.000 101.640 295.600 103.040 ;
        RECT 4.000 101.000 296.000 101.640 ;
        RECT 4.400 100.320 296.000 101.000 ;
        RECT 4.400 99.600 295.600 100.320 ;
        RECT 4.000 98.920 295.600 99.600 ;
        RECT 4.000 97.600 296.000 98.920 ;
        RECT 4.000 96.240 295.600 97.600 ;
        RECT 4.400 96.200 295.600 96.240 ;
        RECT 4.400 95.560 296.000 96.200 ;
        RECT 4.400 94.840 295.600 95.560 ;
        RECT 4.000 94.160 295.600 94.840 ;
        RECT 4.000 92.840 296.000 94.160 ;
        RECT 4.000 91.480 295.600 92.840 ;
        RECT 4.400 91.440 295.600 91.480 ;
        RECT 4.400 90.120 296.000 91.440 ;
        RECT 4.400 90.080 295.600 90.120 ;
        RECT 4.000 88.720 295.600 90.080 ;
        RECT 4.000 87.400 296.000 88.720 ;
        RECT 4.400 86.000 295.600 87.400 ;
        RECT 4.000 84.680 296.000 86.000 ;
        RECT 4.000 83.280 295.600 84.680 ;
        RECT 4.000 82.640 296.000 83.280 ;
        RECT 4.400 81.960 296.000 82.640 ;
        RECT 4.400 81.240 295.600 81.960 ;
        RECT 4.000 80.560 295.600 81.240 ;
        RECT 4.000 79.920 296.000 80.560 ;
        RECT 4.000 78.520 295.600 79.920 ;
        RECT 4.000 77.880 296.000 78.520 ;
        RECT 4.400 77.200 296.000 77.880 ;
        RECT 4.400 76.480 295.600 77.200 ;
        RECT 4.000 75.800 295.600 76.480 ;
        RECT 4.000 74.480 296.000 75.800 ;
        RECT 4.000 73.120 295.600 74.480 ;
        RECT 4.400 73.080 295.600 73.120 ;
        RECT 4.400 71.760 296.000 73.080 ;
        RECT 4.400 71.720 295.600 71.760 ;
        RECT 4.000 70.360 295.600 71.720 ;
        RECT 4.000 69.040 296.000 70.360 ;
        RECT 4.000 68.360 295.600 69.040 ;
        RECT 4.400 67.640 295.600 68.360 ;
        RECT 4.400 66.960 296.000 67.640 ;
        RECT 4.000 66.320 296.000 66.960 ;
        RECT 4.000 64.920 295.600 66.320 ;
        RECT 4.000 64.280 296.000 64.920 ;
        RECT 4.000 63.600 295.600 64.280 ;
        RECT 4.400 62.880 295.600 63.600 ;
        RECT 4.400 62.200 296.000 62.880 ;
        RECT 4.000 61.560 296.000 62.200 ;
        RECT 4.000 60.160 295.600 61.560 ;
        RECT 4.000 58.840 296.000 60.160 ;
        RECT 4.400 57.440 295.600 58.840 ;
        RECT 4.000 56.120 296.000 57.440 ;
        RECT 4.000 54.720 295.600 56.120 ;
        RECT 4.000 54.080 296.000 54.720 ;
        RECT 4.400 53.400 296.000 54.080 ;
        RECT 4.400 52.680 295.600 53.400 ;
        RECT 4.000 52.000 295.600 52.680 ;
        RECT 4.000 50.680 296.000 52.000 ;
        RECT 4.000 49.320 295.600 50.680 ;
        RECT 4.400 49.280 295.600 49.320 ;
        RECT 4.400 48.640 296.000 49.280 ;
        RECT 4.400 47.920 295.600 48.640 ;
        RECT 4.000 47.240 295.600 47.920 ;
        RECT 4.000 45.920 296.000 47.240 ;
        RECT 4.000 45.240 295.600 45.920 ;
        RECT 4.400 44.520 295.600 45.240 ;
        RECT 4.400 43.840 296.000 44.520 ;
        RECT 4.000 43.200 296.000 43.840 ;
        RECT 4.000 41.800 295.600 43.200 ;
        RECT 4.000 40.480 296.000 41.800 ;
        RECT 4.400 39.080 295.600 40.480 ;
        RECT 4.000 37.760 296.000 39.080 ;
        RECT 4.000 36.360 295.600 37.760 ;
        RECT 4.000 35.720 296.000 36.360 ;
        RECT 4.400 35.040 296.000 35.720 ;
        RECT 4.400 34.320 295.600 35.040 ;
        RECT 4.000 33.640 295.600 34.320 ;
        RECT 4.000 33.000 296.000 33.640 ;
        RECT 4.000 31.600 295.600 33.000 ;
        RECT 4.000 30.960 296.000 31.600 ;
        RECT 4.400 30.280 296.000 30.960 ;
        RECT 4.400 29.560 295.600 30.280 ;
        RECT 4.000 28.880 295.600 29.560 ;
        RECT 4.000 27.560 296.000 28.880 ;
        RECT 4.000 26.200 295.600 27.560 ;
        RECT 4.400 26.160 295.600 26.200 ;
        RECT 4.400 24.840 296.000 26.160 ;
        RECT 4.400 24.800 295.600 24.840 ;
        RECT 4.000 23.440 295.600 24.800 ;
        RECT 4.000 22.120 296.000 23.440 ;
        RECT 4.000 21.440 295.600 22.120 ;
        RECT 4.400 20.720 295.600 21.440 ;
        RECT 4.400 20.040 296.000 20.720 ;
        RECT 4.000 19.400 296.000 20.040 ;
        RECT 4.000 18.000 295.600 19.400 ;
        RECT 4.000 17.360 296.000 18.000 ;
        RECT 4.000 16.680 295.600 17.360 ;
        RECT 4.400 15.960 295.600 16.680 ;
        RECT 4.400 15.280 296.000 15.960 ;
        RECT 4.000 14.640 296.000 15.280 ;
        RECT 4.000 13.240 295.600 14.640 ;
        RECT 4.000 11.920 296.000 13.240 ;
        RECT 4.400 10.520 295.600 11.920 ;
        RECT 4.000 9.200 296.000 10.520 ;
        RECT 4.000 7.800 295.600 9.200 ;
        RECT 4.000 7.160 296.000 7.800 ;
        RECT 4.400 6.480 296.000 7.160 ;
        RECT 4.400 5.760 295.600 6.480 ;
        RECT 4.000 5.080 295.600 5.760 ;
        RECT 4.000 3.760 296.000 5.080 ;
        RECT 4.000 3.080 295.600 3.760 ;
        RECT 4.400 2.360 295.600 3.080 ;
        RECT 4.400 1.720 296.000 2.360 ;
        RECT 4.400 1.680 295.600 1.720 ;
        RECT 4.000 0.855 295.600 1.680 ;
      LAYER met4 ;
        RECT 207.295 81.095 251.040 284.745 ;
        RECT 253.440 81.095 254.340 284.745 ;
        RECT 256.740 81.095 257.640 284.745 ;
        RECT 260.040 81.095 260.940 284.745 ;
        RECT 263.340 81.095 289.505 284.745 ;
  END
END wrapper_fibonacci
END LIBRARY

