magic
tech sky130A
magscale 1 2
timestamp 1621533840
<< locali >>
rect 52837 32351 52871 32453
rect 54217 29631 54251 29733
rect 51457 22967 51491 23137
rect 56701 10047 56735 10217
rect 53389 9367 53423 9469
rect 52193 8823 52227 8925
rect 53481 7735 53515 7837
rect 54401 7735 54435 7837
rect 6285 2975 6319 3077
<< viali >>
rect 53941 57545 53975 57579
rect 4537 57477 4571 57511
rect 53297 57477 53331 57511
rect 55505 57477 55539 57511
rect 56333 57477 56367 57511
rect 52561 57409 52595 57443
rect 1409 57341 1443 57375
rect 2053 57341 2087 57375
rect 2697 57341 2731 57375
rect 5089 57341 5123 57375
rect 5825 57341 5859 57375
rect 6929 57341 6963 57375
rect 7573 57341 7607 57375
rect 8217 57341 8251 57375
rect 9597 57341 9631 57375
rect 10241 57341 10275 57375
rect 10885 57341 10919 57375
rect 12265 57341 12299 57375
rect 12909 57341 12943 57375
rect 13553 57341 13587 57375
rect 14933 57341 14967 57375
rect 15577 57341 15611 57375
rect 16221 57341 16255 57375
rect 17601 57341 17635 57375
rect 18245 57341 18279 57375
rect 18889 57341 18923 57375
rect 20269 57341 20303 57375
rect 20913 57341 20947 57375
rect 21557 57341 21591 57375
rect 22937 57341 22971 57375
rect 23581 57341 23615 57375
rect 24225 57341 24259 57375
rect 25605 57341 25639 57375
rect 26249 57341 26283 57375
rect 26893 57341 26927 57375
rect 28273 57341 28307 57375
rect 28917 57341 28951 57375
rect 29561 57341 29595 57375
rect 30941 57341 30975 57375
rect 31585 57341 31619 57375
rect 32229 57341 32263 57375
rect 33609 57341 33643 57375
rect 34253 57341 34287 57375
rect 34897 57341 34931 57375
rect 36277 57341 36311 57375
rect 36921 57341 36955 57375
rect 37565 57341 37599 57375
rect 38945 57341 38979 57375
rect 39589 57341 39623 57375
rect 40233 57341 40267 57375
rect 42165 57341 42199 57375
rect 42993 57341 43027 57375
rect 44281 57341 44315 57375
rect 44925 57341 44959 57375
rect 45569 57341 45603 57375
rect 46949 57341 46983 57375
rect 47593 57341 47627 57375
rect 48237 57341 48271 57375
rect 49617 57341 49651 57375
rect 50261 57341 50295 57375
rect 50905 57341 50939 57375
rect 52377 57341 52411 57375
rect 55965 57341 55999 57375
rect 56149 57341 56183 57375
rect 4353 57273 4387 57307
rect 53113 57273 53147 57307
rect 53849 57273 53883 57307
rect 55321 57273 55355 57307
rect 57989 57273 58023 57307
rect 58173 57273 58207 57307
rect 5273 57205 5307 57239
rect 58173 57001 58207 57035
rect 1409 56865 1443 56899
rect 2513 56865 2547 56899
rect 16129 56865 16163 56899
rect 26433 56865 26467 56899
rect 34253 56865 34287 56899
rect 39773 56865 39807 56899
rect 40969 56865 41003 56899
rect 41613 56865 41647 56899
rect 51457 56865 51491 56899
rect 52101 56865 52135 56899
rect 52745 56865 52779 56899
rect 53665 56865 53699 56899
rect 55781 56865 55815 56899
rect 56885 56865 56919 56899
rect 4537 56797 4571 56831
rect 4721 56797 4755 56831
rect 6377 56797 6411 56831
rect 55137 56797 55171 56831
rect 57529 56797 57563 56831
rect 57713 56797 57747 56831
rect 54493 56729 54527 56763
rect 57069 56729 57103 56763
rect 3341 56661 3375 56695
rect 55597 56661 55631 56695
rect 4169 56457 4203 56491
rect 4813 56457 4847 56491
rect 5457 56457 5491 56491
rect 55045 56457 55079 56491
rect 56609 56457 56643 56491
rect 58081 56457 58115 56491
rect 2881 56389 2915 56423
rect 54401 56389 54435 56423
rect 55505 56389 55539 56423
rect 3525 56321 3559 56355
rect 3709 56321 3743 56355
rect 56333 56321 56367 56355
rect 57529 56321 57563 56355
rect 57713 56321 57747 56355
rect 1409 56253 1443 56287
rect 2053 56253 2087 56287
rect 3065 56253 3099 56287
rect 4629 56253 4663 56287
rect 51641 56253 51675 56287
rect 52285 56253 52319 56287
rect 52929 56253 52963 56287
rect 55689 56253 55723 56287
rect 56149 56253 56183 56287
rect 55597 55913 55631 55947
rect 57253 55845 57287 55879
rect 1409 55777 1443 55811
rect 4261 55777 4295 55811
rect 52377 55777 52411 55811
rect 53021 55777 53055 55811
rect 53665 55777 53699 55811
rect 54309 55777 54343 55811
rect 55781 55777 55815 55811
rect 57989 55777 58023 55811
rect 57437 55709 57471 55743
rect 58173 55641 58207 55675
rect 55137 55573 55171 55607
rect 55045 55301 55079 55335
rect 55689 55233 55723 55267
rect 57529 55233 57563 55267
rect 54217 55165 54251 55199
rect 56333 55165 56367 55199
rect 57713 55165 57747 55199
rect 58173 55165 58207 55199
rect 56885 55097 56919 55131
rect 57069 55097 57103 55131
rect 56149 55029 56183 55063
rect 55781 54825 55815 54859
rect 57345 54825 57379 54859
rect 1409 54689 1443 54723
rect 54309 54689 54343 54723
rect 55137 54689 55171 54723
rect 55597 54689 55631 54723
rect 56885 54689 56919 54723
rect 57989 54689 58023 54723
rect 56701 54621 56735 54655
rect 58173 54553 58207 54587
rect 54953 54485 54987 54519
rect 56149 54281 56183 54315
rect 57897 54281 57931 54315
rect 57529 54145 57563 54179
rect 55505 54077 55539 54111
rect 56333 54077 56367 54111
rect 57713 54077 57747 54111
rect 56885 54009 56919 54043
rect 56977 53941 57011 53975
rect 1409 53601 1443 53635
rect 55597 53601 55631 53635
rect 57069 53533 57103 53567
rect 57253 53533 57287 53567
rect 57437 53465 57471 53499
rect 56425 53193 56459 53227
rect 56885 53193 56919 53227
rect 57989 53193 58023 53227
rect 55781 53057 55815 53091
rect 57529 53057 57563 53091
rect 1409 52989 1443 53023
rect 57069 52989 57103 53023
rect 57713 52989 57747 53023
rect 57253 52649 57287 52683
rect 57437 52513 57471 52547
rect 57989 52513 58023 52547
rect 58173 52445 58207 52479
rect 57989 52105 58023 52139
rect 56149 52037 56183 52071
rect 57713 51969 57747 52003
rect 1409 51901 1443 51935
rect 55505 51901 55539 51935
rect 56333 51901 56367 51935
rect 57529 51901 57563 51935
rect 56885 51833 56919 51867
rect 57069 51833 57103 51867
rect 57713 51561 57747 51595
rect 55137 51425 55171 51459
rect 55781 51357 55815 51391
rect 57069 51357 57103 51391
rect 57253 51357 57287 51391
rect 56609 51017 56643 51051
rect 1409 50813 1443 50847
rect 56149 50813 56183 50847
rect 56793 50813 56827 50847
rect 57437 50813 57471 50847
rect 57989 50745 58023 50779
rect 58173 50745 58207 50779
rect 57253 50677 57287 50711
rect 58173 50473 58207 50507
rect 1409 50337 1443 50371
rect 56885 50337 56919 50371
rect 57529 50337 57563 50371
rect 57713 50337 57747 50371
rect 57069 50201 57103 50235
rect 55781 50133 55815 50167
rect 56701 49929 56735 49963
rect 57529 49929 57563 49963
rect 55873 49861 55907 49895
rect 57161 49793 57195 49827
rect 57345 49793 57379 49827
rect 55229 49725 55263 49759
rect 56057 49725 56091 49759
rect 56517 49725 56551 49759
rect 1409 49249 1443 49283
rect 57437 49249 57471 49283
rect 57989 49249 58023 49283
rect 58173 49249 58207 49283
rect 55781 49045 55815 49079
rect 57253 49045 57287 49079
rect 57989 48841 58023 48875
rect 57069 48773 57103 48807
rect 57529 48705 57563 48739
rect 57713 48705 57747 48739
rect 55505 48637 55539 48671
rect 56333 48637 56367 48671
rect 56885 48569 56919 48603
rect 1409 48161 1443 48195
rect 57069 48161 57103 48195
rect 57253 48093 57287 48127
rect 57437 48025 57471 48059
rect 55781 47957 55815 47991
rect 55505 47753 55539 47787
rect 56149 47685 56183 47719
rect 57069 47617 57103 47651
rect 57529 47617 57563 47651
rect 57713 47617 57747 47651
rect 55689 47549 55723 47583
rect 56333 47549 56367 47583
rect 56885 47481 56919 47515
rect 58173 47481 58207 47515
rect 1409 47073 1443 47107
rect 54309 47073 54343 47107
rect 55597 47073 55631 47107
rect 57253 47073 57287 47107
rect 57437 47073 57471 47107
rect 57989 47073 58023 47107
rect 55137 46937 55171 46971
rect 58173 46937 58207 46971
rect 55781 46869 55815 46903
rect 56977 46665 57011 46699
rect 55689 46597 55723 46631
rect 56333 46529 56367 46563
rect 56517 46529 56551 46563
rect 58173 46529 58207 46563
rect 1409 46461 1443 46495
rect 54401 46461 54435 46495
rect 55229 46461 55263 46495
rect 55873 46461 55907 46495
rect 57529 46393 57563 46427
rect 57621 46393 57655 46427
rect 55045 46121 55079 46155
rect 55597 46121 55631 46155
rect 58173 46121 58207 46155
rect 53665 45985 53699 46019
rect 54953 45985 54987 46019
rect 55137 45985 55171 46019
rect 55781 45985 55815 46019
rect 57253 45985 57287 46019
rect 57989 45985 58023 46019
rect 57437 45849 57471 45883
rect 54493 45781 54527 45815
rect 57069 45509 57103 45543
rect 57989 45509 58023 45543
rect 57529 45441 57563 45475
rect 1409 45373 1443 45407
rect 54033 45373 54067 45407
rect 54217 45373 54251 45407
rect 54861 45373 54895 45407
rect 55045 45373 55079 45407
rect 55689 45373 55723 45407
rect 56333 45373 56367 45407
rect 57713 45373 57747 45407
rect 56885 45305 56919 45339
rect 54125 45237 54159 45271
rect 54953 45237 54987 45271
rect 55505 45237 55539 45271
rect 56149 45237 56183 45271
rect 54033 45033 54067 45067
rect 57345 45033 57379 45067
rect 52265 44897 52299 44931
rect 54033 44897 54067 44931
rect 54401 44897 54435 44931
rect 54861 44897 54895 44931
rect 55597 44897 55631 44931
rect 56885 44897 56919 44931
rect 57989 44897 58023 44931
rect 52009 44829 52043 44863
rect 53849 44829 53883 44863
rect 56701 44829 56735 44863
rect 53389 44761 53423 44795
rect 55689 44761 55723 44795
rect 58173 44761 58207 44795
rect 54953 44693 54987 44727
rect 52009 44489 52043 44523
rect 52929 44489 52963 44523
rect 57989 44489 58023 44523
rect 55873 44421 55907 44455
rect 50169 44353 50203 44387
rect 57529 44353 57563 44387
rect 57713 44353 57747 44387
rect 1409 44285 1443 44319
rect 52009 44285 52043 44319
rect 52193 44285 52227 44319
rect 52929 44285 52963 44319
rect 53113 44285 53147 44319
rect 54493 44285 54527 44319
rect 50436 44217 50470 44251
rect 54760 44217 54794 44251
rect 56885 44217 56919 44251
rect 57069 44217 57103 44251
rect 51549 44149 51583 44183
rect 50445 43945 50479 43979
rect 51549 43945 51583 43979
rect 52561 43945 52595 43979
rect 55137 43945 55171 43979
rect 57529 43945 57563 43979
rect 57989 43945 58023 43979
rect 52653 43877 52687 43911
rect 50353 43809 50387 43843
rect 50537 43809 50571 43843
rect 51457 43809 51491 43843
rect 52377 43809 52411 43843
rect 52745 43809 52779 43843
rect 53481 43809 53515 43843
rect 54125 43809 54159 43843
rect 54309 43809 54343 43843
rect 54401 43809 54435 43843
rect 54585 43809 54619 43843
rect 55045 43809 55079 43843
rect 55229 43809 55263 43843
rect 56885 43809 56919 43843
rect 58173 43809 58207 43843
rect 52193 43741 52227 43775
rect 57069 43741 57103 43775
rect 53297 43673 53331 43707
rect 54217 43673 54251 43707
rect 53941 43605 53975 43639
rect 54033 43401 54067 43435
rect 54401 43333 54435 43367
rect 50537 43265 50571 43299
rect 52837 43265 52871 43299
rect 52929 43265 52963 43299
rect 54493 43265 54527 43299
rect 56977 43265 57011 43299
rect 1409 43197 1443 43231
rect 50445 43197 50479 43231
rect 51089 43197 51123 43231
rect 51273 43197 51307 43231
rect 52101 43197 52135 43231
rect 52741 43197 52775 43231
rect 53021 43197 53055 43231
rect 54217 43197 54251 43231
rect 55045 43197 55079 43231
rect 56885 43197 56919 43231
rect 55312 43129 55346 43163
rect 57989 43129 58023 43163
rect 58173 43129 58207 43163
rect 51181 43061 51215 43095
rect 52561 43061 52595 43095
rect 56425 43061 56459 43095
rect 50353 42857 50387 42891
rect 51641 42857 51675 42891
rect 58173 42857 58207 42891
rect 51457 42789 51491 42823
rect 1409 42721 1443 42755
rect 49240 42721 49274 42755
rect 51733 42721 51767 42755
rect 52929 42721 52963 42755
rect 53021 42721 53055 42755
rect 53113 42721 53147 42755
rect 53297 42721 53331 42755
rect 53757 42721 53791 42755
rect 54677 42721 54711 42755
rect 54769 42721 54803 42755
rect 55045 42721 55079 42755
rect 55505 42721 55539 42755
rect 56885 42721 56919 42755
rect 57529 42721 57563 42755
rect 48973 42653 49007 42687
rect 53849 42653 53883 42687
rect 57713 42653 57747 42687
rect 54493 42585 54527 42619
rect 55597 42585 55631 42619
rect 51457 42517 51491 42551
rect 52653 42517 52687 42551
rect 54953 42517 54987 42551
rect 56977 42517 57011 42551
rect 50997 42313 51031 42347
rect 52837 42313 52871 42347
rect 55413 42313 55447 42347
rect 55873 42313 55907 42347
rect 57161 42313 57195 42347
rect 50445 42245 50479 42279
rect 52193 42245 52227 42279
rect 50537 42177 50571 42211
rect 49433 42109 49467 42143
rect 50261 42109 50295 42143
rect 51227 42109 51261 42143
rect 51362 42109 51396 42143
rect 51478 42109 51512 42143
rect 51653 42109 51687 42143
rect 52101 42109 52135 42143
rect 52745 42109 52779 42143
rect 52929 42109 52963 42143
rect 54033 42109 54067 42143
rect 54289 42109 54323 42143
rect 55873 42109 55907 42143
rect 56057 42109 56091 42143
rect 56793 42109 56827 42143
rect 56977 42109 57011 42143
rect 57989 42041 58023 42075
rect 58173 42041 58207 42075
rect 50077 41973 50111 42007
rect 51641 41769 51675 41803
rect 52561 41769 52595 41803
rect 55597 41769 55631 41803
rect 58173 41769 58207 41803
rect 1409 41633 1443 41667
rect 50353 41633 50387 41667
rect 50537 41633 50571 41667
rect 51457 41633 51491 41667
rect 51641 41633 51675 41667
rect 52745 41633 52779 41667
rect 53389 41633 53423 41667
rect 53481 41633 53515 41667
rect 53757 41633 53791 41667
rect 54217 41633 54251 41667
rect 54861 41633 54895 41667
rect 55045 41633 55079 41667
rect 55781 41633 55815 41667
rect 56885 41633 56919 41667
rect 54309 41565 54343 41599
rect 57529 41565 57563 41599
rect 57713 41565 57747 41599
rect 50353 41497 50387 41531
rect 53205 41497 53239 41531
rect 53665 41497 53699 41531
rect 54861 41429 54895 41463
rect 57069 41429 57103 41463
rect 50905 41225 50939 41259
rect 52745 41225 52779 41259
rect 55965 41225 55999 41259
rect 51365 41021 51399 41055
rect 54585 41021 54619 41055
rect 54852 41021 54886 41055
rect 56425 41021 56459 41055
rect 51610 40953 51644 40987
rect 57253 40953 57287 40987
rect 57437 40953 57471 40987
rect 57989 40953 58023 40987
rect 56517 40885 56551 40919
rect 58081 40885 58115 40919
rect 54493 40681 54527 40715
rect 58173 40681 58207 40715
rect 50445 40613 50479 40647
rect 51917 40613 51951 40647
rect 1409 40545 1443 40579
rect 49709 40545 49743 40579
rect 50353 40545 50387 40579
rect 50537 40545 50571 40579
rect 51641 40545 51675 40579
rect 52009 40545 52043 40579
rect 53021 40545 53055 40579
rect 53481 40545 53515 40579
rect 53849 40545 53883 40579
rect 54677 40545 54711 40579
rect 55137 40545 55171 40579
rect 55321 40545 55355 40579
rect 56701 40545 56735 40579
rect 51457 40477 51491 40511
rect 53573 40477 53607 40511
rect 53757 40477 53791 40511
rect 57529 40477 57563 40511
rect 57713 40477 57747 40511
rect 51733 40409 51767 40443
rect 56793 40409 56827 40443
rect 53113 40341 53147 40375
rect 55137 40341 55171 40375
rect 52193 40137 52227 40171
rect 57529 40137 57563 40171
rect 50261 40069 50295 40103
rect 54033 40069 54067 40103
rect 52561 40001 52595 40035
rect 55321 40001 55355 40035
rect 57161 40001 57195 40035
rect 1409 39933 1443 39967
rect 50261 39933 50295 39967
rect 50445 39933 50479 39967
rect 51089 39933 51123 39967
rect 51549 39933 51583 39967
rect 51733 39933 51767 39967
rect 52377 39933 52411 39967
rect 52653 39933 52687 39967
rect 54217 39933 54251 39967
rect 54309 39933 54343 39967
rect 54493 39933 54527 39967
rect 54585 39933 54619 39967
rect 55577 39933 55611 39967
rect 57345 39933 57379 39967
rect 50905 39797 50939 39831
rect 51733 39797 51767 39831
rect 56701 39797 56735 39831
rect 51825 39593 51859 39627
rect 55689 39593 55723 39627
rect 52285 39525 52319 39559
rect 54002 39525 54036 39559
rect 51641 39457 51675 39491
rect 51825 39457 51859 39491
rect 52561 39457 52595 39491
rect 52653 39457 52687 39491
rect 52745 39457 52779 39491
rect 52929 39457 52963 39491
rect 55597 39457 55631 39491
rect 56793 39457 56827 39491
rect 58081 39457 58115 39491
rect 53757 39389 53791 39423
rect 57437 39389 57471 39423
rect 57621 39389 57655 39423
rect 55137 39321 55171 39355
rect 56977 39321 57011 39355
rect 50537 39253 50571 39287
rect 52101 39049 52135 39083
rect 52561 39049 52595 39083
rect 54861 39049 54895 39083
rect 55321 39049 55355 39083
rect 52837 38913 52871 38947
rect 52929 38913 52963 38947
rect 56701 38913 56735 38947
rect 1409 38845 1443 38879
rect 50629 38845 50663 38879
rect 51457 38845 51491 38879
rect 51917 38845 51951 38879
rect 52745 38845 52779 38879
rect 53021 38845 53055 38879
rect 54033 38845 54067 38879
rect 55045 38845 55079 38879
rect 55137 38845 55171 38879
rect 55413 38845 55447 38879
rect 56425 38845 56459 38879
rect 57989 38777 58023 38811
rect 51273 38709 51307 38743
rect 54125 38709 54159 38743
rect 58081 38709 58115 38743
rect 50445 38505 50479 38539
rect 52745 38505 52779 38539
rect 53113 38505 53147 38539
rect 53297 38505 53331 38539
rect 57253 38505 57287 38539
rect 51917 38437 51951 38471
rect 54309 38437 54343 38471
rect 50353 38369 50387 38403
rect 50537 38369 50571 38403
rect 51641 38369 51675 38403
rect 52009 38369 52043 38403
rect 53021 38369 53055 38403
rect 54493 38369 54527 38403
rect 54585 38369 54619 38403
rect 54861 38369 54895 38403
rect 55321 38369 55355 38403
rect 57437 38369 57471 38403
rect 57989 38369 58023 38403
rect 58173 38369 58207 38403
rect 51457 38301 51491 38335
rect 52929 38301 52963 38335
rect 53389 38301 53423 38335
rect 51733 38165 51767 38199
rect 54769 38165 54803 38199
rect 55413 38165 55447 38199
rect 49617 37961 49651 37995
rect 53021 37961 53055 37995
rect 54493 37961 54527 37995
rect 57989 37961 58023 37995
rect 52101 37893 52135 37927
rect 56977 37893 57011 37927
rect 54033 37825 54067 37859
rect 57529 37825 57563 37859
rect 1409 37757 1443 37791
rect 50077 37757 50111 37791
rect 50261 37757 50295 37791
rect 50721 37757 50755 37791
rect 52929 37757 52963 37791
rect 54217 37757 54251 37791
rect 55045 37757 55079 37791
rect 56885 37757 56919 37791
rect 57713 37757 57747 37791
rect 50169 37689 50203 37723
rect 50966 37689 51000 37723
rect 54585 37689 54619 37723
rect 55312 37689 55346 37723
rect 56425 37621 56459 37655
rect 50353 37417 50387 37451
rect 54953 37417 54987 37451
rect 55505 37417 55539 37451
rect 57713 37417 57747 37451
rect 54677 37349 54711 37383
rect 49065 37281 49099 37315
rect 49709 37281 49743 37315
rect 49893 37281 49927 37315
rect 50537 37281 50571 37315
rect 51917 37281 51951 37315
rect 52101 37281 52135 37315
rect 52817 37281 52851 37315
rect 54401 37281 54435 37315
rect 54585 37281 54619 37315
rect 54769 37281 54803 37315
rect 55413 37281 55447 37315
rect 55597 37281 55631 37315
rect 57253 37281 57287 37315
rect 49801 37213 49835 37247
rect 52561 37213 52595 37247
rect 57069 37213 57103 37247
rect 52009 37145 52043 37179
rect 53941 37077 53975 37111
rect 52285 36873 52319 36907
rect 56149 36873 56183 36907
rect 57253 36873 57287 36907
rect 58173 36737 58207 36771
rect 1409 36669 1443 36703
rect 50077 36669 50111 36703
rect 50333 36669 50367 36703
rect 52541 36669 52575 36703
rect 52653 36669 52687 36703
rect 52750 36669 52784 36703
rect 52929 36669 52963 36703
rect 54033 36669 54067 36703
rect 54769 36669 54803 36703
rect 56609 36669 56643 36703
rect 57437 36669 57471 36703
rect 55014 36601 55048 36635
rect 57989 36601 58023 36635
rect 51457 36533 51491 36567
rect 54125 36533 54159 36567
rect 56701 36533 56735 36567
rect 52469 36329 52503 36363
rect 53573 36329 53607 36363
rect 54677 36329 54711 36363
rect 56977 36329 57011 36363
rect 58173 36329 58207 36363
rect 1409 36193 1443 36227
rect 51549 36193 51583 36227
rect 52653 36193 52687 36227
rect 53757 36193 53791 36227
rect 53849 36193 53883 36227
rect 54125 36193 54159 36227
rect 54585 36193 54619 36227
rect 54769 36193 54803 36227
rect 55597 36193 55631 36227
rect 56885 36193 56919 36227
rect 57713 36193 57747 36227
rect 52837 36125 52871 36159
rect 52929 36125 52963 36159
rect 57529 36125 57563 36159
rect 50537 36057 50571 36091
rect 51641 35989 51675 36023
rect 54033 35989 54067 36023
rect 55689 35989 55723 36023
rect 57253 35785 57287 35819
rect 50353 35717 50387 35751
rect 57069 35649 57103 35683
rect 49709 35581 49743 35615
rect 50537 35581 50571 35615
rect 50997 35581 51031 35615
rect 51733 35581 51767 35615
rect 51917 35581 51951 35615
rect 53113 35581 53147 35615
rect 56885 35581 56919 35615
rect 57989 35581 58023 35615
rect 54493 35513 54527 35547
rect 55229 35513 55263 35547
rect 55413 35513 55447 35547
rect 56241 35513 56275 35547
rect 51089 35445 51123 35479
rect 51825 35445 51859 35479
rect 52929 35445 52963 35479
rect 54585 35445 54619 35479
rect 56333 35445 56367 35479
rect 58173 35445 58207 35479
rect 56977 35241 57011 35275
rect 49801 35173 49835 35207
rect 52070 35173 52104 35207
rect 1409 35105 1443 35139
rect 49709 35105 49743 35139
rect 49893 35105 49927 35139
rect 50537 35105 50571 35139
rect 53665 35105 53699 35139
rect 54576 35105 54610 35139
rect 56885 35105 56919 35139
rect 58173 35105 58207 35139
rect 51825 35037 51859 35071
rect 54309 35037 54343 35071
rect 57529 35037 57563 35071
rect 57713 35037 57747 35071
rect 50353 34969 50387 35003
rect 53205 34969 53239 35003
rect 53757 34901 53791 34935
rect 55689 34901 55723 34935
rect 50353 34697 50387 34731
rect 51273 34697 51307 34731
rect 52009 34697 52043 34731
rect 52929 34697 52963 34731
rect 55045 34697 55079 34731
rect 58081 34697 58115 34731
rect 49709 34629 49743 34663
rect 56425 34629 56459 34663
rect 51733 34561 51767 34595
rect 54493 34561 54527 34595
rect 57069 34561 57103 34595
rect 50169 34493 50203 34527
rect 51917 34493 51951 34527
rect 52285 34493 52319 34527
rect 54033 34493 54067 34527
rect 54217 34493 54251 34527
rect 54309 34493 54343 34527
rect 54585 34493 54619 34527
rect 55045 34493 55079 34527
rect 55241 34493 55275 34527
rect 56885 34493 56919 34527
rect 57529 34493 57563 34527
rect 57989 34493 58023 34527
rect 50905 34425 50939 34459
rect 51089 34425 51123 34459
rect 52193 34425 52227 34459
rect 52837 34425 52871 34459
rect 56241 34425 56275 34459
rect 50445 34153 50479 34187
rect 51917 34153 51951 34187
rect 56885 34153 56919 34187
rect 56793 34085 56827 34119
rect 1409 34017 1443 34051
rect 49709 34017 49743 34051
rect 50353 34017 50387 34051
rect 50537 34017 50571 34051
rect 52101 34017 52135 34051
rect 53022 34017 53056 34051
rect 53113 34017 53147 34051
rect 53389 34017 53423 34051
rect 54668 34017 54702 34051
rect 57529 34017 57563 34051
rect 52377 33949 52411 33983
rect 54401 33949 54435 33983
rect 57713 33949 57747 33983
rect 52837 33881 52871 33915
rect 55781 33881 55815 33915
rect 52285 33813 52319 33847
rect 53297 33813 53331 33847
rect 57989 33813 58023 33847
rect 49801 33609 49835 33643
rect 52009 33609 52043 33643
rect 55505 33609 55539 33643
rect 56057 33609 56091 33643
rect 50261 33541 50295 33575
rect 53113 33541 53147 33575
rect 54493 33541 54527 33575
rect 58173 33541 58207 33575
rect 1409 33405 1443 33439
rect 50261 33405 50295 33439
rect 50445 33405 50479 33439
rect 50997 33405 51031 33439
rect 51917 33405 51951 33439
rect 52561 33405 52595 33439
rect 52837 33405 52871 33439
rect 52929 33405 52963 33439
rect 54217 33405 54251 33439
rect 54355 33405 54389 33439
rect 54585 33405 54619 33439
rect 55229 33405 55263 33439
rect 55321 33405 55355 33439
rect 55597 33405 55631 33439
rect 56057 33405 56091 33439
rect 56241 33405 56275 33439
rect 57989 33405 58023 33439
rect 52745 33337 52779 33371
rect 54033 33337 54067 33371
rect 57253 33337 57287 33371
rect 51089 33269 51123 33303
rect 55045 33269 55079 33303
rect 57345 33269 57379 33303
rect 52837 33065 52871 33099
rect 53573 33065 53607 33099
rect 53481 32997 53515 33031
rect 49709 32929 49743 32963
rect 50537 32929 50571 32963
rect 51713 32929 51747 32963
rect 53665 32929 53699 32963
rect 54309 32929 54343 32963
rect 55137 32929 55171 32963
rect 55229 32929 55263 32963
rect 55505 32929 55539 32963
rect 57161 32929 57195 32963
rect 51457 32861 51491 32895
rect 54401 32861 54435 32895
rect 57345 32861 57379 32895
rect 53297 32793 53331 32827
rect 54953 32793 54987 32827
rect 57529 32793 57563 32827
rect 50353 32725 50387 32759
rect 53849 32725 53883 32759
rect 55413 32725 55447 32759
rect 51549 32521 51583 32555
rect 50997 32453 51031 32487
rect 52837 32453 52871 32487
rect 56701 32453 56735 32487
rect 54033 32385 54067 32419
rect 54309 32385 54343 32419
rect 54493 32385 54527 32419
rect 57713 32385 57747 32419
rect 1409 32317 1443 32351
rect 50905 32317 50939 32351
rect 51089 32317 51123 32351
rect 51825 32317 51859 32351
rect 51917 32317 51951 32351
rect 52009 32317 52043 32351
rect 52193 32317 52227 32351
rect 52837 32317 52871 32351
rect 52929 32317 52963 32351
rect 54217 32317 54251 32351
rect 54401 32317 54435 32351
rect 55321 32317 55355 32351
rect 57529 32317 57563 32351
rect 55566 32249 55600 32283
rect 53021 32181 53055 32215
rect 58173 32181 58207 32215
rect 51733 31977 51767 32011
rect 54125 31977 54159 32011
rect 55045 31909 55079 31943
rect 55137 31909 55171 31943
rect 57989 31909 58023 31943
rect 58173 31909 58207 31943
rect 49893 31841 49927 31875
rect 50537 31841 50571 31875
rect 52009 31841 52043 31875
rect 53001 31841 53035 31875
rect 54861 31841 54895 31875
rect 55229 31841 55263 31875
rect 57253 31841 57287 31875
rect 51917 31773 51951 31807
rect 52101 31773 52135 31807
rect 52193 31773 52227 31807
rect 52745 31773 52779 31807
rect 57437 31773 57471 31807
rect 49709 31705 49743 31739
rect 55413 31637 55447 31671
rect 50813 31433 50847 31467
rect 54401 31433 54435 31467
rect 54769 31433 54803 31467
rect 58081 31433 58115 31467
rect 49341 31365 49375 31399
rect 52929 31365 52963 31399
rect 1409 31229 1443 31263
rect 49525 31229 49559 31263
rect 49985 31229 50019 31263
rect 52285 31229 52319 31263
rect 52469 31229 52503 31263
rect 53113 31229 53147 31263
rect 54585 31229 54619 31263
rect 54861 31229 54895 31263
rect 55321 31229 55355 31263
rect 57437 31229 57471 31263
rect 57621 31229 57655 31263
rect 51365 31161 51399 31195
rect 55588 31161 55622 31195
rect 51457 31093 51491 31127
rect 52469 31093 52503 31127
rect 56701 31093 56735 31127
rect 50445 30889 50479 30923
rect 52193 30889 52227 30923
rect 54309 30889 54343 30923
rect 55413 30889 55447 30923
rect 1409 30753 1443 30787
rect 49709 30753 49743 30787
rect 50353 30753 50387 30787
rect 50537 30753 50571 30787
rect 51733 30753 51767 30787
rect 52423 30753 52457 30787
rect 52542 30753 52576 30787
rect 52653 30753 52687 30787
rect 52837 30753 52871 30787
rect 53573 30753 53607 30787
rect 53757 30753 53791 30787
rect 53849 30753 53883 30787
rect 54493 30753 54527 30787
rect 54585 30753 54619 30787
rect 54861 30753 54895 30787
rect 55321 30753 55355 30787
rect 55505 30753 55539 30787
rect 57253 30753 57287 30787
rect 57989 30753 58023 30787
rect 51549 30617 51583 30651
rect 53389 30617 53423 30651
rect 54769 30617 54803 30651
rect 57437 30617 57471 30651
rect 58173 30617 58207 30651
rect 52929 30345 52963 30379
rect 53113 30345 53147 30379
rect 55137 30345 55171 30379
rect 55689 30345 55723 30379
rect 57989 30345 58023 30379
rect 52009 30277 52043 30311
rect 56793 30277 56827 30311
rect 49525 30209 49559 30243
rect 54033 30209 54067 30243
rect 54585 30209 54619 30243
rect 57529 30209 57563 30243
rect 49065 30141 49099 30175
rect 51917 30141 51951 30175
rect 52561 30141 52595 30175
rect 54217 30141 54251 30175
rect 54447 30141 54481 30175
rect 55045 30141 55079 30175
rect 55689 30141 55723 30175
rect 55873 30141 55907 30175
rect 57713 30141 57747 30175
rect 1869 30073 1903 30107
rect 49770 30073 49804 30107
rect 52929 30073 52963 30107
rect 56609 30073 56643 30107
rect 1961 30005 1995 30039
rect 48881 30005 48915 30039
rect 50905 30005 50939 30039
rect 54401 30005 54435 30039
rect 48697 29801 48731 29835
rect 49433 29801 49467 29835
rect 57989 29801 58023 29835
rect 50445 29733 50479 29767
rect 52653 29733 52687 29767
rect 53297 29733 53331 29767
rect 54217 29733 54251 29767
rect 1869 29665 1903 29699
rect 48881 29665 48915 29699
rect 49341 29665 49375 29699
rect 49525 29665 49559 29699
rect 50169 29665 50203 29699
rect 51457 29665 51491 29699
rect 52377 29665 52411 29699
rect 52745 29665 52779 29699
rect 53205 29665 53239 29699
rect 54565 29665 54599 29699
rect 57069 29665 57103 29699
rect 58173 29665 58207 29699
rect 49985 29597 50019 29631
rect 50537 29597 50571 29631
rect 52285 29597 52319 29631
rect 54217 29597 54251 29631
rect 54309 29597 54343 29631
rect 56885 29597 56919 29631
rect 50261 29529 50295 29563
rect 55689 29529 55723 29563
rect 57253 29529 57287 29563
rect 1961 29461 1995 29495
rect 2697 29461 2731 29495
rect 51549 29461 51583 29495
rect 1961 29257 1995 29291
rect 47685 29257 47719 29291
rect 48973 29257 49007 29291
rect 50077 29257 50111 29291
rect 54033 29257 54067 29291
rect 55781 29257 55815 29291
rect 57253 29257 57287 29291
rect 50537 29189 50571 29223
rect 56517 29189 56551 29223
rect 1593 29121 1627 29155
rect 49525 29121 49559 29155
rect 52469 29121 52503 29155
rect 52745 29121 52779 29155
rect 1777 29053 1811 29087
rect 47869 29053 47903 29087
rect 49433 29053 49467 29087
rect 49617 29053 49651 29087
rect 50261 29053 50295 29087
rect 50353 29053 50387 29087
rect 50629 29053 50663 29087
rect 51457 29053 51491 29087
rect 51549 29053 51583 29087
rect 51733 29053 51767 29087
rect 51825 29053 51859 29087
rect 52285 29053 52319 29087
rect 52837 29053 52871 29087
rect 54033 29053 54067 29087
rect 54217 29053 54251 29087
rect 54953 29053 54987 29087
rect 55137 29053 55171 29087
rect 55965 29053 55999 29087
rect 56425 29053 56459 29087
rect 57437 29053 57471 29087
rect 55045 28985 55079 29019
rect 57989 28985 58023 29019
rect 58173 28985 58207 29019
rect 51273 28917 51307 28951
rect 47777 28713 47811 28747
rect 50445 28713 50479 28747
rect 52469 28713 52503 28747
rect 55229 28713 55263 28747
rect 58173 28713 58207 28747
rect 1777 28577 1811 28611
rect 47317 28577 47351 28611
rect 47961 28577 47995 28611
rect 48421 28577 48455 28611
rect 49065 28577 49099 28611
rect 49249 28577 49283 28611
rect 49709 28577 49743 28611
rect 49893 28577 49927 28611
rect 50353 28577 50387 28611
rect 51733 28577 51767 28611
rect 51917 28577 51951 28611
rect 52101 28577 52135 28611
rect 52285 28577 52319 28611
rect 53553 28577 53587 28611
rect 55137 28577 55171 28611
rect 56885 28577 56919 28611
rect 57069 28577 57103 28611
rect 57529 28577 57563 28611
rect 1961 28509 1995 28543
rect 49801 28509 49835 28543
rect 52009 28509 52043 28543
rect 53297 28509 53331 28543
rect 57713 28509 57747 28543
rect 2145 28441 2179 28475
rect 49065 28441 49099 28475
rect 47133 28373 47167 28407
rect 54677 28373 54711 28407
rect 2513 28169 2547 28203
rect 3157 28169 3191 28203
rect 3985 28169 4019 28203
rect 50169 28169 50203 28203
rect 52469 28169 52503 28203
rect 57437 28169 57471 28203
rect 52009 28101 52043 28135
rect 54401 28101 54435 28135
rect 54493 28033 54527 28067
rect 2697 27965 2731 27999
rect 3341 27965 3375 27999
rect 48789 27965 48823 27999
rect 50629 27965 50663 27999
rect 50813 27965 50847 27999
rect 51825 27965 51859 27999
rect 52745 27965 52779 27999
rect 52834 27965 52868 27999
rect 52929 27965 52963 27999
rect 53113 27965 53147 27999
rect 54217 27965 54251 27999
rect 55137 27965 55171 27999
rect 55393 27965 55427 27999
rect 57069 27965 57103 27999
rect 57253 27965 57287 27999
rect 1869 27897 1903 27931
rect 49056 27897 49090 27931
rect 51641 27897 51675 27931
rect 1961 27829 1995 27863
rect 50721 27829 50755 27863
rect 54033 27829 54067 27863
rect 56517 27829 56551 27863
rect 50537 27625 50571 27659
rect 51457 27625 51491 27659
rect 53481 27625 53515 27659
rect 54125 27557 54159 27591
rect 57069 27557 57103 27591
rect 1685 27489 1719 27523
rect 48605 27489 48639 27523
rect 49065 27489 49099 27523
rect 49249 27489 49283 27523
rect 49893 27489 49927 27523
rect 50353 27489 50387 27523
rect 50537 27489 50571 27523
rect 51641 27489 51675 27523
rect 51917 27489 51951 27523
rect 52561 27489 52595 27523
rect 52653 27489 52687 27523
rect 53389 27489 53423 27523
rect 54309 27489 54343 27523
rect 54401 27489 54435 27523
rect 54677 27489 54711 27523
rect 55321 27489 55355 27523
rect 55505 27489 55539 27523
rect 55689 27489 55723 27523
rect 56885 27489 56919 27523
rect 58173 27489 58207 27523
rect 1869 27421 1903 27455
rect 52745 27421 52779 27455
rect 52837 27421 52871 27455
rect 54585 27421 54619 27455
rect 57529 27421 57563 27455
rect 57713 27421 57747 27455
rect 2053 27353 2087 27387
rect 55321 27353 55355 27387
rect 48421 27285 48455 27319
rect 49065 27285 49099 27319
rect 49709 27285 49743 27319
rect 51825 27285 51859 27319
rect 52377 27285 52411 27319
rect 2513 27081 2547 27115
rect 3341 27081 3375 27115
rect 54125 27081 54159 27115
rect 55321 27081 55355 27115
rect 52561 26945 52595 26979
rect 53113 26945 53147 26979
rect 2697 26877 2731 26911
rect 49249 26877 49283 26911
rect 51365 26877 51399 26911
rect 51454 26877 51488 26911
rect 51549 26877 51583 26911
rect 51733 26877 51767 26911
rect 52745 26877 52779 26911
rect 54033 26877 54067 26911
rect 54769 26877 54803 26911
rect 55137 26877 55171 26911
rect 56149 26877 56183 26911
rect 57161 26877 57195 26911
rect 57345 26877 57379 26911
rect 1869 26809 1903 26843
rect 49516 26809 49550 26843
rect 51089 26809 51123 26843
rect 54953 26809 54987 26843
rect 55045 26809 55079 26843
rect 1961 26741 1995 26775
rect 50629 26741 50663 26775
rect 52929 26741 52963 26775
rect 53021 26741 53055 26775
rect 56241 26741 56275 26775
rect 57805 26741 57839 26775
rect 2329 26537 2363 26571
rect 49709 26537 49743 26571
rect 51457 26537 51491 26571
rect 54309 26537 54343 26571
rect 57345 26537 57379 26571
rect 57253 26469 57287 26503
rect 1685 26401 1719 26435
rect 2973 26401 3007 26435
rect 49893 26401 49927 26435
rect 50353 26401 50387 26435
rect 51641 26401 51675 26435
rect 51733 26401 51767 26435
rect 52009 26401 52043 26435
rect 52929 26401 52963 26435
rect 53196 26401 53230 26435
rect 54953 26401 54987 26435
rect 55045 26401 55079 26435
rect 55321 26401 55355 26435
rect 57989 26401 58023 26435
rect 1869 26333 1903 26367
rect 50445 26333 50479 26367
rect 54769 26333 54803 26367
rect 49249 26265 49283 26299
rect 58173 26265 58207 26299
rect 51917 26197 51951 26231
rect 55229 26197 55263 26231
rect 2513 25993 2547 26027
rect 52009 25993 52043 26027
rect 52561 25993 52595 26027
rect 57989 25993 58023 26027
rect 56333 25925 56367 25959
rect 2697 25789 2731 25823
rect 3341 25789 3375 25823
rect 49341 25789 49375 25823
rect 49985 25789 50019 25823
rect 50169 25789 50203 25823
rect 50629 25789 50663 25823
rect 52469 25789 52503 25823
rect 54309 25789 54343 25823
rect 54953 25789 54987 25823
rect 56793 25789 56827 25823
rect 57529 25789 57563 25823
rect 57713 25789 57747 25823
rect 1869 25721 1903 25755
rect 2053 25721 2087 25755
rect 50077 25721 50111 25755
rect 50874 25721 50908 25755
rect 55198 25721 55232 25755
rect 54401 25653 54435 25687
rect 56885 25653 56919 25687
rect 2513 25449 2547 25483
rect 54125 25449 54159 25483
rect 55137 25449 55171 25483
rect 52837 25381 52871 25415
rect 58173 25381 58207 25415
rect 1869 25313 1903 25347
rect 3157 25313 3191 25347
rect 50353 25313 50387 25347
rect 50537 25313 50571 25347
rect 51733 25313 51767 25347
rect 52377 25313 52411 25347
rect 55045 25313 55079 25347
rect 55229 25313 55263 25347
rect 56793 25313 56827 25347
rect 57437 25313 57471 25347
rect 57989 25313 58023 25347
rect 2053 25245 2087 25279
rect 49893 25245 49927 25279
rect 56977 25245 57011 25279
rect 2973 25177 3007 25211
rect 51549 25177 51583 25211
rect 50353 25109 50387 25143
rect 52193 25109 52227 25143
rect 2789 24769 2823 24803
rect 54125 24769 54159 24803
rect 54953 24769 54987 24803
rect 3433 24701 3467 24735
rect 49525 24701 49559 24735
rect 50169 24701 50203 24735
rect 51733 24701 51767 24735
rect 54033 24701 54067 24735
rect 54217 24701 54251 24735
rect 57253 24701 57287 24735
rect 1869 24633 1903 24667
rect 2605 24633 2639 24667
rect 50905 24633 50939 24667
rect 51089 24633 51123 24667
rect 52000 24633 52034 24667
rect 55198 24633 55232 24667
rect 57989 24633 58023 24667
rect 58173 24633 58207 24667
rect 1961 24565 1995 24599
rect 3249 24565 3283 24599
rect 50353 24565 50387 24599
rect 53113 24565 53147 24599
rect 56333 24565 56367 24599
rect 57437 24565 57471 24599
rect 2329 24361 2363 24395
rect 51917 24361 51951 24395
rect 54401 24361 54435 24395
rect 58173 24361 58207 24395
rect 53021 24293 53055 24327
rect 53665 24293 53699 24327
rect 1685 24225 1719 24259
rect 2973 24225 3007 24259
rect 52101 24225 52135 24259
rect 52745 24225 52779 24259
rect 53573 24225 53607 24259
rect 53757 24225 53791 24259
rect 54401 24225 54435 24259
rect 54769 24225 54803 24259
rect 55229 24225 55263 24259
rect 56885 24225 56919 24259
rect 1869 24157 1903 24191
rect 52561 24157 52595 24191
rect 53113 24157 53147 24191
rect 54217 24157 54251 24191
rect 57529 24157 57563 24191
rect 57713 24157 57747 24191
rect 50537 24089 50571 24123
rect 52837 24021 52871 24055
rect 55321 24021 55355 24055
rect 56977 24021 57011 24055
rect 2053 23817 2087 23851
rect 50537 23817 50571 23851
rect 52469 23817 52503 23851
rect 54033 23817 54067 23851
rect 54953 23817 54987 23851
rect 51825 23749 51859 23783
rect 1685 23681 1719 23715
rect 2973 23681 3007 23715
rect 1869 23613 1903 23647
rect 49249 23613 49283 23647
rect 50077 23613 50111 23647
rect 50721 23613 50755 23647
rect 51181 23613 51215 23647
rect 52009 23613 52043 23647
rect 52469 23613 52503 23647
rect 52653 23613 52687 23647
rect 54217 23613 54251 23647
rect 54401 23613 54435 23647
rect 54493 23613 54527 23647
rect 54953 23613 54987 23647
rect 55137 23613 55171 23647
rect 55965 23613 55999 23647
rect 57253 23545 57287 23579
rect 57437 23545 57471 23579
rect 57989 23545 58023 23579
rect 49893 23477 49927 23511
rect 51365 23477 51399 23511
rect 56057 23477 56091 23511
rect 58081 23477 58115 23511
rect 2513 23273 2547 23307
rect 50445 23205 50479 23239
rect 1869 23137 1903 23171
rect 2697 23137 2731 23171
rect 50353 23137 50387 23171
rect 50537 23137 50571 23171
rect 51457 23137 51491 23171
rect 51733 23137 51767 23171
rect 52449 23137 52483 23171
rect 54493 23137 54527 23171
rect 54769 23137 54803 23171
rect 54953 23137 54987 23171
rect 55597 23137 55631 23171
rect 57161 23137 57195 23171
rect 57345 23137 57379 23171
rect 3341 23001 3375 23035
rect 52193 23069 52227 23103
rect 54677 23069 54711 23103
rect 54309 23001 54343 23035
rect 54585 23001 54619 23035
rect 55689 23001 55723 23035
rect 57529 23001 57563 23035
rect 1961 22933 1995 22967
rect 51457 22933 51491 22967
rect 51549 22933 51583 22967
rect 53573 22933 53607 22967
rect 1961 22729 1995 22763
rect 2881 22729 2915 22763
rect 51549 22729 51583 22763
rect 52101 22729 52135 22763
rect 56241 22729 56275 22763
rect 57345 22729 57379 22763
rect 3341 22661 3375 22695
rect 50813 22661 50847 22695
rect 1593 22593 1627 22627
rect 1777 22593 1811 22627
rect 50261 22593 50295 22627
rect 2697 22525 2731 22559
rect 3525 22525 3559 22559
rect 50169 22525 50203 22559
rect 50353 22525 50387 22559
rect 50997 22525 51031 22559
rect 51457 22525 51491 22559
rect 51641 22525 51675 22559
rect 52377 22525 52411 22559
rect 52466 22525 52500 22559
rect 52561 22525 52595 22559
rect 52745 22525 52779 22559
rect 54125 22525 54159 22559
rect 54861 22525 54895 22559
rect 56977 22525 57011 22559
rect 57161 22525 57195 22559
rect 55106 22457 55140 22491
rect 54217 22389 54251 22423
rect 54953 22185 54987 22219
rect 2605 22117 2639 22151
rect 51549 22117 51583 22151
rect 56885 22117 56919 22151
rect 1869 22049 1903 22083
rect 49249 22049 49283 22083
rect 49709 22049 49743 22083
rect 51733 22049 51767 22083
rect 52653 22049 52687 22083
rect 52837 22049 52871 22083
rect 53849 22049 53883 22083
rect 54033 22049 54067 22083
rect 54125 22049 54159 22083
rect 54401 22049 54435 22083
rect 54861 22049 54895 22083
rect 55045 22049 55079 22083
rect 55505 22049 55539 22083
rect 55689 22049 55723 22083
rect 2881 21981 2915 22015
rect 50537 21981 50571 22015
rect 57529 21981 57563 22015
rect 57713 21981 57747 22015
rect 2053 21913 2087 21947
rect 54309 21913 54343 21947
rect 57989 21913 58023 21947
rect 49065 21845 49099 21879
rect 52745 21845 52779 21879
rect 55505 21845 55539 21879
rect 56977 21845 57011 21879
rect 2053 21641 2087 21675
rect 4261 21641 4295 21675
rect 52469 21641 52503 21675
rect 58081 21641 58115 21675
rect 52837 21573 52871 21607
rect 1685 21505 1719 21539
rect 54309 21505 54343 21539
rect 54493 21505 54527 21539
rect 57713 21505 57747 21539
rect 1869 21437 1903 21471
rect 2973 21437 3007 21471
rect 3617 21437 3651 21471
rect 49893 21437 49927 21471
rect 50077 21437 50111 21471
rect 50537 21437 50571 21471
rect 52653 21437 52687 21471
rect 52745 21437 52779 21471
rect 52929 21437 52963 21471
rect 54217 21437 54251 21471
rect 55137 21437 55171 21471
rect 57529 21437 57563 21471
rect 50782 21369 50816 21403
rect 55404 21369 55438 21403
rect 2789 21301 2823 21335
rect 49985 21301 50019 21335
rect 51917 21301 51951 21335
rect 54493 21301 54527 21335
rect 56517 21301 56551 21335
rect 49065 21097 49099 21131
rect 54493 21097 54527 21131
rect 50445 21029 50479 21063
rect 53297 21029 53331 21063
rect 1869 20961 1903 20995
rect 2605 20961 2639 20995
rect 2789 20961 2823 20995
rect 48605 20961 48639 20995
rect 49249 20961 49283 20995
rect 49893 20961 49927 20995
rect 50353 20961 50387 20995
rect 50537 20961 50571 20995
rect 51917 20961 51951 20995
rect 52653 20961 52687 20995
rect 52837 20961 52871 20995
rect 52929 20961 52963 20995
rect 53757 20961 53791 20995
rect 53941 20961 53975 20995
rect 54309 20961 54343 20995
rect 55229 20961 55263 20995
rect 55321 20961 55355 20995
rect 55597 20961 55631 20995
rect 57069 20961 57103 20995
rect 54033 20893 54067 20927
rect 54125 20893 54159 20927
rect 57253 20893 57287 20927
rect 49709 20825 49743 20859
rect 1961 20757 1995 20791
rect 48421 20757 48455 20791
rect 52009 20757 52043 20791
rect 55045 20757 55079 20791
rect 55505 20757 55539 20791
rect 57437 20757 57471 20791
rect 2421 20553 2455 20587
rect 3249 20553 3283 20587
rect 49893 20553 49927 20587
rect 51273 20553 51307 20587
rect 54861 20553 54895 20587
rect 55413 20553 55447 20587
rect 50353 20485 50387 20519
rect 57437 20485 57471 20519
rect 1961 20417 1995 20451
rect 52837 20417 52871 20451
rect 53021 20417 53055 20451
rect 56149 20417 56183 20451
rect 1777 20349 1811 20383
rect 3433 20349 3467 20383
rect 4077 20349 4111 20383
rect 49065 20349 49099 20383
rect 50537 20349 50571 20383
rect 50997 20349 51031 20383
rect 51181 20349 51215 20383
rect 51549 20349 51583 20383
rect 52745 20349 52779 20383
rect 52920 20349 52954 20383
rect 54309 20349 54343 20383
rect 54585 20349 54619 20383
rect 54677 20349 54711 20383
rect 55321 20349 55355 20383
rect 56057 20349 56091 20383
rect 57253 20349 57287 20383
rect 54493 20281 54527 20315
rect 57989 20281 58023 20315
rect 58173 20281 58207 20315
rect 3893 20213 3927 20247
rect 51457 20213 51491 20247
rect 52561 20213 52595 20247
rect 2421 20009 2455 20043
rect 52193 20009 52227 20043
rect 58173 20009 58207 20043
rect 1961 19873 1995 19907
rect 2881 19873 2915 19907
rect 49249 19873 49283 19907
rect 49893 19873 49927 19907
rect 50537 19873 50571 19907
rect 51549 19873 51583 19907
rect 52377 19873 52411 19907
rect 52561 19873 52595 19907
rect 53113 19873 53147 19907
rect 53380 19873 53414 19907
rect 54953 19873 54987 19907
rect 55137 19873 55171 19907
rect 55597 19873 55631 19907
rect 56885 19873 56919 19907
rect 57529 19873 57563 19907
rect 1777 19805 1811 19839
rect 52653 19805 52687 19839
rect 57713 19805 57747 19839
rect 4445 19737 4479 19771
rect 57069 19737 57103 19771
rect 3065 19669 3099 19703
rect 49065 19669 49099 19703
rect 50353 19669 50387 19703
rect 51641 19669 51675 19703
rect 54493 19669 54527 19703
rect 54953 19669 54987 19703
rect 55689 19669 55723 19703
rect 49617 19465 49651 19499
rect 56333 19465 56367 19499
rect 57345 19465 57379 19499
rect 3433 19261 3467 19295
rect 47869 19261 47903 19295
rect 49157 19261 49191 19295
rect 49801 19261 49835 19295
rect 50261 19261 50295 19295
rect 52745 19261 52779 19295
rect 52834 19261 52868 19295
rect 52929 19261 52963 19295
rect 53113 19261 53147 19295
rect 54309 19261 54343 19295
rect 54953 19261 54987 19295
rect 55220 19261 55254 19295
rect 56977 19261 57011 19295
rect 57161 19261 57195 19295
rect 1869 19193 1903 19227
rect 2605 19193 2639 19227
rect 2789 19193 2823 19227
rect 50528 19193 50562 19227
rect 52469 19193 52503 19227
rect 54401 19193 54435 19227
rect 1961 19125 1995 19159
rect 47685 19125 47719 19159
rect 48973 19125 49007 19159
rect 51641 19125 51675 19159
rect 2605 18921 2639 18955
rect 49065 18921 49099 18955
rect 1961 18785 1995 18819
rect 3249 18785 3283 18819
rect 49249 18785 49283 18819
rect 49709 18785 49743 18819
rect 50353 18785 50387 18819
rect 50537 18785 50571 18819
rect 51641 18785 51675 18819
rect 52561 18785 52595 18819
rect 52929 18785 52963 18819
rect 54125 18785 54159 18819
rect 54217 18785 54251 18819
rect 54493 18785 54527 18819
rect 54953 18785 54987 18819
rect 55597 18785 55631 18819
rect 56793 18785 56827 18819
rect 57989 18785 58023 18819
rect 2145 18717 2179 18751
rect 52377 18717 52411 18751
rect 3065 18649 3099 18683
rect 50353 18649 50387 18683
rect 55137 18649 55171 18683
rect 56977 18649 57011 18683
rect 58173 18649 58207 18683
rect 51733 18581 51767 18615
rect 52837 18581 52871 18615
rect 53941 18581 53975 18615
rect 54401 18581 54435 18615
rect 55689 18581 55723 18615
rect 1961 18377 1995 18411
rect 50629 18377 50663 18411
rect 56149 18377 56183 18411
rect 57989 18377 58023 18411
rect 51917 18309 51951 18343
rect 54125 18309 54159 18343
rect 1593 18241 1627 18275
rect 2881 18241 2915 18275
rect 51365 18241 51399 18275
rect 54769 18241 54803 18275
rect 57713 18241 57747 18275
rect 1777 18173 1811 18207
rect 49985 18173 50019 18207
rect 50169 18173 50203 18207
rect 50813 18173 50847 18207
rect 51273 18173 51307 18207
rect 51917 18173 51951 18207
rect 52101 18173 52135 18207
rect 52561 18173 52595 18207
rect 52745 18173 52779 18207
rect 52837 18173 52871 18207
rect 53021 18173 53055 18207
rect 53113 18173 53147 18207
rect 54033 18173 54067 18207
rect 54217 18173 54251 18207
rect 57529 18173 57563 18207
rect 50077 18105 50111 18139
rect 55014 18105 55048 18139
rect 56885 18105 56919 18139
rect 57069 18105 57103 18139
rect 2513 17833 2547 17867
rect 49709 17833 49743 17867
rect 54861 17833 54895 17867
rect 1869 17697 1903 17731
rect 2697 17697 2731 17731
rect 49893 17697 49927 17731
rect 50353 17697 50387 17731
rect 50537 17697 50571 17731
rect 51641 17697 51675 17731
rect 51733 17697 51767 17731
rect 52009 17697 52043 17731
rect 52469 17697 52503 17731
rect 52653 17697 52687 17731
rect 52837 17697 52871 17731
rect 53021 17697 53055 17731
rect 53205 17697 53239 17731
rect 53941 17697 53975 17731
rect 54030 17697 54064 17731
rect 54125 17697 54159 17731
rect 54309 17697 54343 17731
rect 54769 17697 54803 17731
rect 54953 17697 54987 17731
rect 55505 17697 55539 17731
rect 51917 17629 51951 17663
rect 52745 17629 52779 17663
rect 55597 17629 55631 17663
rect 56977 17629 57011 17663
rect 57161 17629 57195 17663
rect 49249 17561 49283 17595
rect 50445 17561 50479 17595
rect 57345 17561 57379 17595
rect 1961 17493 1995 17527
rect 51457 17493 51491 17527
rect 53665 17493 53699 17527
rect 1961 17289 1995 17323
rect 55505 17289 55539 17323
rect 55965 17289 55999 17323
rect 51181 17221 51215 17255
rect 56425 17221 56459 17255
rect 1593 17153 1627 17187
rect 2881 17153 2915 17187
rect 49801 17153 49835 17187
rect 51641 17153 51675 17187
rect 52193 17153 52227 17187
rect 53113 17153 53147 17187
rect 1777 17085 1811 17119
rect 49157 17085 49191 17119
rect 51825 17085 51859 17119
rect 52837 17085 52871 17119
rect 53021 17085 53055 17119
rect 54125 17085 54159 17119
rect 54381 17085 54415 17119
rect 56149 17085 56183 17119
rect 56241 17085 56275 17119
rect 56517 17085 56551 17119
rect 50068 17017 50102 17051
rect 52101 17017 52135 17051
rect 52653 17017 52687 17051
rect 57253 17017 57287 17051
rect 57437 17017 57471 17051
rect 57989 17017 58023 17051
rect 58173 17017 58207 17051
rect 52009 16949 52043 16983
rect 2513 16745 2547 16779
rect 49709 16745 49743 16779
rect 50445 16745 50479 16779
rect 51641 16745 51675 16779
rect 52929 16745 52963 16779
rect 54677 16745 54711 16779
rect 58173 16745 58207 16779
rect 52101 16677 52135 16711
rect 55321 16677 55355 16711
rect 1869 16609 1903 16643
rect 2697 16609 2731 16643
rect 3341 16609 3375 16643
rect 49893 16609 49927 16643
rect 50353 16609 50387 16643
rect 50537 16609 50571 16643
rect 51457 16609 51491 16643
rect 51641 16609 51675 16643
rect 52285 16609 52319 16643
rect 53113 16609 53147 16643
rect 53389 16609 53423 16643
rect 53941 16609 53975 16643
rect 54585 16609 54619 16643
rect 55229 16609 55263 16643
rect 56701 16609 56735 16643
rect 57713 16609 57747 16643
rect 53205 16541 53239 16575
rect 53297 16541 53331 16575
rect 57529 16541 57563 16575
rect 49249 16473 49283 16507
rect 1961 16405 1995 16439
rect 3157 16405 3191 16439
rect 52469 16405 52503 16439
rect 54033 16405 54067 16439
rect 56885 16405 56919 16439
rect 2237 16201 2271 16235
rect 49617 16201 49651 16235
rect 57437 16201 57471 16235
rect 4721 16133 4755 16167
rect 1869 16065 1903 16099
rect 2053 16065 2087 16099
rect 52561 16065 52595 16099
rect 52653 16065 52687 16099
rect 54033 16065 54067 16099
rect 57253 16065 57287 16099
rect 3433 15997 3467 16031
rect 4077 15997 4111 16031
rect 49801 15997 49835 16031
rect 50261 15997 50295 16031
rect 50997 15997 51031 16031
rect 52101 15997 52135 16031
rect 55965 15997 55999 16031
rect 57069 15997 57103 16031
rect 51181 15929 51215 15963
rect 54278 15929 54312 15963
rect 56333 15929 56367 15963
rect 3249 15861 3283 15895
rect 50445 15861 50479 15895
rect 52285 15861 52319 15895
rect 55413 15861 55447 15895
rect 52837 15657 52871 15691
rect 56885 15657 56919 15691
rect 50445 15589 50479 15623
rect 51917 15589 51951 15623
rect 1869 15521 1903 15555
rect 2605 15521 2639 15555
rect 49709 15521 49743 15555
rect 50353 15521 50387 15555
rect 50537 15521 50571 15555
rect 51641 15521 51675 15555
rect 52009 15521 52043 15555
rect 53067 15521 53101 15555
rect 53202 15521 53236 15555
rect 53297 15521 53331 15555
rect 53481 15521 53515 15555
rect 53941 15521 53975 15555
rect 55045 15521 55079 15555
rect 56701 15521 56735 15555
rect 57989 15521 58023 15555
rect 51457 15453 51491 15487
rect 2789 15385 2823 15419
rect 1961 15317 1995 15351
rect 51733 15317 51767 15351
rect 54033 15317 54067 15351
rect 55137 15317 55171 15351
rect 58081 15317 58115 15351
rect 2421 15113 2455 15147
rect 3065 15113 3099 15147
rect 49985 15113 50019 15147
rect 52285 15113 52319 15147
rect 54585 15113 54619 15147
rect 57989 15113 58023 15147
rect 1777 14977 1811 15011
rect 1961 14977 1995 15011
rect 50445 14977 50479 15011
rect 57713 14977 57747 15011
rect 2881 14909 2915 14943
rect 52469 14909 52503 14943
rect 52653 14909 52687 14943
rect 52745 14909 52779 14943
rect 54309 14909 54343 14943
rect 54493 14909 54527 14943
rect 55137 14909 55171 14943
rect 57529 14909 57563 14943
rect 50712 14841 50746 14875
rect 54677 14841 54711 14875
rect 55382 14841 55416 14875
rect 51825 14773 51859 14807
rect 56517 14773 56551 14807
rect 2513 14569 2547 14603
rect 54217 14569 54251 14603
rect 49801 14501 49835 14535
rect 49709 14433 49743 14467
rect 49893 14433 49927 14467
rect 50537 14433 50571 14467
rect 51457 14433 51491 14467
rect 51641 14433 51675 14467
rect 52377 14433 52411 14467
rect 52644 14433 52678 14467
rect 54401 14433 54435 14467
rect 54493 14433 54527 14467
rect 54769 14433 54803 14467
rect 55413 14433 55447 14467
rect 55505 14433 55539 14467
rect 55781 14433 55815 14467
rect 57253 14433 57287 14467
rect 1869 14365 1903 14399
rect 2053 14365 2087 14399
rect 57437 14365 57471 14399
rect 51457 14297 51491 14331
rect 53757 14297 53791 14331
rect 55689 14297 55723 14331
rect 50353 14229 50387 14263
rect 54677 14229 54711 14263
rect 55229 14229 55263 14263
rect 57621 14229 57655 14263
rect 2513 14025 2547 14059
rect 3985 14025 4019 14059
rect 51917 14025 51951 14059
rect 52561 14025 52595 14059
rect 54769 13957 54803 13991
rect 55505 13957 55539 13991
rect 57897 13957 57931 13991
rect 2697 13821 2731 13855
rect 3341 13821 3375 13855
rect 49157 13821 49191 13855
rect 49801 13821 49835 13855
rect 50445 13821 50479 13855
rect 50629 13821 50663 13855
rect 51365 13821 51399 13855
rect 52101 13821 52135 13855
rect 52561 13821 52595 13855
rect 52745 13821 52779 13855
rect 54217 13821 54251 13855
rect 54401 13821 54435 13855
rect 54585 13821 54619 13855
rect 55321 13821 55355 13855
rect 56057 13821 56091 13855
rect 56885 13821 56919 13855
rect 57069 13821 57103 13855
rect 57529 13821 57563 13855
rect 57713 13821 57747 13855
rect 1869 13753 1903 13787
rect 51181 13753 51215 13787
rect 54493 13753 54527 13787
rect 1961 13685 1995 13719
rect 3157 13685 3191 13719
rect 50537 13685 50571 13719
rect 56149 13685 56183 13719
rect 49709 13481 49743 13515
rect 55321 13481 55355 13515
rect 51917 13413 51951 13447
rect 52653 13413 52687 13447
rect 53941 13413 53975 13447
rect 54677 13413 54711 13447
rect 1685 13345 1719 13379
rect 2973 13345 3007 13379
rect 5089 13345 5123 13379
rect 47869 13345 47903 13379
rect 49893 13345 49927 13379
rect 50353 13345 50387 13379
rect 50537 13345 50571 13379
rect 51641 13345 51675 13379
rect 52837 13345 52871 13379
rect 53849 13345 53883 13379
rect 54585 13345 54619 13379
rect 55229 13345 55263 13379
rect 55413 13345 55447 13379
rect 57253 13345 57287 13379
rect 1869 13277 1903 13311
rect 50445 13277 50479 13311
rect 51457 13277 51491 13311
rect 52009 13277 52043 13311
rect 53113 13277 53147 13311
rect 57069 13277 57103 13311
rect 2053 13209 2087 13243
rect 51733 13209 51767 13243
rect 5089 13141 5123 13175
rect 48145 13141 48179 13175
rect 53021 13141 53055 13175
rect 57437 13141 57471 13175
rect 2973 12937 3007 12971
rect 57345 12937 57379 12971
rect 49801 12801 49835 12835
rect 55045 12801 55079 12835
rect 2881 12733 2915 12767
rect 49341 12733 49375 12767
rect 50068 12733 50102 12767
rect 51641 12733 51675 12767
rect 52745 12733 52779 12767
rect 52837 12733 52871 12767
rect 53021 12733 53055 12767
rect 53113 12733 53147 12767
rect 54033 12733 54067 12767
rect 54217 12733 54251 12767
rect 57253 12733 57287 12767
rect 1869 12665 1903 12699
rect 55312 12665 55346 12699
rect 57989 12665 58023 12699
rect 1961 12597 1995 12631
rect 51181 12597 51215 12631
rect 51733 12597 51767 12631
rect 52561 12597 52595 12631
rect 54125 12597 54159 12631
rect 56425 12597 56459 12631
rect 58081 12597 58115 12631
rect 51457 12393 51491 12427
rect 55597 12393 55631 12427
rect 58173 12393 58207 12427
rect 50445 12325 50479 12359
rect 52561 12325 52595 12359
rect 53910 12325 53944 12359
rect 1593 12257 1627 12291
rect 2697 12257 2731 12291
rect 49893 12257 49927 12291
rect 50353 12257 50387 12291
rect 50537 12257 50571 12291
rect 51641 12257 51675 12291
rect 51733 12257 51767 12291
rect 52009 12257 52043 12291
rect 52791 12257 52825 12291
rect 52929 12257 52963 12291
rect 53021 12257 53055 12291
rect 53205 12257 53239 12291
rect 53665 12257 53699 12291
rect 55505 12257 55539 12291
rect 56701 12257 56735 12291
rect 57529 12257 57563 12291
rect 1777 12189 1811 12223
rect 4445 12189 4479 12223
rect 51917 12189 51951 12223
rect 57713 12189 57747 12223
rect 1961 12121 1995 12155
rect 49709 12121 49743 12155
rect 55045 12121 55079 12155
rect 2881 12053 2915 12087
rect 56793 12053 56827 12087
rect 3249 11849 3283 11883
rect 51273 11849 51307 11883
rect 51825 11849 51859 11883
rect 55045 11849 55079 11883
rect 55597 11849 55631 11883
rect 54585 11781 54619 11815
rect 56701 11781 56735 11815
rect 52745 11713 52779 11747
rect 57345 11713 57379 11747
rect 3433 11645 3467 11679
rect 4077 11645 4111 11679
rect 49249 11645 49283 11679
rect 49433 11645 49467 11679
rect 49893 11645 49927 11679
rect 51733 11645 51767 11679
rect 52377 11645 52411 11679
rect 52549 11645 52583 11679
rect 52653 11645 52687 11679
rect 52929 11645 52963 11679
rect 54769 11645 54803 11679
rect 54861 11645 54895 11679
rect 55137 11645 55171 11679
rect 55597 11645 55631 11679
rect 55781 11645 55815 11679
rect 56517 11645 56551 11679
rect 57161 11645 57195 11679
rect 1869 11577 1903 11611
rect 2605 11577 2639 11611
rect 2789 11577 2823 11611
rect 49341 11577 49375 11611
rect 50160 11577 50194 11611
rect 1961 11509 1995 11543
rect 53113 11509 53147 11543
rect 57805 11509 57839 11543
rect 2513 11305 2547 11339
rect 50445 11305 50479 11339
rect 51549 11305 51583 11339
rect 52653 11305 52687 11339
rect 54677 11237 54711 11271
rect 57989 11237 58023 11271
rect 58173 11237 58207 11271
rect 1869 11169 1903 11203
rect 3157 11169 3191 11203
rect 49065 11169 49099 11203
rect 49893 11169 49927 11203
rect 50353 11169 50387 11203
rect 50537 11169 50571 11203
rect 51457 11169 51491 11203
rect 51641 11169 51675 11203
rect 52887 11169 52921 11203
rect 53021 11169 53055 11203
rect 53113 11169 53147 11203
rect 53389 11169 53423 11203
rect 54033 11169 54067 11203
rect 54125 11169 54159 11203
rect 54309 11169 54343 11203
rect 54585 11169 54619 11203
rect 55321 11169 55355 11203
rect 55505 11169 55539 11203
rect 55689 11169 55723 11203
rect 56701 11169 56735 11203
rect 56885 11169 56919 11203
rect 2053 11101 2087 11135
rect 53205 11101 53239 11135
rect 2973 11033 3007 11067
rect 55321 11033 55355 11067
rect 56701 10965 56735 10999
rect 2053 10761 2087 10795
rect 55045 10761 55079 10795
rect 52193 10693 52227 10727
rect 50169 10625 50203 10659
rect 1685 10557 1719 10591
rect 1869 10557 1903 10591
rect 50813 10557 50847 10591
rect 51457 10557 51491 10591
rect 52009 10557 52043 10591
rect 52929 10557 52963 10591
rect 54493 10557 54527 10591
rect 54861 10557 54895 10591
rect 55505 10557 55539 10591
rect 55772 10557 55806 10591
rect 54677 10489 54711 10523
rect 54769 10489 54803 10523
rect 57989 10489 58023 10523
rect 58173 10489 58207 10523
rect 51273 10421 51307 10455
rect 53021 10421 53055 10455
rect 56885 10421 56919 10455
rect 2513 10217 2547 10251
rect 56701 10217 56735 10251
rect 58173 10217 58207 10251
rect 50169 10149 50203 10183
rect 1869 10081 1903 10115
rect 2697 10081 2731 10115
rect 3341 10081 3375 10115
rect 49341 10081 49375 10115
rect 49985 10081 50019 10115
rect 51713 10081 51747 10115
rect 53527 10081 53561 10115
rect 53665 10081 53699 10115
rect 53757 10081 53791 10115
rect 53941 10081 53975 10115
rect 54585 10081 54619 10115
rect 55229 10081 55263 10115
rect 55367 10081 55401 10115
rect 55505 10081 55539 10115
rect 55643 10081 55677 10115
rect 56885 10081 56919 10115
rect 57713 10081 57747 10115
rect 51457 10013 51491 10047
rect 54677 10013 54711 10047
rect 56701 10013 56735 10047
rect 57529 10013 57563 10047
rect 52837 9945 52871 9979
rect 57069 9945 57103 9979
rect 1961 9877 1995 9911
rect 50353 9877 50387 9911
rect 53297 9877 53331 9911
rect 55781 9877 55815 9911
rect 2145 9673 2179 9707
rect 51181 9673 51215 9707
rect 57161 9673 57195 9707
rect 2881 9605 2915 9639
rect 1961 9537 1995 9571
rect 3709 9537 3743 9571
rect 56793 9537 56827 9571
rect 1777 9469 1811 9503
rect 3065 9469 3099 9503
rect 49065 9469 49099 9503
rect 49332 9469 49366 9503
rect 51181 9469 51215 9503
rect 51365 9469 51399 9503
rect 52098 9469 52132 9503
rect 52469 9469 52503 9503
rect 52561 9469 52595 9503
rect 53389 9469 53423 9503
rect 54033 9469 54067 9503
rect 54289 9469 54323 9503
rect 55873 9469 55907 9503
rect 56977 9469 57011 9503
rect 57989 9401 58023 9435
rect 58173 9401 58207 9435
rect 50445 9333 50479 9367
rect 51917 9333 51951 9367
rect 52101 9333 52135 9367
rect 53389 9333 53423 9367
rect 55413 9333 55447 9367
rect 55965 9333 55999 9367
rect 49985 9129 50019 9163
rect 52377 9129 52411 9163
rect 53297 9129 53331 9163
rect 54493 9129 54527 9163
rect 56885 9129 56919 9163
rect 58173 9129 58207 9163
rect 51549 9061 51583 9095
rect 52929 9061 52963 9095
rect 53113 9061 53147 9095
rect 2973 8993 3007 9027
rect 48053 8993 48087 9027
rect 48697 8993 48731 9027
rect 48881 8993 48915 9027
rect 49525 8993 49559 9027
rect 50169 8993 50203 9027
rect 50261 8993 50295 9027
rect 50537 8993 50571 9027
rect 52285 8993 52319 9027
rect 53757 8993 53791 9027
rect 53941 8993 53975 9027
rect 54677 8993 54711 9027
rect 54769 8993 54803 9027
rect 55045 8993 55079 9027
rect 55505 8993 55539 9027
rect 57069 8993 57103 9027
rect 57529 8993 57563 9027
rect 1685 8925 1719 8959
rect 1869 8925 1903 8959
rect 50445 8925 50479 8959
rect 52193 8925 52227 8959
rect 55597 8925 55631 8959
rect 57713 8925 57747 8959
rect 2789 8857 2823 8891
rect 49341 8857 49375 8891
rect 2329 8789 2363 8823
rect 48697 8789 48731 8823
rect 51641 8789 51675 8823
rect 52193 8789 52227 8823
rect 53757 8789 53791 8823
rect 54953 8789 54987 8823
rect 4353 8585 4387 8619
rect 47685 8585 47719 8619
rect 2789 8517 2823 8551
rect 3617 8517 3651 8551
rect 50261 8517 50295 8551
rect 51457 8517 51491 8551
rect 53021 8517 53055 8551
rect 55413 8517 55447 8551
rect 48881 8449 48915 8483
rect 53113 8449 53147 8483
rect 56425 8449 56459 8483
rect 2605 8381 2639 8415
rect 3157 8381 3191 8415
rect 3341 8381 3375 8415
rect 47041 8381 47075 8415
rect 47685 8381 47719 8415
rect 47869 8381 47903 8415
rect 50721 8381 50755 8415
rect 51365 8381 51399 8415
rect 52009 8381 52043 8415
rect 52193 8381 52227 8415
rect 52837 8381 52871 8415
rect 52929 8381 52963 8415
rect 54033 8381 54067 8415
rect 54289 8381 54323 8415
rect 56609 8381 56643 8415
rect 1869 8313 1903 8347
rect 2053 8313 2087 8347
rect 49148 8313 49182 8347
rect 57069 8313 57103 8347
rect 57989 8313 58023 8347
rect 58173 8313 58207 8347
rect 50813 8245 50847 8279
rect 52101 8245 52135 8279
rect 49341 8041 49375 8075
rect 50077 8041 50111 8075
rect 56701 8041 56735 8075
rect 51908 7973 51942 8007
rect 1869 7905 1903 7939
rect 2513 7905 2547 7939
rect 3341 7905 3375 7939
rect 46949 7905 46983 7939
rect 47409 7905 47443 7939
rect 47593 7905 47627 7939
rect 48053 7905 48087 7939
rect 48881 7905 48915 7939
rect 49525 7905 49559 7939
rect 49985 7905 50019 7939
rect 50169 7905 50203 7939
rect 51641 7905 51675 7939
rect 53573 7905 53607 7939
rect 53733 7905 53767 7939
rect 54677 7905 54711 7939
rect 55137 7905 55171 7939
rect 55229 7905 55263 7939
rect 56885 7905 56919 7939
rect 47501 7837 47535 7871
rect 53481 7837 53515 7871
rect 48697 7769 48731 7803
rect 54401 7837 54435 7871
rect 57345 7837 57379 7871
rect 57529 7837 57563 7871
rect 1961 7701 1995 7735
rect 2697 7701 2731 7735
rect 3157 7701 3191 7735
rect 48237 7701 48271 7735
rect 53021 7701 53055 7735
rect 53481 7701 53515 7735
rect 53573 7701 53607 7735
rect 54401 7701 54435 7735
rect 54493 7701 54527 7735
rect 57713 7701 57747 7735
rect 2053 7497 2087 7531
rect 50721 7497 50755 7531
rect 51457 7497 51491 7531
rect 55781 7497 55815 7531
rect 49801 7429 49835 7463
rect 51733 7429 51767 7463
rect 52745 7429 52779 7463
rect 1685 7361 1719 7395
rect 2973 7361 3007 7395
rect 49893 7361 49927 7395
rect 50353 7361 50387 7395
rect 51457 7361 51491 7395
rect 54125 7361 54159 7395
rect 56425 7361 56459 7395
rect 58173 7361 58207 7395
rect 1869 7293 1903 7327
rect 46581 7293 46615 7327
rect 46949 7293 46983 7327
rect 47225 7293 47259 7327
rect 47869 7293 47903 7327
rect 48973 7293 49007 7327
rect 49617 7293 49651 7327
rect 51365 7293 51399 7327
rect 52561 7293 52595 7327
rect 52837 7293 52871 7327
rect 54033 7293 54067 7327
rect 54677 7293 54711 7327
rect 54861 7293 54895 7327
rect 55965 7293 55999 7327
rect 56609 7293 56643 7327
rect 57989 7225 58023 7259
rect 48789 7157 48823 7191
rect 49433 7157 49467 7191
rect 50721 7157 50755 7191
rect 50905 7157 50939 7191
rect 52377 7157 52411 7191
rect 54769 7157 54803 7191
rect 57069 7157 57103 7191
rect 2329 6953 2363 6987
rect 52101 6953 52135 6987
rect 53389 6953 53423 6987
rect 58173 6953 58207 6987
rect 54484 6885 54518 6919
rect 56885 6885 56919 6919
rect 1685 6817 1719 6851
rect 2973 6817 3007 6851
rect 45109 6817 45143 6851
rect 47593 6817 47627 6851
rect 48964 6817 48998 6851
rect 51825 6817 51859 6851
rect 53205 6817 53239 6851
rect 53389 6817 53423 6851
rect 57713 6817 57747 6851
rect 1869 6749 1903 6783
rect 48697 6749 48731 6783
rect 51641 6749 51675 6783
rect 52193 6749 52227 6783
rect 53757 6749 53791 6783
rect 54217 6749 54251 6783
rect 57069 6749 57103 6783
rect 57529 6749 57563 6783
rect 46949 6681 46983 6715
rect 51917 6681 51951 6715
rect 48237 6613 48271 6647
rect 50077 6613 50111 6647
rect 55597 6613 55631 6647
rect 2513 6409 2547 6443
rect 46581 6409 46615 6443
rect 52377 6409 52411 6443
rect 47777 6273 47811 6307
rect 52745 6273 52779 6307
rect 54401 6273 54435 6307
rect 54493 6273 54527 6307
rect 55321 6273 55355 6307
rect 57529 6273 57563 6307
rect 2697 6205 2731 6239
rect 3341 6205 3375 6239
rect 44465 6205 44499 6239
rect 45017 6205 45051 6239
rect 45293 6205 45327 6239
rect 45661 6205 45695 6239
rect 45937 6205 45971 6239
rect 47225 6205 47259 6239
rect 47685 6205 47719 6239
rect 47869 6205 47903 6239
rect 49065 6205 49099 6239
rect 49525 6205 49559 6239
rect 50169 6205 50203 6239
rect 50445 6205 50479 6239
rect 50537 6205 50571 6239
rect 51181 6205 51215 6239
rect 51365 6205 51399 6239
rect 51641 6205 51675 6239
rect 52561 6205 52595 6239
rect 52653 6205 52687 6239
rect 52837 6205 52871 6239
rect 54217 6205 54251 6239
rect 54309 6205 54343 6239
rect 54677 6205 54711 6239
rect 55229 6205 55263 6239
rect 56425 6205 56459 6239
rect 56609 6205 56643 6239
rect 57713 6205 57747 6239
rect 1869 6137 1903 6171
rect 50353 6137 50387 6171
rect 51733 6137 51767 6171
rect 1961 6069 1995 6103
rect 48881 6069 48915 6103
rect 49709 6069 49743 6103
rect 50721 6069 50755 6103
rect 54033 6069 54067 6103
rect 57069 6069 57103 6103
rect 58173 6069 58207 6103
rect 2329 5865 2363 5899
rect 52745 5865 52779 5899
rect 47685 5797 47719 5831
rect 50261 5797 50295 5831
rect 57989 5797 58023 5831
rect 1685 5729 1719 5763
rect 2973 5729 3007 5763
rect 43821 5729 43855 5763
rect 46489 5729 46523 5763
rect 47593 5729 47627 5763
rect 47777 5729 47811 5763
rect 48421 5729 48455 5763
rect 49065 5729 49099 5763
rect 49709 5729 49743 5763
rect 50169 5729 50203 5763
rect 51779 5729 51813 5763
rect 51898 5729 51932 5763
rect 51998 5729 52032 5763
rect 52193 5729 52227 5763
rect 52929 5729 52963 5763
rect 53021 5729 53055 5763
rect 53297 5729 53331 5763
rect 53757 5729 53791 5763
rect 53849 5729 53883 5763
rect 54493 5729 54527 5763
rect 55597 5729 55631 5763
rect 58173 5729 58207 5763
rect 1869 5661 1903 5695
rect 4445 5661 4479 5695
rect 56701 5661 56735 5695
rect 56885 5661 56919 5695
rect 2789 5593 2823 5627
rect 49525 5593 49559 5627
rect 44373 5525 44407 5559
rect 44649 5525 44683 5559
rect 44925 5525 44959 5559
rect 45293 5525 45327 5559
rect 47133 5525 47167 5559
rect 48237 5525 48271 5559
rect 48881 5525 48915 5559
rect 51549 5525 51583 5559
rect 53205 5525 53239 5559
rect 54585 5525 54619 5559
rect 55689 5525 55723 5559
rect 57069 5525 57103 5559
rect 47685 5321 47719 5355
rect 50721 5321 50755 5355
rect 51273 5321 51307 5355
rect 52009 5321 52043 5355
rect 53021 5321 53055 5355
rect 56977 5321 57011 5355
rect 55781 5253 55815 5287
rect 57897 5253 57931 5287
rect 2053 5185 2087 5219
rect 4077 5185 4111 5219
rect 44373 5185 44407 5219
rect 57713 5185 57747 5219
rect 2789 5117 2823 5151
rect 3433 5117 3467 5151
rect 43545 5117 43579 5151
rect 45017 5117 45051 5151
rect 45661 5117 45695 5151
rect 46581 5117 46615 5151
rect 47041 5117 47075 5151
rect 47225 5117 47259 5151
rect 47869 5117 47903 5151
rect 49341 5117 49375 5151
rect 51181 5117 51215 5151
rect 51917 5117 51951 5151
rect 52101 5117 52135 5151
rect 52929 5117 52963 5151
rect 54039 5117 54073 5151
rect 54217 5117 54251 5151
rect 55413 5117 55447 5151
rect 55597 5117 55631 5151
rect 56885 5117 56919 5151
rect 57529 5117 57563 5151
rect 1869 5049 1903 5083
rect 2605 5049 2639 5083
rect 47133 5049 47167 5083
rect 49608 5049 49642 5083
rect 54769 5049 54803 5083
rect 3249 4981 3283 5015
rect 54125 4981 54159 5015
rect 54861 4981 54895 5015
rect 57345 4981 57379 5015
rect 2605 4777 2639 4811
rect 48789 4777 48823 4811
rect 49985 4777 50019 4811
rect 51794 4709 51828 4743
rect 53656 4709 53690 4743
rect 56885 4709 56919 4743
rect 2145 4641 2179 4675
rect 3249 4641 3283 4675
rect 38117 4641 38151 4675
rect 46857 4641 46891 4675
rect 47501 4641 47535 4675
rect 48145 4641 48179 4675
rect 48605 4641 48639 4675
rect 49433 4641 49467 4675
rect 49893 4641 49927 4675
rect 50077 4641 50111 4675
rect 55321 4641 55355 4675
rect 1961 4573 1995 4607
rect 51549 4573 51583 4607
rect 53389 4573 53423 4607
rect 57345 4573 57379 4607
rect 57529 4573 57563 4607
rect 57713 4573 57747 4607
rect 46673 4505 46707 4539
rect 52929 4505 52963 4539
rect 55505 4505 55539 4539
rect 3065 4437 3099 4471
rect 4445 4437 4479 4471
rect 34529 4437 34563 4471
rect 35909 4437 35943 4471
rect 36737 4437 36771 4471
rect 37933 4437 37967 4471
rect 38761 4437 38795 4471
rect 42809 4437 42843 4471
rect 43545 4437 43579 4471
rect 44189 4437 44223 4471
rect 45109 4437 45143 4471
rect 47317 4437 47351 4471
rect 47961 4437 47995 4471
rect 49249 4437 49283 4471
rect 54769 4437 54803 4471
rect 56977 4437 57011 4471
rect 57989 4437 58023 4471
rect 2881 4233 2915 4267
rect 52193 4233 52227 4267
rect 56885 4233 56919 4267
rect 39773 4165 39807 4199
rect 41153 4165 41187 4199
rect 41981 4165 42015 4199
rect 46581 4165 46615 4199
rect 47041 4165 47075 4199
rect 1777 4097 1811 4131
rect 56333 4097 56367 4131
rect 56517 4097 56551 4131
rect 56701 4097 56735 4131
rect 1593 4029 1627 4063
rect 3617 4029 3651 4063
rect 4261 4029 4295 4063
rect 4721 4029 4755 4063
rect 33333 4029 33367 4063
rect 33977 4029 34011 4063
rect 34621 4029 34655 4063
rect 35725 4029 35759 4063
rect 36369 4029 36403 4063
rect 36829 4029 36863 4063
rect 38485 4029 38519 4063
rect 39129 4029 39163 4063
rect 40509 4029 40543 4063
rect 42625 4029 42659 4063
rect 44189 4029 44223 4063
rect 45293 4029 45327 4063
rect 45937 4029 45971 4063
rect 46397 4029 46431 4063
rect 47225 4029 47259 4063
rect 47869 4029 47903 4063
rect 49157 4029 49191 4063
rect 49801 4029 49835 4063
rect 50445 4029 50479 4063
rect 50905 4029 50939 4063
rect 51733 4029 51767 4063
rect 52377 4029 52411 4063
rect 52929 4029 52963 4063
rect 55873 4029 55907 4063
rect 57989 4029 58023 4063
rect 2237 3961 2271 3995
rect 2789 3961 2823 3995
rect 53113 3961 53147 3995
rect 54401 3961 54435 3995
rect 55137 3961 55171 3995
rect 56057 3961 56091 3995
rect 58173 3961 58207 3995
rect 3433 3893 3467 3927
rect 33149 3893 33183 3927
rect 34437 3893 34471 3927
rect 35541 3893 35575 3927
rect 36185 3893 36219 3927
rect 37013 3893 37047 3927
rect 38301 3893 38335 3927
rect 42441 3893 42475 3927
rect 44005 3893 44039 3927
rect 45109 3893 45143 3927
rect 45753 3893 45787 3927
rect 47685 3893 47719 3927
rect 48973 3893 49007 3927
rect 49617 3893 49651 3927
rect 50261 3893 50295 3927
rect 51089 3893 51123 3927
rect 51549 3893 51583 3927
rect 54493 3893 54527 3927
rect 55229 3893 55263 3927
rect 44465 3689 44499 3723
rect 50537 3621 50571 3655
rect 55597 3621 55631 3655
rect 56885 3621 56919 3655
rect 1961 3553 1995 3587
rect 3157 3553 3191 3587
rect 5549 3553 5583 3587
rect 6193 3553 6227 3587
rect 28549 3553 28583 3587
rect 29377 3553 29411 3587
rect 30757 3553 30791 3587
rect 33333 3553 33367 3587
rect 34253 3553 34287 3587
rect 35817 3553 35851 3587
rect 37105 3553 37139 3587
rect 38025 3553 38059 3587
rect 38945 3553 38979 3587
rect 39773 3553 39807 3587
rect 41153 3553 41187 3587
rect 42165 3553 42199 3587
rect 42717 3553 42751 3587
rect 43353 3553 43387 3587
rect 44649 3553 44683 3587
rect 45293 3553 45327 3587
rect 46305 3553 46339 3587
rect 47041 3553 47075 3587
rect 47777 3553 47811 3587
rect 48513 3553 48547 3587
rect 49801 3553 49835 3587
rect 50353 3553 50387 3587
rect 52101 3553 52135 3587
rect 53021 3553 53055 3587
rect 53941 3553 53975 3587
rect 55045 3553 55079 3587
rect 57713 3553 57747 3587
rect 2145 3485 2179 3519
rect 53757 3485 53791 3519
rect 57345 3485 57379 3519
rect 57529 3485 57563 3519
rect 2329 3417 2363 3451
rect 43545 3417 43579 3451
rect 45109 3417 45143 3451
rect 55781 3417 55815 3451
rect 3249 3349 3283 3383
rect 4445 3349 4479 3383
rect 5089 3349 5123 3383
rect 30573 3349 30607 3383
rect 31401 3349 31435 3383
rect 32045 3349 32079 3383
rect 32781 3349 32815 3383
rect 33425 3349 33459 3383
rect 34345 3349 34379 3383
rect 35909 3349 35943 3383
rect 37197 3349 37231 3383
rect 38117 3349 38151 3383
rect 39037 3349 39071 3383
rect 39589 3349 39623 3383
rect 40969 3349 41003 3383
rect 41981 3349 42015 3383
rect 42809 3349 42843 3383
rect 46397 3349 46431 3383
rect 47133 3349 47167 3383
rect 47869 3349 47903 3383
rect 48605 3349 48639 3383
rect 49617 3349 49651 3383
rect 52193 3349 52227 3383
rect 53113 3349 53147 3383
rect 54401 3349 54435 3383
rect 54861 3349 54895 3383
rect 56977 3349 57011 3383
rect 57989 3349 58023 3383
rect 3157 3145 3191 3179
rect 4629 3145 4663 3179
rect 34253 3145 34287 3179
rect 37381 3145 37415 3179
rect 38669 3145 38703 3179
rect 46213 3145 46247 3179
rect 47869 3145 47903 3179
rect 53021 3145 53055 3179
rect 55965 3145 55999 3179
rect 57989 3145 58023 3179
rect 6285 3077 6319 3111
rect 29285 3077 29319 3111
rect 57253 3077 57287 3111
rect 1685 3009 1719 3043
rect 2789 3009 2823 3043
rect 2973 3009 3007 3043
rect 28825 3009 28859 3043
rect 29929 3009 29963 3043
rect 30113 3009 30147 3043
rect 33701 3009 33735 3043
rect 35541 3009 35575 3043
rect 38485 3009 38519 3043
rect 40049 3009 40083 3043
rect 43729 3009 43763 3043
rect 44189 3009 44223 3043
rect 45569 3009 45603 3043
rect 45753 3009 45787 3043
rect 47225 3009 47259 3043
rect 47409 3009 47443 3043
rect 48789 3009 48823 3043
rect 48973 3009 49007 3043
rect 52561 3009 52595 3043
rect 55597 3009 55631 3043
rect 56885 3009 56919 3043
rect 57069 3009 57103 3043
rect 1409 2941 1443 2975
rect 4813 2941 4847 2975
rect 5457 2941 5491 2975
rect 6285 2941 6319 2975
rect 6837 2941 6871 2975
rect 7481 2941 7515 2975
rect 8861 2941 8895 2975
rect 29469 2941 29503 2975
rect 31309 2941 31343 2975
rect 33241 2941 33275 2975
rect 33885 2941 33919 2975
rect 35357 2941 35391 2975
rect 37197 2941 37231 2975
rect 38301 2941 38335 2975
rect 39589 2941 39623 2975
rect 40233 2941 40267 2975
rect 43545 2941 43579 2975
rect 52377 2941 52411 2975
rect 54861 2941 54895 2975
rect 55781 2941 55815 2975
rect 58173 2941 58207 2975
rect 3985 2873 4019 2907
rect 4169 2873 4203 2907
rect 31953 2873 31987 2907
rect 32137 2873 32171 2907
rect 36001 2873 36035 2907
rect 36553 2873 36587 2907
rect 40693 2873 40727 2907
rect 41245 2873 41279 2907
rect 41981 2873 42015 2907
rect 44741 2873 44775 2907
rect 49433 2873 49467 2907
rect 49985 2873 50019 2907
rect 50721 2873 50755 2907
rect 51457 2873 51491 2907
rect 54125 2873 54159 2907
rect 5273 2805 5307 2839
rect 30573 2805 30607 2839
rect 31125 2805 31159 2839
rect 33057 2805 33091 2839
rect 36645 2805 36679 2839
rect 39405 2805 39439 2839
rect 41337 2805 41371 2839
rect 42073 2805 42107 2839
rect 44833 2805 44867 2839
rect 50077 2805 50111 2839
rect 50813 2805 50847 2839
rect 51549 2805 51583 2839
rect 54217 2805 54251 2839
rect 54953 2805 54987 2839
rect 2329 2601 2363 2635
rect 35357 2601 35391 2635
rect 36921 2601 36955 2635
rect 39589 2601 39623 2635
rect 44925 2601 44959 2635
rect 46029 2601 46063 2635
rect 47593 2601 47627 2635
rect 50261 2601 50295 2635
rect 51365 2601 51399 2635
rect 54033 2601 54067 2635
rect 55597 2601 55631 2635
rect 56701 2601 56735 2635
rect 2881 2533 2915 2567
rect 4905 2533 4939 2567
rect 29837 2533 29871 2567
rect 37841 2533 37875 2567
rect 40693 2533 40727 2567
rect 48145 2533 48179 2567
rect 57989 2533 58023 2567
rect 1685 2465 1719 2499
rect 4261 2465 4295 2499
rect 5549 2465 5583 2499
rect 6929 2465 6963 2499
rect 7573 2465 7607 2499
rect 8217 2465 8251 2499
rect 9781 2465 9815 2499
rect 10793 2465 10827 2499
rect 12265 2465 12299 2499
rect 12909 2465 12943 2499
rect 13553 2465 13587 2499
rect 14933 2465 14967 2499
rect 15577 2465 15611 2499
rect 16405 2465 16439 2499
rect 17601 2465 17635 2499
rect 18245 2465 18279 2499
rect 19165 2465 19199 2499
rect 20269 2465 20303 2499
rect 21097 2465 21131 2499
rect 21833 2465 21867 2499
rect 22937 2465 22971 2499
rect 23857 2465 23891 2499
rect 25605 2465 25639 2499
rect 26249 2465 26283 2499
rect 26893 2465 26927 2499
rect 28273 2465 28307 2499
rect 29101 2465 29135 2499
rect 30941 2465 30975 2499
rect 32045 2465 32079 2499
rect 32229 2465 32263 2499
rect 33609 2465 33643 2499
rect 33793 2465 33827 2499
rect 34713 2465 34747 2499
rect 34897 2465 34931 2499
rect 36461 2465 36495 2499
rect 38945 2465 38979 2499
rect 39129 2465 39163 2499
rect 40049 2465 40083 2499
rect 40233 2465 40267 2499
rect 41613 2465 41647 2499
rect 41797 2465 41831 2499
rect 42717 2465 42751 2499
rect 42901 2465 42935 2499
rect 44281 2465 44315 2499
rect 44465 2465 44499 2499
rect 45385 2465 45419 2499
rect 45569 2465 45603 2499
rect 46949 2465 46983 2499
rect 47133 2465 47167 2499
rect 49617 2465 49651 2499
rect 49801 2465 49835 2499
rect 52285 2465 52319 2499
rect 53389 2465 53423 2499
rect 53573 2465 53607 2499
rect 56057 2465 56091 2499
rect 1869 2397 1903 2431
rect 4445 2397 4479 2431
rect 31125 2397 31159 2431
rect 36277 2397 36311 2431
rect 50721 2397 50755 2431
rect 50905 2397 50939 2431
rect 52469 2397 52503 2431
rect 54953 2397 54987 2431
rect 55137 2397 55171 2431
rect 56241 2397 56275 2431
rect 5365 2329 5399 2363
rect 30021 2329 30055 2363
rect 31309 2329 31343 2363
rect 32413 2329 32447 2363
rect 33977 2329 34011 2363
rect 38025 2329 38059 2363
rect 41981 2329 42015 2363
rect 43085 2329 43119 2363
rect 48329 2329 48363 2363
rect 52653 2329 52687 2363
rect 2973 2261 3007 2295
rect 29193 2261 29227 2295
rect 54769 2261 54803 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 55214 58284 55220 58336
rect 55272 58324 55278 58336
rect 56410 58324 56416 58336
rect 55272 58296 56416 58324
rect 55272 58284 55278 58296
rect 56410 58284 56416 58296
rect 56468 58284 56474 58336
rect 1104 57690 58880 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 58880 57690
rect 1104 57616 58880 57638
rect 53929 57579 53987 57585
rect 53929 57545 53941 57579
rect 53975 57576 53987 57579
rect 59538 57576 59544 57588
rect 53975 57548 59544 57576
rect 53975 57545 53987 57548
rect 53929 57539 53987 57545
rect 59538 57536 59544 57548
rect 59596 57536 59602 57588
rect 4525 57511 4583 57517
rect 4525 57477 4537 57511
rect 4571 57508 4583 57511
rect 4614 57508 4620 57520
rect 4571 57480 4620 57508
rect 4571 57477 4583 57480
rect 4525 57471 4583 57477
rect 4614 57468 4620 57480
rect 4672 57468 4678 57520
rect 24026 57468 24032 57520
rect 24084 57508 24090 57520
rect 24084 57480 25636 57508
rect 24084 57468 24090 57480
rect 6638 57400 6644 57452
rect 6696 57440 6702 57452
rect 6696 57412 6960 57440
rect 6696 57400 6702 57412
rect 1394 57372 1400 57384
rect 1355 57344 1400 57372
rect 1394 57332 1400 57344
rect 1452 57332 1458 57384
rect 2038 57372 2044 57384
rect 1999 57344 2044 57372
rect 2038 57332 2044 57344
rect 2096 57332 2102 57384
rect 2685 57375 2743 57381
rect 2685 57341 2697 57375
rect 2731 57372 2743 57375
rect 2774 57372 2780 57384
rect 2731 57344 2780 57372
rect 2731 57341 2743 57344
rect 2685 57335 2743 57341
rect 2774 57332 2780 57344
rect 2832 57332 2838 57384
rect 5074 57372 5080 57384
rect 5035 57344 5080 57372
rect 5074 57332 5080 57344
rect 5132 57332 5138 57384
rect 5813 57375 5871 57381
rect 5813 57341 5825 57375
rect 5859 57372 5871 57375
rect 5902 57372 5908 57384
rect 5859 57344 5908 57372
rect 5859 57341 5871 57344
rect 5813 57335 5871 57341
rect 5902 57332 5908 57344
rect 5960 57332 5966 57384
rect 6932 57381 6960 57412
rect 14550 57400 14556 57452
rect 14608 57440 14614 57452
rect 14608 57412 15240 57440
rect 14608 57400 14614 57412
rect 6917 57375 6975 57381
rect 6917 57341 6929 57375
rect 6963 57341 6975 57375
rect 6917 57335 6975 57341
rect 7466 57332 7472 57384
rect 7524 57372 7530 57384
rect 7561 57375 7619 57381
rect 7561 57372 7573 57375
rect 7524 57344 7573 57372
rect 7524 57332 7530 57344
rect 7561 57341 7573 57344
rect 7607 57341 7619 57375
rect 8202 57372 8208 57384
rect 8163 57344 8208 57372
rect 7561 57335 7619 57341
rect 8202 57332 8208 57344
rect 8260 57332 8266 57384
rect 9030 57332 9036 57384
rect 9088 57372 9094 57384
rect 9585 57375 9643 57381
rect 9585 57372 9597 57375
rect 9088 57344 9597 57372
rect 9088 57332 9094 57344
rect 9585 57341 9597 57344
rect 9631 57341 9643 57375
rect 9585 57335 9643 57341
rect 9766 57332 9772 57384
rect 9824 57372 9830 57384
rect 10229 57375 10287 57381
rect 10229 57372 10241 57375
rect 9824 57344 10241 57372
rect 9824 57332 9830 57344
rect 10229 57341 10241 57344
rect 10275 57341 10287 57375
rect 10229 57335 10287 57341
rect 10594 57332 10600 57384
rect 10652 57372 10658 57384
rect 10873 57375 10931 57381
rect 10873 57372 10885 57375
rect 10652 57344 10885 57372
rect 10652 57332 10658 57344
rect 10873 57341 10885 57344
rect 10919 57341 10931 57375
rect 10873 57335 10931 57341
rect 11422 57332 11428 57384
rect 11480 57372 11486 57384
rect 12253 57375 12311 57381
rect 12253 57372 12265 57375
rect 11480 57344 12265 57372
rect 11480 57332 11486 57344
rect 12253 57341 12265 57344
rect 12299 57341 12311 57375
rect 12253 57335 12311 57341
rect 12434 57332 12440 57384
rect 12492 57372 12498 57384
rect 12897 57375 12955 57381
rect 12897 57372 12909 57375
rect 12492 57344 12909 57372
rect 12492 57332 12498 57344
rect 12897 57341 12909 57344
rect 12943 57341 12955 57375
rect 12897 57335 12955 57341
rect 12986 57332 12992 57384
rect 13044 57372 13050 57384
rect 13541 57375 13599 57381
rect 13541 57372 13553 57375
rect 13044 57344 13553 57372
rect 13044 57332 13050 57344
rect 13541 57341 13553 57344
rect 13587 57341 13599 57375
rect 13541 57335 13599 57341
rect 13814 57332 13820 57384
rect 13872 57372 13878 57384
rect 14921 57375 14979 57381
rect 14921 57372 14933 57375
rect 13872 57344 14933 57372
rect 13872 57332 13878 57344
rect 14921 57341 14933 57344
rect 14967 57341 14979 57375
rect 15212 57372 15240 57412
rect 15378 57400 15384 57452
rect 15436 57440 15442 57452
rect 15436 57412 16252 57440
rect 15436 57400 15442 57412
rect 16224 57381 16252 57412
rect 20070 57400 20076 57452
rect 20128 57440 20134 57452
rect 20128 57412 20944 57440
rect 20128 57400 20134 57412
rect 15565 57375 15623 57381
rect 15565 57372 15577 57375
rect 15212 57344 15577 57372
rect 14921 57335 14979 57341
rect 15565 57341 15577 57344
rect 15611 57341 15623 57375
rect 15565 57335 15623 57341
rect 16209 57375 16267 57381
rect 16209 57341 16221 57375
rect 16255 57341 16267 57375
rect 16209 57335 16267 57341
rect 16942 57332 16948 57384
rect 17000 57372 17006 57384
rect 17589 57375 17647 57381
rect 17589 57372 17601 57375
rect 17000 57344 17601 57372
rect 17000 57332 17006 57344
rect 17589 57341 17601 57344
rect 17635 57341 17647 57375
rect 17589 57335 17647 57341
rect 17678 57332 17684 57384
rect 17736 57372 17742 57384
rect 18233 57375 18291 57381
rect 18233 57372 18245 57375
rect 17736 57344 18245 57372
rect 17736 57332 17742 57344
rect 18233 57341 18245 57344
rect 18279 57341 18291 57375
rect 18233 57335 18291 57341
rect 18506 57332 18512 57384
rect 18564 57372 18570 57384
rect 18877 57375 18935 57381
rect 18877 57372 18889 57375
rect 18564 57344 18889 57372
rect 18564 57332 18570 57344
rect 18877 57341 18889 57344
rect 18923 57341 18935 57375
rect 18877 57335 18935 57341
rect 19334 57332 19340 57384
rect 19392 57372 19398 57384
rect 20916 57381 20944 57412
rect 22462 57400 22468 57452
rect 22520 57440 22526 57452
rect 22520 57412 23060 57440
rect 22520 57400 22526 57412
rect 20257 57375 20315 57381
rect 20257 57372 20269 57375
rect 19392 57344 20269 57372
rect 19392 57332 19398 57344
rect 20257 57341 20269 57344
rect 20303 57341 20315 57375
rect 20257 57335 20315 57341
rect 20901 57375 20959 57381
rect 20901 57341 20913 57375
rect 20947 57341 20959 57375
rect 20901 57335 20959 57341
rect 20990 57332 20996 57384
rect 21048 57372 21054 57384
rect 21545 57375 21603 57381
rect 21545 57372 21557 57375
rect 21048 57344 21557 57372
rect 21048 57332 21054 57344
rect 21545 57341 21557 57344
rect 21591 57341 21603 57375
rect 21545 57335 21603 57341
rect 21634 57332 21640 57384
rect 21692 57372 21698 57384
rect 22925 57375 22983 57381
rect 22925 57372 22937 57375
rect 21692 57344 22937 57372
rect 21692 57332 21698 57344
rect 22925 57341 22937 57344
rect 22971 57341 22983 57375
rect 23032 57372 23060 57412
rect 23198 57400 23204 57452
rect 23256 57440 23262 57452
rect 23256 57412 24256 57440
rect 23256 57400 23262 57412
rect 24228 57381 24256 57412
rect 25608 57381 25636 57480
rect 31938 57468 31944 57520
rect 31996 57508 32002 57520
rect 53285 57511 53343 57517
rect 31996 57480 33180 57508
rect 31996 57468 32002 57480
rect 25682 57400 25688 57452
rect 25740 57440 25746 57452
rect 25740 57412 26924 57440
rect 25740 57400 25746 57412
rect 26896 57381 26924 57412
rect 27982 57400 27988 57452
rect 28040 57440 28046 57452
rect 28040 57412 28948 57440
rect 28040 57400 28046 57412
rect 23569 57375 23627 57381
rect 23569 57372 23581 57375
rect 23032 57344 23581 57372
rect 22925 57335 22983 57341
rect 23569 57341 23581 57344
rect 23615 57341 23627 57375
rect 23569 57335 23627 57341
rect 24213 57375 24271 57381
rect 24213 57341 24225 57375
rect 24259 57341 24271 57375
rect 24213 57335 24271 57341
rect 25593 57375 25651 57381
rect 25593 57341 25605 57375
rect 25639 57341 25651 57375
rect 25593 57335 25651 57341
rect 26237 57375 26295 57381
rect 26237 57341 26249 57375
rect 26283 57341 26295 57375
rect 26237 57335 26295 57341
rect 26881 57375 26939 57381
rect 26881 57341 26893 57375
rect 26927 57341 26939 57375
rect 26881 57335 26939 57341
rect 4341 57307 4399 57313
rect 4341 57273 4353 57307
rect 4387 57304 4399 57307
rect 4614 57304 4620 57316
rect 4387 57276 4620 57304
rect 4387 57273 4399 57276
rect 4341 57267 4399 57273
rect 4614 57264 4620 57276
rect 4672 57264 4678 57316
rect 5074 57196 5080 57248
rect 5132 57236 5138 57248
rect 5261 57239 5319 57245
rect 5261 57236 5273 57239
rect 5132 57208 5273 57236
rect 5132 57196 5138 57208
rect 5261 57205 5273 57208
rect 5307 57205 5319 57239
rect 5261 57199 5319 57205
rect 24854 57196 24860 57248
rect 24912 57236 24918 57248
rect 26252 57236 26280 57335
rect 27154 57332 27160 57384
rect 27212 57372 27218 57384
rect 28920 57381 28948 57412
rect 30374 57400 30380 57452
rect 30432 57440 30438 57452
rect 30432 57412 31064 57440
rect 30432 57400 30438 57412
rect 28261 57375 28319 57381
rect 28261 57372 28273 57375
rect 27212 57344 28273 57372
rect 27212 57332 27218 57344
rect 28261 57341 28273 57344
rect 28307 57341 28319 57375
rect 28261 57335 28319 57341
rect 28905 57375 28963 57381
rect 28905 57341 28917 57375
rect 28951 57341 28963 57375
rect 28905 57335 28963 57341
rect 28994 57332 29000 57384
rect 29052 57372 29058 57384
rect 29549 57375 29607 57381
rect 29549 57372 29561 57375
rect 29052 57344 29561 57372
rect 29052 57332 29058 57344
rect 29549 57341 29561 57344
rect 29595 57341 29607 57375
rect 29549 57335 29607 57341
rect 29638 57332 29644 57384
rect 29696 57372 29702 57384
rect 30929 57375 30987 57381
rect 30929 57372 30941 57375
rect 29696 57344 30941 57372
rect 29696 57332 29702 57344
rect 30929 57341 30941 57344
rect 30975 57341 30987 57375
rect 31036 57372 31064 57412
rect 31110 57400 31116 57452
rect 31168 57440 31174 57452
rect 31168 57412 32260 57440
rect 31168 57400 31174 57412
rect 32232 57381 32260 57412
rect 31573 57375 31631 57381
rect 31573 57372 31585 57375
rect 31036 57344 31585 57372
rect 30929 57335 30987 57341
rect 31573 57341 31585 57344
rect 31619 57341 31631 57375
rect 31573 57335 31631 57341
rect 32217 57375 32275 57381
rect 32217 57341 32229 57375
rect 32263 57341 32275 57375
rect 33152 57372 33180 57480
rect 53285 57477 53297 57511
rect 53331 57508 53343 57511
rect 55030 57508 55036 57520
rect 53331 57480 55036 57508
rect 53331 57477 53343 57480
rect 53285 57471 53343 57477
rect 55030 57468 55036 57480
rect 55088 57468 55094 57520
rect 55490 57508 55496 57520
rect 55451 57480 55496 57508
rect 55490 57468 55496 57480
rect 55548 57468 55554 57520
rect 56321 57511 56379 57517
rect 56321 57477 56333 57511
rect 56367 57477 56379 57511
rect 56321 57471 56379 57477
rect 33502 57400 33508 57452
rect 33560 57440 33566 57452
rect 33560 57412 34928 57440
rect 33560 57400 33566 57412
rect 34900 57381 34928 57412
rect 36630 57400 36636 57452
rect 36688 57440 36694 57452
rect 36688 57412 37596 57440
rect 36688 57400 36694 57412
rect 33597 57375 33655 57381
rect 33597 57372 33609 57375
rect 33152 57344 33609 57372
rect 32217 57335 32275 57341
rect 33597 57341 33609 57344
rect 33643 57341 33655 57375
rect 33597 57335 33655 57341
rect 34241 57375 34299 57381
rect 34241 57341 34253 57375
rect 34287 57341 34299 57375
rect 34241 57335 34299 57341
rect 34885 57375 34943 57381
rect 34885 57341 34897 57375
rect 34931 57341 34943 57375
rect 34885 57335 34943 57341
rect 32674 57264 32680 57316
rect 32732 57304 32738 57316
rect 34256 57304 34284 57335
rect 35250 57332 35256 57384
rect 35308 57372 35314 57384
rect 37568 57381 37596 57412
rect 39022 57400 39028 57452
rect 39080 57440 39086 57452
rect 39080 57412 40264 57440
rect 39080 57400 39086 57412
rect 36265 57375 36323 57381
rect 36265 57372 36277 57375
rect 35308 57344 36277 57372
rect 35308 57332 35314 57344
rect 36265 57341 36277 57344
rect 36311 57341 36323 57375
rect 36265 57335 36323 57341
rect 36909 57375 36967 57381
rect 36909 57341 36921 57375
rect 36955 57341 36967 57375
rect 36909 57335 36967 57341
rect 37553 57375 37611 57381
rect 37553 57341 37565 57375
rect 37599 57341 37611 57375
rect 37553 57335 37611 57341
rect 32732 57276 34284 57304
rect 32732 57264 32738 57276
rect 35894 57264 35900 57316
rect 35952 57304 35958 57316
rect 36924 57304 36952 57335
rect 37642 57332 37648 57384
rect 37700 57372 37706 57384
rect 40236 57381 40264 57412
rect 45370 57400 45376 57452
rect 45428 57440 45434 57452
rect 45428 57412 45600 57440
rect 45428 57400 45434 57412
rect 38933 57375 38991 57381
rect 38933 57372 38945 57375
rect 37700 57344 38945 57372
rect 37700 57332 37706 57344
rect 38933 57341 38945 57344
rect 38979 57341 38991 57375
rect 38933 57335 38991 57341
rect 39577 57375 39635 57381
rect 39577 57341 39589 57375
rect 39623 57341 39635 57375
rect 39577 57335 39635 57341
rect 40221 57375 40279 57381
rect 40221 57341 40233 57375
rect 40267 57341 40279 57375
rect 42150 57372 42156 57384
rect 42111 57344 42156 57372
rect 40221 57335 40279 57341
rect 35952 57276 36952 57304
rect 35952 57264 35958 57276
rect 38194 57264 38200 57316
rect 38252 57304 38258 57316
rect 39592 57304 39620 57335
rect 42150 57332 42156 57344
rect 42208 57332 42214 57384
rect 42978 57372 42984 57384
rect 42939 57344 42984 57372
rect 42978 57332 42984 57344
rect 43036 57332 43042 57384
rect 43714 57332 43720 57384
rect 43772 57372 43778 57384
rect 44269 57375 44327 57381
rect 44269 57372 44281 57375
rect 43772 57344 44281 57372
rect 43772 57332 43778 57344
rect 44269 57341 44281 57344
rect 44315 57341 44327 57375
rect 44269 57335 44327 57341
rect 44542 57332 44548 57384
rect 44600 57372 44606 57384
rect 45572 57381 45600 57412
rect 49234 57400 49240 57452
rect 49292 57440 49298 57452
rect 49292 57412 49832 57440
rect 49292 57400 49298 57412
rect 44913 57375 44971 57381
rect 44913 57372 44925 57375
rect 44600 57344 44925 57372
rect 44600 57332 44606 57344
rect 44913 57341 44925 57344
rect 44959 57341 44971 57375
rect 44913 57335 44971 57341
rect 45557 57375 45615 57381
rect 45557 57341 45569 57375
rect 45603 57341 45615 57375
rect 45557 57335 45615 57341
rect 46106 57332 46112 57384
rect 46164 57372 46170 57384
rect 46937 57375 46995 57381
rect 46937 57372 46949 57375
rect 46164 57344 46949 57372
rect 46164 57332 46170 57344
rect 46937 57341 46949 57344
rect 46983 57341 46995 57375
rect 46937 57335 46995 57341
rect 47026 57332 47032 57384
rect 47084 57372 47090 57384
rect 47581 57375 47639 57381
rect 47581 57372 47593 57375
rect 47084 57344 47593 57372
rect 47084 57332 47090 57344
rect 47581 57341 47593 57344
rect 47627 57341 47639 57375
rect 47581 57335 47639 57341
rect 47670 57332 47676 57384
rect 47728 57372 47734 57384
rect 48225 57375 48283 57381
rect 48225 57372 48237 57375
rect 47728 57344 48237 57372
rect 47728 57332 47734 57344
rect 48225 57341 48237 57344
rect 48271 57341 48283 57375
rect 48225 57335 48283 57341
rect 48498 57332 48504 57384
rect 48556 57372 48562 57384
rect 49605 57375 49663 57381
rect 49605 57372 49617 57375
rect 48556 57344 49617 57372
rect 48556 57332 48562 57344
rect 49605 57341 49617 57344
rect 49651 57341 49663 57375
rect 49804 57372 49832 57412
rect 50062 57400 50068 57452
rect 50120 57440 50126 57452
rect 52549 57443 52607 57449
rect 50120 57412 50936 57440
rect 50120 57400 50126 57412
rect 50908 57381 50936 57412
rect 52549 57409 52561 57443
rect 52595 57440 52607 57443
rect 54938 57440 54944 57452
rect 52595 57412 54944 57440
rect 52595 57409 52607 57412
rect 52549 57403 52607 57409
rect 54938 57400 54944 57412
rect 54996 57400 55002 57452
rect 56336 57440 56364 57471
rect 55324 57412 56364 57440
rect 50249 57375 50307 57381
rect 50249 57372 50261 57375
rect 49804 57344 50261 57372
rect 49605 57335 49663 57341
rect 50249 57341 50261 57344
rect 50295 57341 50307 57375
rect 50249 57335 50307 57341
rect 50893 57375 50951 57381
rect 50893 57341 50905 57375
rect 50939 57341 50951 57375
rect 50893 57335 50951 57341
rect 52365 57375 52423 57381
rect 52365 57341 52377 57375
rect 52411 57372 52423 57375
rect 55324 57372 55352 57412
rect 52411 57344 55352 57372
rect 52411 57341 52423 57344
rect 52365 57335 52423 57341
rect 55398 57332 55404 57384
rect 55456 57372 55462 57384
rect 55953 57375 56011 57381
rect 55953 57372 55965 57375
rect 55456 57344 55965 57372
rect 55456 57332 55462 57344
rect 55953 57341 55965 57344
rect 55999 57341 56011 57375
rect 55953 57335 56011 57341
rect 56137 57375 56195 57381
rect 56137 57341 56149 57375
rect 56183 57341 56195 57375
rect 56137 57335 56195 57341
rect 53098 57304 53104 57316
rect 38252 57276 39620 57304
rect 53059 57276 53104 57304
rect 38252 57264 38258 57276
rect 53098 57264 53104 57276
rect 53156 57264 53162 57316
rect 53834 57304 53840 57316
rect 53795 57276 53840 57304
rect 53834 57264 53840 57276
rect 53892 57264 53898 57316
rect 55309 57307 55367 57313
rect 55309 57273 55321 57307
rect 55355 57273 55367 57307
rect 55309 57267 55367 57273
rect 24912 57208 26280 57236
rect 55324 57236 55352 57267
rect 55766 57264 55772 57316
rect 55824 57304 55830 57316
rect 56152 57304 56180 57335
rect 57974 57304 57980 57316
rect 55824 57276 56180 57304
rect 57935 57276 57980 57304
rect 55824 57264 55830 57276
rect 57974 57264 57980 57276
rect 58032 57264 58038 57316
rect 58158 57304 58164 57316
rect 58119 57276 58164 57304
rect 58158 57264 58164 57276
rect 58216 57264 58222 57316
rect 58066 57236 58072 57248
rect 55324 57208 58072 57236
rect 24912 57196 24918 57208
rect 58066 57196 58072 57208
rect 58124 57196 58130 57248
rect 1104 57146 58880 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 50326 57146
rect 50378 57094 50390 57146
rect 50442 57094 50454 57146
rect 50506 57094 50518 57146
rect 50570 57094 58880 57146
rect 1104 57072 58880 57094
rect 53098 56992 53104 57044
rect 53156 57032 53162 57044
rect 56594 57032 56600 57044
rect 53156 57004 56600 57032
rect 53156 56992 53162 57004
rect 56594 56992 56600 57004
rect 56652 56992 56658 57044
rect 57974 56992 57980 57044
rect 58032 57032 58038 57044
rect 58161 57035 58219 57041
rect 58161 57032 58173 57035
rect 58032 57004 58173 57032
rect 58032 56992 58038 57004
rect 58161 57001 58173 57004
rect 58207 57001 58219 57035
rect 58161 56995 58219 57001
rect 1394 56896 1400 56908
rect 1355 56868 1400 56896
rect 1394 56856 1400 56868
rect 1452 56856 1458 56908
rect 2501 56899 2559 56905
rect 2501 56865 2513 56899
rect 2547 56896 2559 56899
rect 2682 56896 2688 56908
rect 2547 56868 2688 56896
rect 2547 56865 2559 56868
rect 2501 56859 2559 56865
rect 2682 56856 2688 56868
rect 2740 56856 2746 56908
rect 16114 56896 16120 56908
rect 16075 56868 16120 56896
rect 16114 56856 16120 56868
rect 16172 56856 16178 56908
rect 26418 56896 26424 56908
rect 26379 56868 26424 56896
rect 26418 56856 26424 56868
rect 26476 56856 26482 56908
rect 34238 56896 34244 56908
rect 34199 56868 34244 56896
rect 34238 56856 34244 56868
rect 34296 56856 34302 56908
rect 39758 56896 39764 56908
rect 39719 56868 39764 56896
rect 39758 56856 39764 56868
rect 39816 56856 39822 56908
rect 40586 56856 40592 56908
rect 40644 56896 40650 56908
rect 40957 56899 41015 56905
rect 40957 56896 40969 56899
rect 40644 56868 40969 56896
rect 40644 56856 40650 56868
rect 40957 56865 40969 56868
rect 41003 56865 41015 56899
rect 40957 56859 41015 56865
rect 41414 56856 41420 56908
rect 41472 56896 41478 56908
rect 41601 56899 41659 56905
rect 41601 56896 41613 56899
rect 41472 56868 41613 56896
rect 41472 56856 41478 56868
rect 41601 56865 41613 56868
rect 41647 56865 41659 56899
rect 41601 56859 41659 56865
rect 51074 56856 51080 56908
rect 51132 56896 51138 56908
rect 51445 56899 51503 56905
rect 51445 56896 51457 56899
rect 51132 56868 51457 56896
rect 51132 56856 51138 56868
rect 51445 56865 51457 56868
rect 51491 56865 51503 56899
rect 51445 56859 51503 56865
rect 51626 56856 51632 56908
rect 51684 56896 51690 56908
rect 52089 56899 52147 56905
rect 52089 56896 52101 56899
rect 51684 56868 52101 56896
rect 51684 56856 51690 56868
rect 52089 56865 52101 56868
rect 52135 56865 52147 56899
rect 52089 56859 52147 56865
rect 52454 56856 52460 56908
rect 52512 56896 52518 56908
rect 52733 56899 52791 56905
rect 52733 56896 52745 56899
rect 52512 56868 52745 56896
rect 52512 56856 52518 56868
rect 52733 56865 52745 56868
rect 52779 56865 52791 56899
rect 52733 56859 52791 56865
rect 53653 56899 53711 56905
rect 53653 56865 53665 56899
rect 53699 56896 53711 56899
rect 55582 56896 55588 56908
rect 53699 56868 55588 56896
rect 53699 56865 53711 56868
rect 53653 56859 53711 56865
rect 55582 56856 55588 56868
rect 55640 56856 55646 56908
rect 55766 56896 55772 56908
rect 55727 56868 55772 56896
rect 55766 56856 55772 56868
rect 55824 56856 55830 56908
rect 56873 56899 56931 56905
rect 56873 56865 56885 56899
rect 56919 56896 56931 56899
rect 57974 56896 57980 56908
rect 56919 56868 57980 56896
rect 56919 56865 56931 56868
rect 56873 56859 56931 56865
rect 57974 56856 57980 56868
rect 58032 56856 58038 56908
rect 4525 56831 4583 56837
rect 4525 56797 4537 56831
rect 4571 56797 4583 56831
rect 4706 56828 4712 56840
rect 4667 56800 4712 56828
rect 4525 56791 4583 56797
rect 4540 56760 4568 56791
rect 4706 56788 4712 56800
rect 4764 56788 4770 56840
rect 6365 56831 6423 56837
rect 6365 56797 6377 56831
rect 6411 56828 6423 56831
rect 53834 56828 53840 56840
rect 6411 56800 53840 56828
rect 6411 56797 6423 56800
rect 6365 56791 6423 56797
rect 53834 56788 53840 56800
rect 53892 56788 53898 56840
rect 55125 56831 55183 56837
rect 55125 56797 55137 56831
rect 55171 56828 55183 56831
rect 55171 56800 56272 56828
rect 55171 56797 55183 56800
rect 55125 56791 55183 56797
rect 5442 56760 5448 56772
rect 4540 56732 5448 56760
rect 5442 56720 5448 56732
rect 5500 56720 5506 56772
rect 54481 56763 54539 56769
rect 54481 56729 54493 56763
rect 54527 56760 54539 56763
rect 56134 56760 56140 56772
rect 54527 56732 56140 56760
rect 54527 56729 54539 56732
rect 54481 56723 54539 56729
rect 56134 56720 56140 56732
rect 56192 56720 56198 56772
rect 56244 56760 56272 56800
rect 56318 56788 56324 56840
rect 56376 56828 56382 56840
rect 57517 56831 57575 56837
rect 57517 56828 57529 56831
rect 56376 56800 57529 56828
rect 56376 56788 56382 56800
rect 57517 56797 57529 56800
rect 57563 56797 57575 56831
rect 57517 56791 57575 56797
rect 57606 56788 57612 56840
rect 57664 56828 57670 56840
rect 57701 56831 57759 56837
rect 57701 56828 57713 56831
rect 57664 56800 57713 56828
rect 57664 56788 57670 56800
rect 57701 56797 57713 56800
rect 57747 56797 57759 56831
rect 57701 56791 57759 56797
rect 56870 56760 56876 56772
rect 56244 56732 56876 56760
rect 56870 56720 56876 56732
rect 56928 56720 56934 56772
rect 57054 56760 57060 56772
rect 57015 56732 57060 56760
rect 57054 56720 57060 56732
rect 57112 56720 57118 56772
rect 3326 56692 3332 56704
rect 3287 56664 3332 56692
rect 3326 56652 3332 56664
rect 3384 56652 3390 56704
rect 55585 56695 55643 56701
rect 55585 56661 55597 56695
rect 55631 56692 55643 56695
rect 57698 56692 57704 56704
rect 55631 56664 57704 56692
rect 55631 56661 55643 56664
rect 55585 56655 55643 56661
rect 57698 56652 57704 56664
rect 57756 56652 57762 56704
rect 1104 56602 58880 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 58880 56602
rect 1104 56528 58880 56550
rect 382 56448 388 56500
rect 440 56488 446 56500
rect 1302 56488 1308 56500
rect 440 56460 1308 56488
rect 440 56448 446 56460
rect 1302 56448 1308 56460
rect 1360 56448 1366 56500
rect 4157 56491 4215 56497
rect 4157 56457 4169 56491
rect 4203 56488 4215 56491
rect 4614 56488 4620 56500
rect 4203 56460 4620 56488
rect 4203 56457 4215 56460
rect 4157 56451 4215 56457
rect 4614 56448 4620 56460
rect 4672 56448 4678 56500
rect 4706 56448 4712 56500
rect 4764 56488 4770 56500
rect 4801 56491 4859 56497
rect 4801 56488 4813 56491
rect 4764 56460 4813 56488
rect 4764 56448 4770 56460
rect 4801 56457 4813 56460
rect 4847 56457 4859 56491
rect 5442 56488 5448 56500
rect 5403 56460 5448 56488
rect 4801 56451 4859 56457
rect 5442 56448 5448 56460
rect 5500 56448 5506 56500
rect 53926 56448 53932 56500
rect 53984 56488 53990 56500
rect 54754 56488 54760 56500
rect 53984 56460 54760 56488
rect 53984 56448 53990 56460
rect 54754 56448 54760 56460
rect 54812 56448 54818 56500
rect 55033 56491 55091 56497
rect 55033 56457 55045 56491
rect 55079 56488 55091 56491
rect 56318 56488 56324 56500
rect 55079 56460 56324 56488
rect 55079 56457 55091 56460
rect 55033 56451 55091 56457
rect 56318 56448 56324 56460
rect 56376 56448 56382 56500
rect 56594 56488 56600 56500
rect 56555 56460 56600 56488
rect 56594 56448 56600 56460
rect 56652 56448 56658 56500
rect 58066 56488 58072 56500
rect 58027 56460 58072 56488
rect 58066 56448 58072 56460
rect 58124 56448 58130 56500
rect 2869 56423 2927 56429
rect 2869 56389 2881 56423
rect 2915 56420 2927 56423
rect 54389 56423 54447 56429
rect 2915 56392 3740 56420
rect 2915 56389 2927 56392
rect 2869 56383 2927 56389
rect 3326 56312 3332 56364
rect 3384 56352 3390 56364
rect 3712 56361 3740 56392
rect 54389 56389 54401 56423
rect 54435 56420 54447 56423
rect 55398 56420 55404 56432
rect 54435 56392 55404 56420
rect 54435 56389 54447 56392
rect 54389 56383 54447 56389
rect 55398 56380 55404 56392
rect 55456 56380 55462 56432
rect 55493 56423 55551 56429
rect 55493 56389 55505 56423
rect 55539 56389 55551 56423
rect 55493 56383 55551 56389
rect 3513 56355 3571 56361
rect 3513 56352 3525 56355
rect 3384 56324 3525 56352
rect 3384 56312 3390 56324
rect 3513 56321 3525 56324
rect 3559 56321 3571 56355
rect 3513 56315 3571 56321
rect 3697 56355 3755 56361
rect 3697 56321 3709 56355
rect 3743 56321 3755 56355
rect 55122 56352 55128 56364
rect 3697 56315 3755 56321
rect 52288 56324 55128 56352
rect 1118 56244 1124 56296
rect 1176 56284 1182 56296
rect 1397 56287 1455 56293
rect 1397 56284 1409 56287
rect 1176 56256 1409 56284
rect 1176 56244 1182 56256
rect 1397 56253 1409 56256
rect 1443 56253 1455 56287
rect 1397 56247 1455 56253
rect 1946 56244 1952 56296
rect 2004 56284 2010 56296
rect 52288 56293 52316 56324
rect 55122 56312 55128 56324
rect 55180 56312 55186 56364
rect 55508 56352 55536 56383
rect 56226 56380 56232 56432
rect 56284 56420 56290 56432
rect 58250 56420 58256 56432
rect 56284 56392 58256 56420
rect 56284 56380 56290 56392
rect 58250 56380 58256 56392
rect 58308 56380 58314 56432
rect 56321 56355 56379 56361
rect 56321 56352 56333 56355
rect 55508 56324 56333 56352
rect 56321 56321 56333 56324
rect 56367 56321 56379 56355
rect 56321 56315 56379 56321
rect 56870 56312 56876 56364
rect 56928 56352 56934 56364
rect 57517 56355 57575 56361
rect 57517 56352 57529 56355
rect 56928 56324 57529 56352
rect 56928 56312 56934 56324
rect 57517 56321 57529 56324
rect 57563 56321 57575 56355
rect 57698 56352 57704 56364
rect 57659 56324 57704 56352
rect 57517 56315 57575 56321
rect 57698 56312 57704 56324
rect 57756 56312 57762 56364
rect 2041 56287 2099 56293
rect 2041 56284 2053 56287
rect 2004 56256 2053 56284
rect 2004 56244 2010 56256
rect 2041 56253 2053 56256
rect 2087 56253 2099 56287
rect 2041 56247 2099 56253
rect 3053 56287 3111 56293
rect 3053 56253 3065 56287
rect 3099 56284 3111 56287
rect 4617 56287 4675 56293
rect 4617 56284 4629 56287
rect 3099 56256 4629 56284
rect 3099 56253 3111 56256
rect 3053 56247 3111 56253
rect 3712 56228 3740 56256
rect 4617 56253 4629 56256
rect 4663 56253 4675 56287
rect 4617 56247 4675 56253
rect 51629 56287 51687 56293
rect 51629 56253 51641 56287
rect 51675 56253 51687 56287
rect 51629 56247 51687 56253
rect 52273 56287 52331 56293
rect 52273 56253 52285 56287
rect 52319 56253 52331 56287
rect 52273 56247 52331 56253
rect 52917 56287 52975 56293
rect 52917 56253 52929 56287
rect 52963 56284 52975 56287
rect 53190 56284 53196 56296
rect 52963 56256 53196 56284
rect 52963 56253 52975 56256
rect 52917 56247 52975 56253
rect 3694 56176 3700 56228
rect 3752 56176 3758 56228
rect 51644 56216 51672 56247
rect 53190 56244 53196 56256
rect 53248 56244 53254 56296
rect 55677 56287 55735 56293
rect 55677 56253 55689 56287
rect 55723 56284 55735 56287
rect 55766 56284 55772 56296
rect 55723 56256 55772 56284
rect 55723 56253 55735 56256
rect 55677 56247 55735 56253
rect 55766 56244 55772 56256
rect 55824 56244 55830 56296
rect 56134 56284 56140 56296
rect 56095 56256 56140 56284
rect 56134 56244 56140 56256
rect 56192 56244 56198 56296
rect 57146 56216 57152 56228
rect 51644 56188 57152 56216
rect 57146 56176 57152 56188
rect 57204 56176 57210 56228
rect 1104 56058 58880 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 50326 56058
rect 50378 56006 50390 56058
rect 50442 56006 50454 56058
rect 50506 56006 50518 56058
rect 50570 56006 58880 56058
rect 1104 55984 58880 56006
rect 55585 55947 55643 55953
rect 55585 55913 55597 55947
rect 55631 55944 55643 55947
rect 57606 55944 57612 55956
rect 55631 55916 57612 55944
rect 55631 55913 55643 55916
rect 55585 55907 55643 55913
rect 57606 55904 57612 55916
rect 57664 55904 57670 55956
rect 57241 55879 57299 55885
rect 52380 55848 56456 55876
rect 1394 55808 1400 55820
rect 1355 55780 1400 55808
rect 1394 55768 1400 55780
rect 1452 55768 1458 55820
rect 3510 55768 3516 55820
rect 3568 55808 3574 55820
rect 52380 55817 52408 55848
rect 4249 55811 4307 55817
rect 4249 55808 4261 55811
rect 3568 55780 4261 55808
rect 3568 55768 3574 55780
rect 4249 55777 4261 55780
rect 4295 55777 4307 55811
rect 4249 55771 4307 55777
rect 52365 55811 52423 55817
rect 52365 55777 52377 55811
rect 52411 55777 52423 55811
rect 52365 55771 52423 55777
rect 53009 55811 53067 55817
rect 53009 55777 53021 55811
rect 53055 55777 53067 55811
rect 53009 55771 53067 55777
rect 53653 55811 53711 55817
rect 53653 55777 53665 55811
rect 53699 55808 53711 55811
rect 54018 55808 54024 55820
rect 53699 55780 54024 55808
rect 53699 55777 53711 55780
rect 53653 55771 53711 55777
rect 53024 55740 53052 55771
rect 54018 55768 54024 55780
rect 54076 55768 54082 55820
rect 54297 55811 54355 55817
rect 54297 55777 54309 55811
rect 54343 55808 54355 55811
rect 55674 55808 55680 55820
rect 54343 55780 55680 55808
rect 54343 55777 54355 55780
rect 54297 55771 54355 55777
rect 55674 55768 55680 55780
rect 55732 55768 55738 55820
rect 55766 55768 55772 55820
rect 55824 55808 55830 55820
rect 55824 55780 55869 55808
rect 55824 55768 55830 55780
rect 55306 55740 55312 55752
rect 53024 55712 55312 55740
rect 55306 55700 55312 55712
rect 55364 55700 55370 55752
rect 56428 55672 56456 55848
rect 57241 55845 57253 55879
rect 57287 55876 57299 55879
rect 58250 55876 58256 55888
rect 57287 55848 58256 55876
rect 57287 55845 57299 55848
rect 57241 55839 57299 55845
rect 58250 55836 58256 55848
rect 58308 55836 58314 55888
rect 57330 55768 57336 55820
rect 57388 55808 57394 55820
rect 57977 55811 58035 55817
rect 57977 55808 57989 55811
rect 57388 55780 57989 55808
rect 57388 55768 57394 55780
rect 57977 55777 57989 55780
rect 58023 55777 58035 55811
rect 57977 55771 58035 55777
rect 56502 55700 56508 55752
rect 56560 55740 56566 55752
rect 57425 55743 57483 55749
rect 57425 55740 57437 55743
rect 56560 55712 57437 55740
rect 56560 55700 56566 55712
rect 57425 55709 57437 55712
rect 57471 55709 57483 55743
rect 58710 55740 58716 55752
rect 57425 55703 57483 55709
rect 57532 55712 58716 55740
rect 57532 55672 57560 55712
rect 58710 55700 58716 55712
rect 58768 55700 58774 55752
rect 58158 55672 58164 55684
rect 56428 55644 57560 55672
rect 58119 55644 58164 55672
rect 58158 55632 58164 55644
rect 58216 55632 58222 55684
rect 55125 55607 55183 55613
rect 55125 55573 55137 55607
rect 55171 55604 55183 55607
rect 55490 55604 55496 55616
rect 55171 55576 55496 55604
rect 55171 55573 55183 55576
rect 55125 55567 55183 55573
rect 55490 55564 55496 55576
rect 55548 55564 55554 55616
rect 1104 55514 58880 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 58880 55514
rect 1104 55440 58880 55462
rect 55033 55335 55091 55341
rect 55033 55301 55045 55335
rect 55079 55332 55091 55335
rect 55079 55304 57560 55332
rect 55079 55301 55091 55304
rect 55033 55295 55091 55301
rect 55677 55267 55735 55273
rect 55677 55233 55689 55267
rect 55723 55264 55735 55267
rect 57238 55264 57244 55276
rect 55723 55236 57244 55264
rect 55723 55233 55735 55236
rect 55677 55227 55735 55233
rect 57238 55224 57244 55236
rect 57296 55224 57302 55276
rect 57532 55273 57560 55304
rect 57517 55267 57575 55273
rect 57517 55233 57529 55267
rect 57563 55233 57575 55267
rect 57517 55227 57575 55233
rect 53926 55156 53932 55208
rect 53984 55196 53990 55208
rect 54205 55199 54263 55205
rect 54205 55196 54217 55199
rect 53984 55168 54217 55196
rect 53984 55156 53990 55168
rect 54205 55165 54217 55168
rect 54251 55165 54263 55199
rect 56318 55196 56324 55208
rect 56279 55168 56324 55196
rect 54205 55159 54263 55165
rect 56318 55156 56324 55168
rect 56376 55156 56382 55208
rect 56594 55156 56600 55208
rect 56652 55196 56658 55208
rect 57701 55199 57759 55205
rect 57701 55196 57713 55199
rect 56652 55168 57713 55196
rect 56652 55156 56658 55168
rect 57701 55165 57713 55168
rect 57747 55165 57759 55199
rect 57701 55159 57759 55165
rect 57974 55156 57980 55208
rect 58032 55196 58038 55208
rect 58161 55199 58219 55205
rect 58161 55196 58173 55199
rect 58032 55168 58173 55196
rect 58032 55156 58038 55168
rect 58161 55165 58173 55168
rect 58207 55165 58219 55199
rect 58161 55159 58219 55165
rect 56870 55128 56876 55140
rect 56831 55100 56876 55128
rect 56870 55088 56876 55100
rect 56928 55088 56934 55140
rect 57054 55128 57060 55140
rect 57015 55100 57060 55128
rect 57054 55088 57060 55100
rect 57112 55088 57118 55140
rect 56134 55060 56140 55072
rect 56095 55032 56140 55060
rect 56134 55020 56140 55032
rect 56192 55020 56198 55072
rect 1104 54970 58880 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 50326 54970
rect 50378 54918 50390 54970
rect 50442 54918 50454 54970
rect 50506 54918 50518 54970
rect 50570 54918 58880 54970
rect 1104 54896 58880 54918
rect 55766 54856 55772 54868
rect 55679 54828 55772 54856
rect 55766 54816 55772 54828
rect 55824 54856 55830 54868
rect 56318 54856 56324 54868
rect 55824 54828 56324 54856
rect 55824 54816 55830 54828
rect 56318 54816 56324 54828
rect 56376 54816 56382 54868
rect 57330 54856 57336 54868
rect 57291 54828 57336 54856
rect 57330 54816 57336 54828
rect 57388 54816 57394 54868
rect 56226 54788 56232 54800
rect 54312 54760 56232 54788
rect 1394 54720 1400 54732
rect 1355 54692 1400 54720
rect 1394 54680 1400 54692
rect 1452 54680 1458 54732
rect 54312 54729 54340 54760
rect 56226 54748 56232 54760
rect 56284 54748 56290 54800
rect 54297 54723 54355 54729
rect 54297 54689 54309 54723
rect 54343 54689 54355 54723
rect 54297 54683 54355 54689
rect 55125 54723 55183 54729
rect 55125 54689 55137 54723
rect 55171 54689 55183 54723
rect 55125 54683 55183 54689
rect 55140 54584 55168 54683
rect 55306 54680 55312 54732
rect 55364 54720 55370 54732
rect 55585 54723 55643 54729
rect 55585 54720 55597 54723
rect 55364 54692 55597 54720
rect 55364 54680 55370 54692
rect 55585 54689 55597 54692
rect 55631 54689 55643 54723
rect 55585 54683 55643 54689
rect 56134 54680 56140 54732
rect 56192 54720 56198 54732
rect 56873 54723 56931 54729
rect 56873 54720 56885 54723
rect 56192 54692 56885 54720
rect 56192 54680 56198 54692
rect 56873 54689 56885 54692
rect 56919 54689 56931 54723
rect 57974 54720 57980 54732
rect 57935 54692 57980 54720
rect 56873 54683 56931 54689
rect 57974 54680 57980 54692
rect 58032 54680 58038 54732
rect 55490 54612 55496 54664
rect 55548 54652 55554 54664
rect 56689 54655 56747 54661
rect 56689 54652 56701 54655
rect 55548 54624 56701 54652
rect 55548 54612 55554 54624
rect 56689 54621 56701 54624
rect 56735 54621 56747 54655
rect 56689 54615 56747 54621
rect 56318 54584 56324 54596
rect 55140 54556 56324 54584
rect 56318 54544 56324 54556
rect 56376 54544 56382 54596
rect 58158 54584 58164 54596
rect 58119 54556 58164 54584
rect 58158 54544 58164 54556
rect 58216 54544 58222 54596
rect 54938 54516 54944 54528
rect 54899 54488 54944 54516
rect 54938 54476 54944 54488
rect 54996 54476 55002 54528
rect 1104 54426 58880 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 58880 54426
rect 1104 54352 58880 54374
rect 56137 54315 56195 54321
rect 56137 54281 56149 54315
rect 56183 54312 56195 54315
rect 56594 54312 56600 54324
rect 56183 54284 56600 54312
rect 56183 54281 56195 54284
rect 56137 54275 56195 54281
rect 56594 54272 56600 54284
rect 56652 54272 56658 54324
rect 56870 54272 56876 54324
rect 56928 54312 56934 54324
rect 57885 54315 57943 54321
rect 57885 54312 57897 54315
rect 56928 54284 57897 54312
rect 56928 54272 56934 54284
rect 57885 54281 57897 54284
rect 57931 54281 57943 54315
rect 57885 54275 57943 54281
rect 54938 54136 54944 54188
rect 54996 54176 55002 54188
rect 54996 54148 56456 54176
rect 54996 54136 55002 54148
rect 55490 54108 55496 54120
rect 55451 54080 55496 54108
rect 55490 54068 55496 54080
rect 55548 54068 55554 54120
rect 56318 54108 56324 54120
rect 56279 54080 56324 54108
rect 56318 54068 56324 54080
rect 56376 54068 56382 54120
rect 56428 54108 56456 54148
rect 57238 54136 57244 54188
rect 57296 54176 57302 54188
rect 57517 54179 57575 54185
rect 57517 54176 57529 54179
rect 57296 54148 57529 54176
rect 57296 54136 57302 54148
rect 57517 54145 57529 54148
rect 57563 54145 57575 54179
rect 57517 54139 57575 54145
rect 57701 54111 57759 54117
rect 57701 54108 57713 54111
rect 56428 54080 57713 54108
rect 57701 54077 57713 54080
rect 57747 54077 57759 54111
rect 57701 54071 57759 54077
rect 56873 54043 56931 54049
rect 56873 54009 56885 54043
rect 56919 54040 56931 54043
rect 57422 54040 57428 54052
rect 56919 54012 57428 54040
rect 56919 54009 56931 54012
rect 56873 54003 56931 54009
rect 57422 54000 57428 54012
rect 57480 54000 57486 54052
rect 56962 53972 56968 53984
rect 56923 53944 56968 53972
rect 56962 53932 56968 53944
rect 57020 53932 57026 53984
rect 1104 53882 58880 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 50326 53882
rect 50378 53830 50390 53882
rect 50442 53830 50454 53882
rect 50506 53830 50518 53882
rect 50570 53830 58880 53882
rect 1104 53808 58880 53830
rect 1394 53632 1400 53644
rect 1355 53604 1400 53632
rect 1394 53592 1400 53604
rect 1452 53592 1458 53644
rect 55582 53632 55588 53644
rect 55543 53604 55588 53632
rect 55582 53592 55588 53604
rect 55640 53592 55646 53644
rect 56410 53524 56416 53576
rect 56468 53564 56474 53576
rect 57057 53567 57115 53573
rect 57057 53564 57069 53567
rect 56468 53536 57069 53564
rect 56468 53524 56474 53536
rect 57057 53533 57069 53536
rect 57103 53533 57115 53567
rect 57238 53564 57244 53576
rect 57199 53536 57244 53564
rect 57057 53527 57115 53533
rect 57238 53524 57244 53536
rect 57296 53524 57302 53576
rect 57422 53496 57428 53508
rect 57383 53468 57428 53496
rect 57422 53456 57428 53468
rect 57480 53456 57486 53508
rect 1104 53338 58880 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 58880 53338
rect 1104 53264 58880 53286
rect 56410 53224 56416 53236
rect 56371 53196 56416 53224
rect 56410 53184 56416 53196
rect 56468 53184 56474 53236
rect 56873 53227 56931 53233
rect 56873 53193 56885 53227
rect 56919 53224 56931 53227
rect 57238 53224 57244 53236
rect 56919 53196 57244 53224
rect 56919 53193 56931 53196
rect 56873 53187 56931 53193
rect 57238 53184 57244 53196
rect 57296 53184 57302 53236
rect 57974 53224 57980 53236
rect 57935 53196 57980 53224
rect 57974 53184 57980 53196
rect 58032 53184 58038 53236
rect 55769 53091 55827 53097
rect 55769 53057 55781 53091
rect 55815 53088 55827 53091
rect 57517 53091 57575 53097
rect 57517 53088 57529 53091
rect 55815 53060 57529 53088
rect 55815 53057 55827 53060
rect 55769 53051 55827 53057
rect 57517 53057 57529 53060
rect 57563 53057 57575 53091
rect 57517 53051 57575 53057
rect 1394 53020 1400 53032
rect 1355 52992 1400 53020
rect 1394 52980 1400 52992
rect 1452 52980 1458 53032
rect 56318 52980 56324 53032
rect 56376 53020 56382 53032
rect 57057 53023 57115 53029
rect 57057 53020 57069 53023
rect 56376 52992 57069 53020
rect 56376 52980 56382 52992
rect 57057 52989 57069 52992
rect 57103 52989 57115 53023
rect 57057 52983 57115 52989
rect 57238 52980 57244 53032
rect 57296 53020 57302 53032
rect 57701 53023 57759 53029
rect 57701 53020 57713 53023
rect 57296 52992 57713 53020
rect 57296 52980 57302 52992
rect 57701 52989 57713 52992
rect 57747 52989 57759 53023
rect 57701 52983 57759 52989
rect 1104 52794 58880 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 50326 52794
rect 50378 52742 50390 52794
rect 50442 52742 50454 52794
rect 50506 52742 50518 52794
rect 50570 52742 58880 52794
rect 1104 52720 58880 52742
rect 57238 52680 57244 52692
rect 57199 52652 57244 52680
rect 57238 52640 57244 52652
rect 57296 52640 57302 52692
rect 57422 52544 57428 52556
rect 57383 52516 57428 52544
rect 57422 52504 57428 52516
rect 57480 52504 57486 52556
rect 57974 52544 57980 52556
rect 57935 52516 57980 52544
rect 57974 52504 57980 52516
rect 58032 52504 58038 52556
rect 57882 52436 57888 52488
rect 57940 52476 57946 52488
rect 58161 52479 58219 52485
rect 58161 52476 58173 52479
rect 57940 52448 58173 52476
rect 57940 52436 57946 52448
rect 58161 52445 58173 52448
rect 58207 52445 58219 52479
rect 58161 52439 58219 52445
rect 1104 52250 58880 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 58880 52250
rect 1104 52176 58880 52198
rect 57974 52136 57980 52148
rect 57935 52108 57980 52136
rect 57974 52096 57980 52108
rect 58032 52096 58038 52148
rect 56137 52071 56195 52077
rect 56137 52037 56149 52071
rect 56183 52037 56195 52071
rect 56137 52031 56195 52037
rect 56152 52000 56180 52031
rect 57701 52003 57759 52009
rect 57701 52000 57713 52003
rect 56152 51972 57713 52000
rect 57701 51969 57713 51972
rect 57747 51969 57759 52003
rect 57701 51963 57759 51969
rect 1394 51932 1400 51944
rect 1355 51904 1400 51932
rect 1394 51892 1400 51904
rect 1452 51892 1458 51944
rect 55490 51932 55496 51944
rect 55451 51904 55496 51932
rect 55490 51892 55496 51904
rect 55548 51892 55554 51944
rect 56321 51935 56379 51941
rect 56321 51901 56333 51935
rect 56367 51932 56379 51935
rect 57514 51932 57520 51944
rect 56367 51904 57192 51932
rect 57475 51904 57520 51932
rect 56367 51901 56379 51904
rect 56321 51895 56379 51901
rect 56870 51864 56876 51876
rect 56831 51836 56876 51864
rect 56870 51824 56876 51836
rect 56928 51824 56934 51876
rect 57054 51864 57060 51876
rect 57015 51836 57060 51864
rect 57054 51824 57060 51836
rect 57112 51824 57118 51876
rect 57164 51864 57192 51904
rect 57514 51892 57520 51904
rect 57572 51892 57578 51944
rect 57422 51864 57428 51876
rect 57164 51836 57428 51864
rect 57422 51824 57428 51836
rect 57480 51824 57486 51876
rect 1104 51706 58880 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 50326 51706
rect 50378 51654 50390 51706
rect 50442 51654 50454 51706
rect 50506 51654 50518 51706
rect 50570 51654 58880 51706
rect 1104 51632 58880 51654
rect 56870 51552 56876 51604
rect 56928 51592 56934 51604
rect 57701 51595 57759 51601
rect 57701 51592 57713 51595
rect 56928 51564 57713 51592
rect 56928 51552 56934 51564
rect 57701 51561 57713 51564
rect 57747 51561 57759 51595
rect 57701 51555 57759 51561
rect 55125 51459 55183 51465
rect 55125 51425 55137 51459
rect 55171 51456 55183 51459
rect 57514 51456 57520 51468
rect 55171 51428 57520 51456
rect 55171 51425 55183 51428
rect 55125 51419 55183 51425
rect 57514 51416 57520 51428
rect 57572 51416 57578 51468
rect 55769 51391 55827 51397
rect 55769 51357 55781 51391
rect 55815 51388 55827 51391
rect 57057 51391 57115 51397
rect 57057 51388 57069 51391
rect 55815 51360 57069 51388
rect 55815 51357 55827 51360
rect 55769 51351 55827 51357
rect 57057 51357 57069 51360
rect 57103 51357 57115 51391
rect 57238 51388 57244 51400
rect 57199 51360 57244 51388
rect 57057 51351 57115 51357
rect 57238 51348 57244 51360
rect 57296 51348 57302 51400
rect 1104 51162 58880 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 58880 51162
rect 1104 51088 58880 51110
rect 56597 51051 56655 51057
rect 56597 51017 56609 51051
rect 56643 51048 56655 51051
rect 57238 51048 57244 51060
rect 56643 51020 57244 51048
rect 56643 51017 56655 51020
rect 56597 51011 56655 51017
rect 57238 51008 57244 51020
rect 57296 51008 57302 51060
rect 1394 50844 1400 50856
rect 1355 50816 1400 50844
rect 1394 50804 1400 50816
rect 1452 50804 1458 50856
rect 56137 50847 56195 50853
rect 56137 50813 56149 50847
rect 56183 50813 56195 50847
rect 56137 50807 56195 50813
rect 56152 50776 56180 50807
rect 56318 50804 56324 50856
rect 56376 50844 56382 50856
rect 56781 50847 56839 50853
rect 56781 50844 56793 50847
rect 56376 50816 56793 50844
rect 56376 50804 56382 50816
rect 56781 50813 56793 50816
rect 56827 50813 56839 50847
rect 57422 50844 57428 50856
rect 57383 50816 57428 50844
rect 56781 50807 56839 50813
rect 57422 50804 57428 50816
rect 57480 50804 57486 50856
rect 57514 50776 57520 50788
rect 56152 50748 57520 50776
rect 57514 50736 57520 50748
rect 57572 50736 57578 50788
rect 57974 50776 57980 50788
rect 57935 50748 57980 50776
rect 57974 50736 57980 50748
rect 58032 50736 58038 50788
rect 58158 50776 58164 50788
rect 58119 50748 58164 50776
rect 58158 50736 58164 50748
rect 58216 50736 58222 50788
rect 57241 50711 57299 50717
rect 57241 50677 57253 50711
rect 57287 50708 57299 50711
rect 57698 50708 57704 50720
rect 57287 50680 57704 50708
rect 57287 50677 57299 50680
rect 57241 50671 57299 50677
rect 57698 50668 57704 50680
rect 57756 50668 57762 50720
rect 1104 50618 58880 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 50326 50618
rect 50378 50566 50390 50618
rect 50442 50566 50454 50618
rect 50506 50566 50518 50618
rect 50570 50566 58880 50618
rect 1104 50544 58880 50566
rect 57974 50464 57980 50516
rect 58032 50504 58038 50516
rect 58161 50507 58219 50513
rect 58161 50504 58173 50507
rect 58032 50476 58173 50504
rect 58032 50464 58038 50476
rect 58161 50473 58173 50476
rect 58207 50473 58219 50507
rect 58161 50467 58219 50473
rect 1394 50368 1400 50380
rect 1355 50340 1400 50368
rect 1394 50328 1400 50340
rect 1452 50328 1458 50380
rect 56870 50368 56876 50380
rect 56831 50340 56876 50368
rect 56870 50328 56876 50340
rect 56928 50328 56934 50380
rect 57514 50368 57520 50380
rect 57475 50340 57520 50368
rect 57514 50328 57520 50340
rect 57572 50328 57578 50380
rect 57698 50368 57704 50380
rect 57659 50340 57704 50368
rect 57698 50328 57704 50340
rect 57756 50328 57762 50380
rect 57054 50232 57060 50244
rect 57015 50204 57060 50232
rect 57054 50192 57060 50204
rect 57112 50192 57118 50244
rect 55769 50167 55827 50173
rect 55769 50133 55781 50167
rect 55815 50164 55827 50167
rect 57146 50164 57152 50176
rect 55815 50136 57152 50164
rect 55815 50133 55827 50136
rect 55769 50127 55827 50133
rect 57146 50124 57152 50136
rect 57204 50124 57210 50176
rect 1104 50074 58880 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 58880 50074
rect 1104 50000 58880 50022
rect 56318 49920 56324 49972
rect 56376 49960 56382 49972
rect 56689 49963 56747 49969
rect 56689 49960 56701 49963
rect 56376 49932 56701 49960
rect 56376 49920 56382 49932
rect 56689 49929 56701 49932
rect 56735 49929 56747 49963
rect 56689 49923 56747 49929
rect 56870 49920 56876 49972
rect 56928 49960 56934 49972
rect 57517 49963 57575 49969
rect 57517 49960 57529 49963
rect 56928 49932 57529 49960
rect 56928 49920 56934 49932
rect 57517 49929 57529 49932
rect 57563 49929 57575 49963
rect 57517 49923 57575 49929
rect 55861 49895 55919 49901
rect 55861 49861 55873 49895
rect 55907 49892 55919 49895
rect 55907 49864 57376 49892
rect 55907 49861 55919 49864
rect 55861 49855 55919 49861
rect 55950 49784 55956 49836
rect 56008 49824 56014 49836
rect 57146 49824 57152 49836
rect 56008 49796 56548 49824
rect 57107 49796 57152 49824
rect 56008 49784 56014 49796
rect 55214 49756 55220 49768
rect 55175 49728 55220 49756
rect 55214 49716 55220 49728
rect 55272 49716 55278 49768
rect 56045 49759 56103 49765
rect 56045 49725 56057 49759
rect 56091 49756 56103 49759
rect 56318 49756 56324 49768
rect 56091 49728 56324 49756
rect 56091 49725 56103 49728
rect 56045 49719 56103 49725
rect 56318 49716 56324 49728
rect 56376 49716 56382 49768
rect 56520 49765 56548 49796
rect 57146 49784 57152 49796
rect 57204 49784 57210 49836
rect 57348 49833 57376 49864
rect 57333 49827 57391 49833
rect 57333 49793 57345 49827
rect 57379 49793 57391 49827
rect 57333 49787 57391 49793
rect 56505 49759 56563 49765
rect 56505 49725 56517 49759
rect 56551 49725 56563 49759
rect 56505 49719 56563 49725
rect 1104 49530 58880 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 50326 49530
rect 50378 49478 50390 49530
rect 50442 49478 50454 49530
rect 50506 49478 50518 49530
rect 50570 49478 58880 49530
rect 1104 49456 58880 49478
rect 1394 49280 1400 49292
rect 1355 49252 1400 49280
rect 1394 49240 1400 49252
rect 1452 49240 1458 49292
rect 57422 49280 57428 49292
rect 57335 49252 57428 49280
rect 57422 49240 57428 49252
rect 57480 49280 57486 49292
rect 57790 49280 57796 49292
rect 57480 49252 57796 49280
rect 57480 49240 57486 49252
rect 57790 49240 57796 49252
rect 57848 49240 57854 49292
rect 57974 49280 57980 49292
rect 57935 49252 57980 49280
rect 57974 49240 57980 49252
rect 58032 49240 58038 49292
rect 58158 49280 58164 49292
rect 58119 49252 58164 49280
rect 58158 49240 58164 49252
rect 58216 49240 58222 49292
rect 55766 49076 55772 49088
rect 55727 49048 55772 49076
rect 55766 49036 55772 49048
rect 55824 49036 55830 49088
rect 57241 49079 57299 49085
rect 57241 49045 57253 49079
rect 57287 49076 57299 49079
rect 57698 49076 57704 49088
rect 57287 49048 57704 49076
rect 57287 49045 57299 49048
rect 57241 49039 57299 49045
rect 57698 49036 57704 49048
rect 57756 49036 57762 49088
rect 1104 48986 58880 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 58880 48986
rect 1104 48912 58880 48934
rect 57974 48872 57980 48884
rect 57935 48844 57980 48872
rect 57974 48832 57980 48844
rect 58032 48832 58038 48884
rect 57054 48804 57060 48816
rect 57015 48776 57060 48804
rect 57054 48764 57060 48776
rect 57112 48764 57118 48816
rect 55766 48696 55772 48748
rect 55824 48736 55830 48748
rect 57517 48739 57575 48745
rect 57517 48736 57529 48739
rect 55824 48708 57529 48736
rect 55824 48696 55830 48708
rect 57517 48705 57529 48708
rect 57563 48705 57575 48739
rect 57698 48736 57704 48748
rect 57659 48708 57704 48736
rect 57517 48699 57575 48705
rect 57698 48696 57704 48708
rect 57756 48696 57762 48748
rect 55490 48668 55496 48680
rect 55451 48640 55496 48668
rect 55490 48628 55496 48640
rect 55548 48628 55554 48680
rect 56321 48671 56379 48677
rect 56321 48637 56333 48671
rect 56367 48668 56379 48671
rect 57054 48668 57060 48680
rect 56367 48640 57060 48668
rect 56367 48637 56379 48640
rect 56321 48631 56379 48637
rect 57054 48628 57060 48640
rect 57112 48628 57118 48680
rect 56873 48603 56931 48609
rect 56873 48569 56885 48603
rect 56919 48600 56931 48603
rect 57422 48600 57428 48612
rect 56919 48572 57428 48600
rect 56919 48569 56931 48572
rect 56873 48563 56931 48569
rect 57422 48560 57428 48572
rect 57480 48560 57486 48612
rect 1104 48442 58880 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 50326 48442
rect 50378 48390 50390 48442
rect 50442 48390 50454 48442
rect 50506 48390 50518 48442
rect 50570 48390 58880 48442
rect 1104 48368 58880 48390
rect 1394 48192 1400 48204
rect 1355 48164 1400 48192
rect 1394 48152 1400 48164
rect 1452 48152 1458 48204
rect 57054 48192 57060 48204
rect 57015 48164 57060 48192
rect 57054 48152 57060 48164
rect 57112 48152 57118 48204
rect 55490 48084 55496 48136
rect 55548 48124 55554 48136
rect 57241 48127 57299 48133
rect 57241 48124 57253 48127
rect 55548 48096 57253 48124
rect 55548 48084 55554 48096
rect 57241 48093 57253 48096
rect 57287 48093 57299 48127
rect 57241 48087 57299 48093
rect 57422 48056 57428 48068
rect 57383 48028 57428 48056
rect 57422 48016 57428 48028
rect 57480 48016 57486 48068
rect 55769 47991 55827 47997
rect 55769 47957 55781 47991
rect 55815 47988 55827 47991
rect 57514 47988 57520 48000
rect 55815 47960 57520 47988
rect 55815 47957 55827 47960
rect 55769 47951 55827 47957
rect 57514 47948 57520 47960
rect 57572 47948 57578 48000
rect 1104 47898 58880 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 58880 47898
rect 1104 47824 58880 47846
rect 55490 47784 55496 47796
rect 55451 47756 55496 47784
rect 55490 47744 55496 47756
rect 55548 47744 55554 47796
rect 56137 47719 56195 47725
rect 56137 47685 56149 47719
rect 56183 47716 56195 47719
rect 56183 47688 57744 47716
rect 56183 47685 56195 47688
rect 56137 47679 56195 47685
rect 57054 47648 57060 47660
rect 57015 47620 57060 47648
rect 57054 47608 57060 47620
rect 57112 47608 57118 47660
rect 57514 47648 57520 47660
rect 57475 47620 57520 47648
rect 57514 47608 57520 47620
rect 57572 47608 57578 47660
rect 57716 47657 57744 47688
rect 57701 47651 57759 47657
rect 57701 47617 57713 47651
rect 57747 47617 57759 47651
rect 57701 47611 57759 47617
rect 55674 47580 55680 47592
rect 55635 47552 55680 47580
rect 55674 47540 55680 47552
rect 55732 47540 55738 47592
rect 56321 47583 56379 47589
rect 56321 47549 56333 47583
rect 56367 47580 56379 47583
rect 57790 47580 57796 47592
rect 56367 47552 57796 47580
rect 56367 47549 56379 47552
rect 56321 47543 56379 47549
rect 57790 47540 57796 47552
rect 57848 47540 57854 47592
rect 56873 47515 56931 47521
rect 56873 47481 56885 47515
rect 56919 47512 56931 47515
rect 58161 47515 58219 47521
rect 58161 47512 58173 47515
rect 56919 47484 58173 47512
rect 56919 47481 56931 47484
rect 56873 47475 56931 47481
rect 58161 47481 58173 47484
rect 58207 47481 58219 47515
rect 58161 47475 58219 47481
rect 1104 47354 58880 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 50326 47354
rect 50378 47302 50390 47354
rect 50442 47302 50454 47354
rect 50506 47302 50518 47354
rect 50570 47302 58880 47354
rect 1104 47280 58880 47302
rect 1394 47104 1400 47116
rect 1355 47076 1400 47104
rect 1394 47064 1400 47076
rect 1452 47064 1458 47116
rect 54297 47107 54355 47113
rect 54297 47073 54309 47107
rect 54343 47104 54355 47107
rect 55214 47104 55220 47116
rect 54343 47076 55220 47104
rect 54343 47073 54355 47076
rect 54297 47067 54355 47073
rect 55214 47064 55220 47076
rect 55272 47064 55278 47116
rect 55585 47107 55643 47113
rect 55585 47073 55597 47107
rect 55631 47104 55643 47107
rect 55950 47104 55956 47116
rect 55631 47076 55956 47104
rect 55631 47073 55643 47076
rect 55585 47067 55643 47073
rect 55950 47064 55956 47076
rect 56008 47064 56014 47116
rect 57238 47104 57244 47116
rect 57199 47076 57244 47104
rect 57238 47064 57244 47076
rect 57296 47064 57302 47116
rect 57422 47104 57428 47116
rect 57383 47076 57428 47104
rect 57422 47064 57428 47076
rect 57480 47064 57486 47116
rect 57974 47104 57980 47116
rect 57935 47076 57980 47104
rect 57974 47064 57980 47076
rect 58032 47064 58038 47116
rect 55125 46971 55183 46977
rect 55125 46937 55137 46971
rect 55171 46968 55183 46971
rect 57514 46968 57520 46980
rect 55171 46940 57520 46968
rect 55171 46937 55183 46940
rect 55125 46931 55183 46937
rect 57514 46928 57520 46940
rect 57572 46928 57578 46980
rect 57882 46928 57888 46980
rect 57940 46968 57946 46980
rect 58161 46971 58219 46977
rect 58161 46968 58173 46971
rect 57940 46940 58173 46968
rect 57940 46928 57946 46940
rect 58161 46937 58173 46940
rect 58207 46937 58219 46971
rect 58161 46931 58219 46937
rect 55674 46860 55680 46912
rect 55732 46900 55738 46912
rect 55769 46903 55827 46909
rect 55769 46900 55781 46903
rect 55732 46872 55781 46900
rect 55732 46860 55738 46872
rect 55769 46869 55781 46872
rect 55815 46869 55827 46903
rect 55769 46863 55827 46869
rect 1104 46810 58880 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 58880 46810
rect 1104 46736 58880 46758
rect 56965 46699 57023 46705
rect 56965 46665 56977 46699
rect 57011 46696 57023 46699
rect 57238 46696 57244 46708
rect 57011 46668 57244 46696
rect 57011 46665 57023 46668
rect 56965 46659 57023 46665
rect 57238 46656 57244 46668
rect 57296 46656 57302 46708
rect 55677 46631 55735 46637
rect 55677 46597 55689 46631
rect 55723 46628 55735 46631
rect 55723 46600 56548 46628
rect 55723 46597 55735 46600
rect 55677 46591 55735 46597
rect 55030 46520 55036 46572
rect 55088 46560 55094 46572
rect 56520 46569 56548 46600
rect 56321 46563 56379 46569
rect 56321 46560 56333 46563
rect 55088 46532 56333 46560
rect 55088 46520 55094 46532
rect 56321 46529 56333 46532
rect 56367 46529 56379 46563
rect 56321 46523 56379 46529
rect 56505 46563 56563 46569
rect 56505 46529 56517 46563
rect 56551 46529 56563 46563
rect 56505 46523 56563 46529
rect 58161 46563 58219 46569
rect 58161 46529 58173 46563
rect 58207 46560 58219 46563
rect 58250 46560 58256 46572
rect 58207 46532 58256 46560
rect 58207 46529 58219 46532
rect 58161 46523 58219 46529
rect 58250 46520 58256 46532
rect 58308 46520 58314 46572
rect 1394 46492 1400 46504
rect 1355 46464 1400 46492
rect 1394 46452 1400 46464
rect 1452 46452 1458 46504
rect 54389 46495 54447 46501
rect 54389 46461 54401 46495
rect 54435 46492 54447 46495
rect 54754 46492 54760 46504
rect 54435 46464 54760 46492
rect 54435 46461 54447 46464
rect 54389 46455 54447 46461
rect 54754 46452 54760 46464
rect 54812 46452 54818 46504
rect 55217 46495 55275 46501
rect 55217 46461 55229 46495
rect 55263 46461 55275 46495
rect 55217 46455 55275 46461
rect 55232 46424 55260 46455
rect 55674 46452 55680 46504
rect 55732 46492 55738 46504
rect 55861 46495 55919 46501
rect 55861 46492 55873 46495
rect 55732 46464 55873 46492
rect 55732 46452 55738 46464
rect 55861 46461 55873 46464
rect 55907 46461 55919 46495
rect 55861 46455 55919 46461
rect 57517 46427 57575 46433
rect 57517 46424 57529 46427
rect 55232 46396 57529 46424
rect 57517 46393 57529 46396
rect 57563 46393 57575 46427
rect 57517 46387 57575 46393
rect 57606 46384 57612 46436
rect 57664 46424 57670 46436
rect 57664 46396 57709 46424
rect 57664 46384 57670 46396
rect 1104 46266 58880 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 50326 46266
rect 50378 46214 50390 46266
rect 50442 46214 50454 46266
rect 50506 46214 50518 46266
rect 50570 46214 58880 46266
rect 1104 46192 58880 46214
rect 55030 46152 55036 46164
rect 54991 46124 55036 46152
rect 55030 46112 55036 46124
rect 55088 46112 55094 46164
rect 55585 46155 55643 46161
rect 55585 46121 55597 46155
rect 55631 46152 55643 46155
rect 57606 46152 57612 46164
rect 55631 46124 57612 46152
rect 55631 46121 55643 46124
rect 55585 46115 55643 46121
rect 57606 46112 57612 46124
rect 57664 46112 57670 46164
rect 57790 46112 57796 46164
rect 57848 46152 57854 46164
rect 58161 46155 58219 46161
rect 58161 46152 58173 46155
rect 57848 46124 58173 46152
rect 57848 46112 57854 46124
rect 58161 46121 58173 46124
rect 58207 46121 58219 46155
rect 58161 46115 58219 46121
rect 53653 46019 53711 46025
rect 53653 45985 53665 46019
rect 53699 45985 53711 46019
rect 54938 46016 54944 46028
rect 54899 45988 54944 46016
rect 53653 45979 53711 45985
rect 53668 45948 53696 45979
rect 54938 45976 54944 45988
rect 54996 45976 55002 46028
rect 55125 46019 55183 46025
rect 55125 45985 55137 46019
rect 55171 45985 55183 46019
rect 55766 46016 55772 46028
rect 55727 45988 55772 46016
rect 55125 45979 55183 45985
rect 55030 45948 55036 45960
rect 53668 45920 55036 45948
rect 55030 45908 55036 45920
rect 55088 45908 55094 45960
rect 51534 45840 51540 45892
rect 51592 45880 51598 45892
rect 55140 45880 55168 45979
rect 55766 45976 55772 45988
rect 55824 45976 55830 46028
rect 55950 45976 55956 46028
rect 56008 46016 56014 46028
rect 57241 46019 57299 46025
rect 57241 46016 57253 46019
rect 56008 45988 57253 46016
rect 56008 45976 56014 45988
rect 57241 45985 57253 45988
rect 57287 45985 57299 46019
rect 57241 45979 57299 45985
rect 57977 46019 58035 46025
rect 57977 45985 57989 46019
rect 58023 46016 58035 46019
rect 58250 46016 58256 46028
rect 58023 45988 58256 46016
rect 58023 45985 58035 45988
rect 57977 45979 58035 45985
rect 58250 45976 58256 45988
rect 58308 45976 58314 46028
rect 51592 45852 55168 45880
rect 51592 45840 51598 45852
rect 55766 45840 55772 45892
rect 55824 45880 55830 45892
rect 57425 45883 57483 45889
rect 57425 45880 57437 45883
rect 55824 45852 57437 45880
rect 55824 45840 55830 45852
rect 57425 45849 57437 45852
rect 57471 45849 57483 45883
rect 57425 45843 57483 45849
rect 54481 45815 54539 45821
rect 54481 45781 54493 45815
rect 54527 45812 54539 45815
rect 56502 45812 56508 45824
rect 54527 45784 56508 45812
rect 54527 45781 54539 45784
rect 54481 45775 54539 45781
rect 56502 45772 56508 45784
rect 56560 45772 56566 45824
rect 1104 45722 58880 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 58880 45722
rect 1104 45648 58880 45670
rect 57054 45540 57060 45552
rect 57015 45512 57060 45540
rect 57054 45500 57060 45512
rect 57112 45500 57118 45552
rect 57974 45540 57980 45552
rect 57935 45512 57980 45540
rect 57974 45500 57980 45512
rect 58032 45500 58038 45552
rect 57514 45472 57520 45484
rect 57475 45444 57520 45472
rect 57514 45432 57520 45444
rect 57572 45432 57578 45484
rect 1394 45404 1400 45416
rect 1355 45376 1400 45404
rect 1394 45364 1400 45376
rect 1452 45364 1458 45416
rect 53926 45364 53932 45416
rect 53984 45404 53990 45416
rect 54021 45407 54079 45413
rect 54021 45404 54033 45407
rect 53984 45376 54033 45404
rect 53984 45364 53990 45376
rect 54021 45373 54033 45376
rect 54067 45373 54079 45407
rect 54202 45404 54208 45416
rect 54163 45376 54208 45404
rect 54021 45367 54079 45373
rect 54202 45364 54208 45376
rect 54260 45364 54266 45416
rect 54849 45407 54907 45413
rect 54849 45373 54861 45407
rect 54895 45404 54907 45407
rect 54938 45404 54944 45416
rect 54895 45376 54944 45404
rect 54895 45373 54907 45376
rect 54849 45367 54907 45373
rect 52914 45296 52920 45348
rect 52972 45336 52978 45348
rect 54864 45336 54892 45367
rect 54938 45364 54944 45376
rect 54996 45364 55002 45416
rect 55033 45407 55091 45413
rect 55033 45373 55045 45407
rect 55079 45404 55091 45407
rect 55122 45404 55128 45416
rect 55079 45376 55128 45404
rect 55079 45373 55091 45376
rect 55033 45367 55091 45373
rect 55122 45364 55128 45376
rect 55180 45364 55186 45416
rect 55674 45404 55680 45416
rect 55635 45376 55680 45404
rect 55674 45364 55680 45376
rect 55732 45364 55738 45416
rect 56321 45407 56379 45413
rect 56321 45373 56333 45407
rect 56367 45404 56379 45407
rect 57606 45404 57612 45416
rect 56367 45376 57612 45404
rect 56367 45373 56379 45376
rect 56321 45367 56379 45373
rect 57606 45364 57612 45376
rect 57664 45364 57670 45416
rect 57701 45407 57759 45413
rect 57701 45373 57713 45407
rect 57747 45404 57759 45407
rect 58066 45404 58072 45416
rect 57747 45376 58072 45404
rect 57747 45373 57759 45376
rect 57701 45367 57759 45373
rect 58066 45364 58072 45376
rect 58124 45364 58130 45416
rect 52972 45308 54892 45336
rect 56873 45339 56931 45345
rect 52972 45296 52978 45308
rect 56873 45305 56885 45339
rect 56919 45336 56931 45339
rect 57330 45336 57336 45348
rect 56919 45308 57336 45336
rect 56919 45305 56931 45308
rect 56873 45299 56931 45305
rect 57330 45296 57336 45308
rect 57388 45296 57394 45348
rect 54110 45268 54116 45280
rect 54071 45240 54116 45268
rect 54110 45228 54116 45240
rect 54168 45228 54174 45280
rect 54941 45271 54999 45277
rect 54941 45237 54953 45271
rect 54987 45268 54999 45271
rect 55398 45268 55404 45280
rect 54987 45240 55404 45268
rect 54987 45237 54999 45240
rect 54941 45231 54999 45237
rect 55398 45228 55404 45240
rect 55456 45228 55462 45280
rect 55493 45271 55551 45277
rect 55493 45237 55505 45271
rect 55539 45268 55551 45271
rect 56042 45268 56048 45280
rect 55539 45240 56048 45268
rect 55539 45237 55551 45240
rect 55493 45231 55551 45237
rect 56042 45228 56048 45240
rect 56100 45228 56106 45280
rect 56137 45271 56195 45277
rect 56137 45237 56149 45271
rect 56183 45268 56195 45271
rect 57698 45268 57704 45280
rect 56183 45240 57704 45268
rect 56183 45237 56195 45240
rect 56137 45231 56195 45237
rect 57698 45228 57704 45240
rect 57756 45228 57762 45280
rect 1104 45178 58880 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 50326 45178
rect 50378 45126 50390 45178
rect 50442 45126 50454 45178
rect 50506 45126 50518 45178
rect 50570 45126 58880 45178
rect 1104 45104 58880 45126
rect 52730 45024 52736 45076
rect 52788 45064 52794 45076
rect 54021 45067 54079 45073
rect 54021 45064 54033 45067
rect 52788 45036 54033 45064
rect 52788 45024 52794 45036
rect 54021 45033 54033 45036
rect 54067 45033 54079 45067
rect 57330 45064 57336 45076
rect 57291 45036 57336 45064
rect 54021 45027 54079 45033
rect 57330 45024 57336 45036
rect 57388 45024 57394 45076
rect 54202 44996 54208 45008
rect 54036 44968 54208 44996
rect 52086 44888 52092 44940
rect 52144 44928 52150 44940
rect 54036 44937 54064 44968
rect 54202 44956 54208 44968
rect 54260 44996 54266 45008
rect 54260 44968 54892 44996
rect 54260 44956 54266 44968
rect 52253 44931 52311 44937
rect 52253 44928 52265 44931
rect 52144 44900 52265 44928
rect 52144 44888 52150 44900
rect 52253 44897 52265 44900
rect 52299 44897 52311 44931
rect 54021 44931 54079 44937
rect 54021 44928 54033 44931
rect 52253 44891 52311 44897
rect 53392 44900 54033 44928
rect 51258 44820 51264 44872
rect 51316 44860 51322 44872
rect 51997 44863 52055 44869
rect 51997 44860 52009 44863
rect 51316 44832 52009 44860
rect 51316 44820 51322 44832
rect 51997 44829 52009 44832
rect 52043 44829 52055 44863
rect 51997 44823 52055 44829
rect 53392 44801 53420 44900
rect 54021 44897 54033 44900
rect 54067 44897 54079 44931
rect 54021 44891 54079 44897
rect 54110 44888 54116 44940
rect 54168 44928 54174 44940
rect 54294 44928 54300 44940
rect 54168 44900 54300 44928
rect 54168 44888 54174 44900
rect 54294 44888 54300 44900
rect 54352 44928 54358 44940
rect 54864 44937 54892 44968
rect 54389 44931 54447 44937
rect 54389 44928 54401 44931
rect 54352 44900 54401 44928
rect 54352 44888 54358 44900
rect 54389 44897 54401 44900
rect 54435 44897 54447 44931
rect 54389 44891 54447 44897
rect 54849 44931 54907 44937
rect 54849 44897 54861 44931
rect 54895 44897 54907 44931
rect 55582 44928 55588 44940
rect 55543 44900 55588 44928
rect 54849 44891 54907 44897
rect 55582 44888 55588 44900
rect 55640 44888 55646 44940
rect 56042 44888 56048 44940
rect 56100 44928 56106 44940
rect 56873 44931 56931 44937
rect 56873 44928 56885 44931
rect 56100 44900 56885 44928
rect 56100 44888 56106 44900
rect 56873 44897 56885 44900
rect 56919 44897 56931 44931
rect 57974 44928 57980 44940
rect 57935 44900 57980 44928
rect 56873 44891 56931 44897
rect 57974 44888 57980 44900
rect 58032 44888 58038 44940
rect 53837 44863 53895 44869
rect 53837 44829 53849 44863
rect 53883 44860 53895 44863
rect 53926 44860 53932 44872
rect 53883 44832 53932 44860
rect 53883 44829 53895 44832
rect 53837 44823 53895 44829
rect 53926 44820 53932 44832
rect 53984 44860 53990 44872
rect 55600 44860 55628 44888
rect 56686 44860 56692 44872
rect 53984 44832 55628 44860
rect 56647 44832 56692 44860
rect 53984 44820 53990 44832
rect 56686 44820 56692 44832
rect 56744 44820 56750 44872
rect 53377 44795 53435 44801
rect 53377 44761 53389 44795
rect 53423 44761 53435 44795
rect 53377 44755 53435 44761
rect 54386 44752 54392 44804
rect 54444 44792 54450 44804
rect 55677 44795 55735 44801
rect 55677 44792 55689 44795
rect 54444 44764 55689 44792
rect 54444 44752 54450 44764
rect 55677 44761 55689 44764
rect 55723 44761 55735 44795
rect 58158 44792 58164 44804
rect 58119 44764 58164 44792
rect 55677 44755 55735 44761
rect 58158 44752 58164 44764
rect 58216 44752 58222 44804
rect 54938 44724 54944 44736
rect 54899 44696 54944 44724
rect 54938 44684 54944 44696
rect 54996 44684 55002 44736
rect 1104 44634 58880 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 58880 44634
rect 1104 44560 58880 44582
rect 51074 44520 51080 44532
rect 50172 44492 51080 44520
rect 50172 44393 50200 44492
rect 51074 44480 51080 44492
rect 51132 44520 51138 44532
rect 51258 44520 51264 44532
rect 51132 44492 51264 44520
rect 51132 44480 51138 44492
rect 51258 44480 51264 44492
rect 51316 44480 51322 44532
rect 51997 44523 52055 44529
rect 51997 44489 52009 44523
rect 52043 44520 52055 44523
rect 52086 44520 52092 44532
rect 52043 44492 52092 44520
rect 52043 44489 52055 44492
rect 51997 44483 52055 44489
rect 52086 44480 52092 44492
rect 52144 44480 52150 44532
rect 52917 44523 52975 44529
rect 52917 44489 52929 44523
rect 52963 44520 52975 44523
rect 56686 44520 56692 44532
rect 52963 44492 56692 44520
rect 52963 44489 52975 44492
rect 52917 44483 52975 44489
rect 56686 44480 56692 44492
rect 56744 44480 56750 44532
rect 57974 44520 57980 44532
rect 57935 44492 57980 44520
rect 57974 44480 57980 44492
rect 58032 44480 58038 44532
rect 55582 44412 55588 44464
rect 55640 44452 55646 44464
rect 55861 44455 55919 44461
rect 55861 44452 55873 44455
rect 55640 44424 55873 44452
rect 55640 44412 55646 44424
rect 55861 44421 55873 44424
rect 55907 44421 55919 44455
rect 55861 44415 55919 44421
rect 50157 44387 50215 44393
rect 50157 44353 50169 44387
rect 50203 44353 50215 44387
rect 52546 44384 52552 44396
rect 50157 44347 50215 44353
rect 52012 44356 52552 44384
rect 1394 44316 1400 44328
rect 1355 44288 1400 44316
rect 1394 44276 1400 44288
rect 1452 44276 1458 44328
rect 50706 44276 50712 44328
rect 50764 44316 50770 44328
rect 52012 44325 52040 44356
rect 52546 44344 52552 44356
rect 52604 44344 52610 44396
rect 56502 44344 56508 44396
rect 56560 44384 56566 44396
rect 57517 44387 57575 44393
rect 57517 44384 57529 44387
rect 56560 44356 57529 44384
rect 56560 44344 56566 44356
rect 57517 44353 57529 44356
rect 57563 44353 57575 44387
rect 57698 44384 57704 44396
rect 57659 44356 57704 44384
rect 57517 44347 57575 44353
rect 57698 44344 57704 44356
rect 57756 44344 57762 44396
rect 51997 44319 52055 44325
rect 50764 44288 51074 44316
rect 50764 44276 50770 44288
rect 50424 44251 50482 44257
rect 50424 44217 50436 44251
rect 50470 44248 50482 44251
rect 50614 44248 50620 44260
rect 50470 44220 50620 44248
rect 50470 44217 50482 44220
rect 50424 44211 50482 44217
rect 50614 44208 50620 44220
rect 50672 44208 50678 44260
rect 51046 44248 51074 44288
rect 51997 44285 52009 44319
rect 52043 44285 52055 44319
rect 51997 44279 52055 44285
rect 52181 44319 52239 44325
rect 52181 44285 52193 44319
rect 52227 44285 52239 44319
rect 52181 44279 52239 44285
rect 52196 44248 52224 44279
rect 52454 44276 52460 44328
rect 52512 44316 52518 44328
rect 52914 44316 52920 44328
rect 52512 44288 52920 44316
rect 52512 44276 52518 44288
rect 52914 44276 52920 44288
rect 52972 44276 52978 44328
rect 53101 44319 53159 44325
rect 53101 44285 53113 44319
rect 53147 44316 53159 44319
rect 54386 44316 54392 44328
rect 53147 44288 54392 44316
rect 53147 44285 53159 44288
rect 53101 44279 53159 44285
rect 54386 44276 54392 44288
rect 54444 44276 54450 44328
rect 54478 44276 54484 44328
rect 54536 44316 54542 44328
rect 54536 44288 54581 44316
rect 54536 44276 54542 44288
rect 51046 44220 52224 44248
rect 54748 44251 54806 44257
rect 54748 44217 54760 44251
rect 54794 44248 54806 44251
rect 55122 44248 55128 44260
rect 54794 44220 55128 44248
rect 54794 44217 54806 44220
rect 54748 44211 54806 44217
rect 55122 44208 55128 44220
rect 55180 44208 55186 44260
rect 56870 44248 56876 44260
rect 56831 44220 56876 44248
rect 56870 44208 56876 44220
rect 56928 44208 56934 44260
rect 57054 44248 57060 44260
rect 57015 44220 57060 44248
rect 57054 44208 57060 44220
rect 57112 44208 57118 44260
rect 51442 44140 51448 44192
rect 51500 44180 51506 44192
rect 51537 44183 51595 44189
rect 51537 44180 51549 44183
rect 51500 44152 51549 44180
rect 51500 44140 51506 44152
rect 51537 44149 51549 44152
rect 51583 44149 51595 44183
rect 51537 44143 51595 44149
rect 1104 44090 58880 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 58880 44090
rect 1104 44016 58880 44038
rect 50433 43979 50491 43985
rect 50433 43945 50445 43979
rect 50479 43976 50491 43979
rect 50614 43976 50620 43988
rect 50479 43948 50620 43976
rect 50479 43945 50491 43948
rect 50433 43939 50491 43945
rect 50614 43936 50620 43948
rect 50672 43936 50678 43988
rect 51534 43976 51540 43988
rect 51495 43948 51540 43976
rect 51534 43936 51540 43948
rect 51592 43936 51598 43988
rect 52546 43976 52552 43988
rect 52507 43948 52552 43976
rect 52546 43936 52552 43948
rect 52604 43936 52610 43988
rect 55122 43976 55128 43988
rect 55083 43948 55128 43976
rect 55122 43936 55128 43948
rect 55180 43936 55186 43988
rect 56870 43936 56876 43988
rect 56928 43976 56934 43988
rect 57517 43979 57575 43985
rect 57517 43976 57529 43979
rect 56928 43948 57529 43976
rect 56928 43936 56934 43948
rect 57517 43945 57529 43948
rect 57563 43945 57575 43979
rect 57517 43939 57575 43945
rect 57977 43979 58035 43985
rect 57977 43945 57989 43979
rect 58023 43976 58035 43979
rect 58066 43976 58072 43988
rect 58023 43948 58072 43976
rect 58023 43945 58035 43948
rect 57977 43939 58035 43945
rect 58066 43936 58072 43948
rect 58124 43936 58130 43988
rect 50706 43908 50712 43920
rect 50356 43880 50712 43908
rect 50356 43849 50384 43880
rect 50706 43868 50712 43880
rect 50764 43868 50770 43920
rect 52638 43908 52644 43920
rect 52380 43880 52644 43908
rect 50341 43843 50399 43849
rect 50341 43809 50353 43843
rect 50387 43809 50399 43843
rect 50341 43803 50399 43809
rect 50525 43843 50583 43849
rect 50525 43809 50537 43843
rect 50571 43840 50583 43843
rect 51166 43840 51172 43852
rect 50571 43812 51172 43840
rect 50571 43809 50583 43812
rect 50525 43803 50583 43809
rect 51166 43800 51172 43812
rect 51224 43800 51230 43852
rect 51442 43840 51448 43852
rect 51403 43812 51448 43840
rect 51442 43800 51448 43812
rect 51500 43800 51506 43852
rect 52380 43849 52408 43880
rect 52638 43868 52644 43880
rect 52696 43868 52702 43920
rect 54938 43868 54944 43920
rect 54996 43908 55002 43920
rect 54996 43880 55260 43908
rect 54996 43868 55002 43880
rect 52365 43843 52423 43849
rect 52365 43809 52377 43843
rect 52411 43809 52423 43843
rect 52730 43840 52736 43852
rect 52691 43812 52736 43840
rect 52365 43803 52423 43809
rect 52730 43800 52736 43812
rect 52788 43800 52794 43852
rect 53190 43800 53196 43852
rect 53248 43840 53254 43852
rect 53469 43843 53527 43849
rect 53469 43840 53481 43843
rect 53248 43812 53481 43840
rect 53248 43800 53254 43812
rect 53469 43809 53481 43812
rect 53515 43809 53527 43843
rect 54110 43840 54116 43852
rect 54071 43812 54116 43840
rect 53469 43803 53527 43809
rect 52181 43775 52239 43781
rect 52181 43741 52193 43775
rect 52227 43772 52239 43775
rect 52748 43772 52776 43800
rect 52227 43744 52776 43772
rect 53484 43772 53512 43803
rect 54110 43800 54116 43812
rect 54168 43800 54174 43852
rect 54294 43840 54300 43852
rect 54255 43812 54300 43840
rect 54294 43800 54300 43812
rect 54352 43800 54358 43852
rect 54386 43800 54392 43852
rect 54444 43840 54450 43852
rect 54573 43843 54631 43849
rect 54444 43812 54489 43840
rect 54444 43800 54450 43812
rect 54573 43809 54585 43843
rect 54619 43840 54631 43843
rect 54956 43840 54984 43868
rect 55232 43849 55260 43880
rect 54619 43812 54984 43840
rect 55033 43843 55091 43849
rect 54619 43809 54631 43812
rect 54573 43803 54631 43809
rect 55033 43809 55045 43843
rect 55079 43809 55091 43843
rect 55033 43803 55091 43809
rect 55217 43843 55275 43849
rect 55217 43809 55229 43843
rect 55263 43809 55275 43843
rect 55217 43803 55275 43809
rect 53484 43744 54800 43772
rect 52227 43741 52239 43744
rect 52181 43735 52239 43741
rect 53285 43707 53343 43713
rect 53285 43673 53297 43707
rect 53331 43704 53343 43707
rect 53331 43676 54156 43704
rect 53331 43673 53343 43676
rect 53285 43667 53343 43673
rect 53926 43636 53932 43648
rect 53887 43608 53932 43636
rect 53926 43596 53932 43608
rect 53984 43596 53990 43648
rect 54128 43636 54156 43676
rect 54202 43664 54208 43716
rect 54260 43704 54266 43716
rect 54772 43704 54800 43744
rect 54846 43732 54852 43784
rect 54904 43772 54910 43784
rect 55048 43772 55076 43803
rect 55398 43800 55404 43852
rect 55456 43840 55462 43852
rect 56873 43843 56931 43849
rect 56873 43840 56885 43843
rect 55456 43812 56885 43840
rect 55456 43800 55462 43812
rect 56873 43809 56885 43812
rect 56919 43809 56931 43843
rect 56873 43803 56931 43809
rect 57606 43800 57612 43852
rect 57664 43840 57670 43852
rect 58161 43843 58219 43849
rect 58161 43840 58173 43843
rect 57664 43812 58173 43840
rect 57664 43800 57670 43812
rect 58161 43809 58173 43812
rect 58207 43809 58219 43843
rect 58161 43803 58219 43809
rect 54904 43744 55076 43772
rect 57057 43775 57115 43781
rect 54904 43732 54910 43744
rect 57057 43741 57069 43775
rect 57103 43741 57115 43775
rect 57057 43735 57115 43741
rect 55674 43704 55680 43716
rect 54260 43676 54305 43704
rect 54772 43676 55680 43704
rect 54260 43664 54266 43676
rect 55674 43664 55680 43676
rect 55732 43664 55738 43716
rect 57072 43636 57100 43735
rect 54128 43608 57100 43636
rect 1104 43546 58880 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 58880 43546
rect 1104 43472 58880 43494
rect 52638 43392 52644 43444
rect 52696 43432 52702 43444
rect 54021 43435 54079 43441
rect 54021 43432 54033 43435
rect 52696 43404 54033 43432
rect 52696 43392 52702 43404
rect 54021 43401 54033 43404
rect 54067 43401 54079 43435
rect 54021 43395 54079 43401
rect 52730 43324 52736 43376
rect 52788 43364 52794 43376
rect 52788 43336 52960 43364
rect 52788 43324 52794 43336
rect 50525 43299 50583 43305
rect 50525 43265 50537 43299
rect 50571 43296 50583 43299
rect 51166 43296 51172 43308
rect 50571 43268 51172 43296
rect 50571 43265 50583 43268
rect 50525 43259 50583 43265
rect 51166 43256 51172 43268
rect 51224 43296 51230 43308
rect 51224 43268 51304 43296
rect 51224 43256 51230 43268
rect 1394 43228 1400 43240
rect 1355 43200 1400 43228
rect 1394 43188 1400 43200
rect 1452 43188 1458 43240
rect 50433 43231 50491 43237
rect 50433 43197 50445 43231
rect 50479 43228 50491 43231
rect 50614 43228 50620 43240
rect 50479 43200 50620 43228
rect 50479 43197 50491 43200
rect 50433 43191 50491 43197
rect 50614 43188 50620 43200
rect 50672 43188 50678 43240
rect 51276 43237 51304 43268
rect 52638 43256 52644 43308
rect 52696 43296 52702 43308
rect 52932 43305 52960 43336
rect 54202 43324 54208 43376
rect 54260 43364 54266 43376
rect 54389 43367 54447 43373
rect 54389 43364 54401 43367
rect 54260 43336 54401 43364
rect 54260 43324 54266 43336
rect 54389 43333 54401 43336
rect 54435 43364 54447 43367
rect 55030 43364 55036 43376
rect 54435 43336 55036 43364
rect 54435 43333 54447 43336
rect 54389 43327 54447 43333
rect 55030 43324 55036 43336
rect 55088 43324 55094 43376
rect 52825 43299 52883 43305
rect 52825 43296 52837 43299
rect 52696 43268 52837 43296
rect 52696 43256 52702 43268
rect 52825 43265 52837 43268
rect 52871 43265 52883 43299
rect 52825 43259 52883 43265
rect 52917 43299 52975 43305
rect 52917 43265 52929 43299
rect 52963 43265 52975 43299
rect 52917 43259 52975 43265
rect 54110 43256 54116 43308
rect 54168 43296 54174 43308
rect 54481 43299 54539 43305
rect 54481 43296 54493 43299
rect 54168 43268 54493 43296
rect 54168 43256 54174 43268
rect 54481 43265 54493 43268
rect 54527 43296 54539 43299
rect 54938 43296 54944 43308
rect 54527 43268 54944 43296
rect 54527 43265 54539 43268
rect 54481 43259 54539 43265
rect 54938 43256 54944 43268
rect 54996 43256 55002 43308
rect 55048 43296 55076 43324
rect 56965 43299 57023 43305
rect 56965 43296 56977 43299
rect 55048 43268 55168 43296
rect 55140 43240 55168 43268
rect 56060 43268 56977 43296
rect 51077 43231 51135 43237
rect 51077 43197 51089 43231
rect 51123 43197 51135 43231
rect 51077 43191 51135 43197
rect 51261 43231 51319 43237
rect 51261 43197 51273 43231
rect 51307 43228 51319 43231
rect 51626 43228 51632 43240
rect 51307 43200 51632 43228
rect 51307 43197 51319 43200
rect 51261 43191 51319 43197
rect 51092 43160 51120 43191
rect 51626 43188 51632 43200
rect 51684 43188 51690 43240
rect 52086 43228 52092 43240
rect 52047 43200 52092 43228
rect 52086 43188 52092 43200
rect 52144 43188 52150 43240
rect 52729 43231 52787 43237
rect 52729 43197 52741 43231
rect 52775 43197 52787 43231
rect 52729 43191 52787 43197
rect 53009 43231 53067 43237
rect 53009 43197 53021 43231
rect 53055 43228 53067 43231
rect 53834 43228 53840 43240
rect 53055 43200 53840 43228
rect 53055 43197 53067 43200
rect 53009 43191 53067 43197
rect 51534 43160 51540 43172
rect 51092 43132 51540 43160
rect 51534 43120 51540 43132
rect 51592 43120 51598 43172
rect 52748 43160 52776 43191
rect 53834 43188 53840 43200
rect 53892 43188 53898 43240
rect 54202 43228 54208 43240
rect 54163 43200 54208 43228
rect 54202 43188 54208 43200
rect 54260 43188 54266 43240
rect 55033 43231 55091 43237
rect 55033 43197 55045 43231
rect 55079 43197 55091 43231
rect 55033 43191 55091 43197
rect 52914 43160 52920 43172
rect 52748 43132 52920 43160
rect 52914 43120 52920 43132
rect 52972 43120 52978 43172
rect 54018 43120 54024 43172
rect 54076 43160 54082 43172
rect 54478 43160 54484 43172
rect 54076 43132 54484 43160
rect 54076 43120 54082 43132
rect 54478 43120 54484 43132
rect 54536 43160 54542 43172
rect 55048 43160 55076 43191
rect 55122 43188 55128 43240
rect 55180 43228 55186 43240
rect 56060 43228 56088 43268
rect 56965 43265 56977 43268
rect 57011 43265 57023 43299
rect 56965 43259 57023 43265
rect 56873 43231 56931 43237
rect 56873 43228 56885 43231
rect 55180 43200 56088 43228
rect 56428 43200 56885 43228
rect 55180 43188 55186 43200
rect 54536 43132 55076 43160
rect 55300 43163 55358 43169
rect 54536 43120 54542 43132
rect 55300 43129 55312 43163
rect 55346 43160 55358 43163
rect 55858 43160 55864 43172
rect 55346 43132 55864 43160
rect 55346 43129 55358 43132
rect 55300 43123 55358 43129
rect 55858 43120 55864 43132
rect 55916 43120 55922 43172
rect 56428 43104 56456 43200
rect 56873 43197 56885 43200
rect 56919 43197 56931 43231
rect 56873 43191 56931 43197
rect 57974 43160 57980 43172
rect 57935 43132 57980 43160
rect 57974 43120 57980 43132
rect 58032 43120 58038 43172
rect 58158 43160 58164 43172
rect 58119 43132 58164 43160
rect 58158 43120 58164 43132
rect 58216 43120 58222 43172
rect 51166 43092 51172 43104
rect 51127 43064 51172 43092
rect 51166 43052 51172 43064
rect 51224 43052 51230 43104
rect 51442 43052 51448 43104
rect 51500 43092 51506 43104
rect 52549 43095 52607 43101
rect 52549 43092 52561 43095
rect 51500 43064 52561 43092
rect 51500 43052 51506 43064
rect 52549 43061 52561 43064
rect 52595 43061 52607 43095
rect 56410 43092 56416 43104
rect 56371 43064 56416 43092
rect 52549 43055 52607 43061
rect 56410 43052 56416 43064
rect 56468 43052 56474 43104
rect 1104 43002 58880 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 58880 43002
rect 1104 42928 58880 42950
rect 50341 42891 50399 42897
rect 50341 42857 50353 42891
rect 50387 42888 50399 42891
rect 50614 42888 50620 42900
rect 50387 42860 50620 42888
rect 50387 42857 50399 42860
rect 50341 42851 50399 42857
rect 50614 42848 50620 42860
rect 50672 42848 50678 42900
rect 51626 42888 51632 42900
rect 51587 42860 51632 42888
rect 51626 42848 51632 42860
rect 51684 42848 51690 42900
rect 52086 42848 52092 42900
rect 52144 42888 52150 42900
rect 52144 42860 57560 42888
rect 52144 42848 52150 42860
rect 50522 42780 50528 42832
rect 50580 42820 50586 42832
rect 51166 42820 51172 42832
rect 50580 42792 51172 42820
rect 50580 42780 50586 42792
rect 51166 42780 51172 42792
rect 51224 42820 51230 42832
rect 51445 42823 51503 42829
rect 51445 42820 51457 42823
rect 51224 42792 51457 42820
rect 51224 42780 51230 42792
rect 51445 42789 51457 42792
rect 51491 42789 51503 42823
rect 51445 42783 51503 42789
rect 52822 42780 52828 42832
rect 52880 42820 52886 42832
rect 54202 42820 54208 42832
rect 52880 42792 53144 42820
rect 52880 42780 52886 42792
rect 1394 42752 1400 42764
rect 1355 42724 1400 42752
rect 1394 42712 1400 42724
rect 1452 42712 1458 42764
rect 49228 42755 49286 42761
rect 49228 42721 49240 42755
rect 49274 42752 49286 42755
rect 50982 42752 50988 42764
rect 49274 42724 50988 42752
rect 49274 42721 49286 42724
rect 49228 42715 49286 42721
rect 50982 42712 50988 42724
rect 51040 42712 51046 42764
rect 51534 42712 51540 42764
rect 51592 42752 51598 42764
rect 51721 42755 51779 42761
rect 51721 42752 51733 42755
rect 51592 42724 51733 42752
rect 51592 42712 51598 42724
rect 51721 42721 51733 42724
rect 51767 42721 51779 42755
rect 52914 42752 52920 42764
rect 52875 42724 52920 42752
rect 51721 42715 51779 42721
rect 52914 42712 52920 42724
rect 52972 42712 52978 42764
rect 53116 42761 53144 42792
rect 53668 42792 54208 42820
rect 53009 42755 53067 42761
rect 53009 42721 53021 42755
rect 53055 42721 53067 42755
rect 53009 42715 53067 42721
rect 53101 42755 53159 42761
rect 53101 42721 53113 42755
rect 53147 42721 53159 42755
rect 53101 42715 53159 42721
rect 53285 42755 53343 42761
rect 53285 42721 53297 42755
rect 53331 42752 53343 42755
rect 53668 42752 53696 42792
rect 54202 42780 54208 42792
rect 54260 42780 54266 42832
rect 56410 42820 56416 42832
rect 54956 42792 56416 42820
rect 53331 42724 53696 42752
rect 53745 42755 53803 42761
rect 53331 42721 53343 42724
rect 53285 42715 53343 42721
rect 53745 42721 53757 42755
rect 53791 42752 53803 42755
rect 53926 42752 53932 42764
rect 53791 42724 53932 42752
rect 53791 42721 53803 42724
rect 53745 42715 53803 42721
rect 48961 42687 49019 42693
rect 48961 42653 48973 42687
rect 49007 42653 49019 42687
rect 48961 42647 49019 42653
rect 48976 42548 49004 42647
rect 52730 42576 52736 42628
rect 52788 42616 52794 42628
rect 53024 42616 53052 42715
rect 53926 42712 53932 42724
rect 53984 42712 53990 42764
rect 54665 42755 54723 42761
rect 54665 42721 54677 42755
rect 54711 42721 54723 42755
rect 54665 42715 54723 42721
rect 54757 42755 54815 42761
rect 54757 42721 54769 42755
rect 54803 42752 54815 42755
rect 54956 42752 54984 42792
rect 56410 42780 56416 42792
rect 56468 42780 56474 42832
rect 54803 42724 54984 42752
rect 54803 42721 54815 42724
rect 54757 42715 54815 42721
rect 53834 42684 53840 42696
rect 53795 42656 53840 42684
rect 53834 42644 53840 42656
rect 53892 42644 53898 42696
rect 54680 42684 54708 42715
rect 55030 42712 55036 42764
rect 55088 42752 55094 42764
rect 55493 42755 55551 42761
rect 55088 42724 55133 42752
rect 55088 42712 55094 42724
rect 55493 42721 55505 42755
rect 55539 42721 55551 42755
rect 55493 42715 55551 42721
rect 56873 42755 56931 42761
rect 56873 42721 56885 42755
rect 56919 42752 56931 42755
rect 57146 42752 57152 42764
rect 56919 42724 57152 42752
rect 56919 42721 56931 42724
rect 56873 42715 56931 42721
rect 55398 42684 55404 42696
rect 54680 42656 55404 42684
rect 55398 42644 55404 42656
rect 55456 42684 55462 42696
rect 55508 42684 55536 42715
rect 57146 42712 57152 42724
rect 57204 42712 57210 42764
rect 57532 42761 57560 42860
rect 57974 42848 57980 42900
rect 58032 42888 58038 42900
rect 58161 42891 58219 42897
rect 58161 42888 58173 42891
rect 58032 42860 58173 42888
rect 58032 42848 58038 42860
rect 58161 42857 58173 42860
rect 58207 42857 58219 42891
rect 58161 42851 58219 42857
rect 57517 42755 57575 42761
rect 57517 42721 57529 42755
rect 57563 42721 57575 42755
rect 57517 42715 57575 42721
rect 57698 42684 57704 42696
rect 55456 42656 55536 42684
rect 57659 42656 57704 42684
rect 55456 42644 55462 42656
rect 57698 42644 57704 42656
rect 57756 42644 57762 42696
rect 54481 42619 54539 42625
rect 54481 42616 54493 42619
rect 52788 42588 54493 42616
rect 52788 42576 52794 42588
rect 54481 42585 54493 42588
rect 54527 42585 54539 42619
rect 54481 42579 54539 42585
rect 55030 42576 55036 42628
rect 55088 42616 55094 42628
rect 55585 42619 55643 42625
rect 55585 42616 55597 42619
rect 55088 42588 55597 42616
rect 55088 42576 55094 42588
rect 55585 42585 55597 42588
rect 55631 42585 55643 42619
rect 55585 42579 55643 42585
rect 51074 42548 51080 42560
rect 48976 42520 51080 42548
rect 51074 42508 51080 42520
rect 51132 42508 51138 42560
rect 51166 42508 51172 42560
rect 51224 42548 51230 42560
rect 51445 42551 51503 42557
rect 51445 42548 51457 42551
rect 51224 42520 51457 42548
rect 51224 42508 51230 42520
rect 51445 42517 51457 42520
rect 51491 42548 51503 42551
rect 51626 42548 51632 42560
rect 51491 42520 51632 42548
rect 51491 42517 51503 42520
rect 51445 42511 51503 42517
rect 51626 42508 51632 42520
rect 51684 42508 51690 42560
rect 52641 42551 52699 42557
rect 52641 42517 52653 42551
rect 52687 42548 52699 42551
rect 54110 42548 54116 42560
rect 52687 42520 54116 42548
rect 52687 42517 52699 42520
rect 52641 42511 52699 42517
rect 54110 42508 54116 42520
rect 54168 42508 54174 42560
rect 54941 42551 54999 42557
rect 54941 42517 54953 42551
rect 54987 42548 54999 42551
rect 55122 42548 55128 42560
rect 54987 42520 55128 42548
rect 54987 42517 54999 42520
rect 54941 42511 54999 42517
rect 55122 42508 55128 42520
rect 55180 42508 55186 42560
rect 56962 42548 56968 42560
rect 56923 42520 56968 42548
rect 56962 42508 56968 42520
rect 57020 42508 57026 42560
rect 1104 42458 58880 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 58880 42458
rect 1104 42384 58880 42406
rect 50982 42344 50988 42356
rect 50943 42316 50988 42344
rect 50982 42304 50988 42316
rect 51040 42304 51046 42356
rect 52825 42347 52883 42353
rect 52825 42313 52837 42347
rect 52871 42344 52883 42347
rect 54202 42344 54208 42356
rect 52871 42316 54208 42344
rect 52871 42313 52883 42316
rect 52825 42307 52883 42313
rect 54202 42304 54208 42316
rect 54260 42304 54266 42356
rect 55398 42344 55404 42356
rect 55359 42316 55404 42344
rect 55398 42304 55404 42316
rect 55456 42304 55462 42356
rect 55858 42344 55864 42356
rect 55819 42316 55864 42344
rect 55858 42304 55864 42316
rect 55916 42304 55922 42356
rect 57146 42344 57152 42356
rect 57107 42316 57152 42344
rect 57146 42304 57152 42316
rect 57204 42304 57210 42356
rect 50430 42276 50436 42288
rect 50391 42248 50436 42276
rect 50430 42236 50436 42248
rect 50488 42236 50494 42288
rect 52178 42276 52184 42288
rect 52139 42248 52184 42276
rect 52178 42236 52184 42248
rect 52236 42236 52242 42288
rect 50522 42168 50528 42220
rect 50580 42208 50586 42220
rect 50580 42180 50625 42208
rect 50580 42168 50586 42180
rect 55030 42168 55036 42220
rect 55088 42208 55094 42220
rect 55088 42180 56088 42208
rect 55088 42168 55094 42180
rect 49418 42140 49424 42152
rect 49379 42112 49424 42140
rect 49418 42100 49424 42112
rect 49476 42100 49482 42152
rect 50249 42143 50307 42149
rect 50249 42109 50261 42143
rect 50295 42109 50307 42143
rect 50249 42103 50307 42109
rect 50065 42007 50123 42013
rect 50065 41973 50077 42007
rect 50111 42004 50123 42007
rect 50154 42004 50160 42016
rect 50111 41976 50160 42004
rect 50111 41973 50123 41976
rect 50065 41967 50123 41973
rect 50154 41964 50160 41976
rect 50212 41964 50218 42016
rect 50264 42004 50292 42103
rect 51166 42100 51172 42152
rect 51224 42149 51230 42152
rect 51224 42143 51273 42149
rect 51224 42109 51227 42143
rect 51261 42109 51273 42143
rect 51224 42103 51273 42109
rect 51224 42100 51230 42103
rect 51331 42100 51337 42152
rect 51389 42149 51395 42152
rect 51389 42143 51408 42149
rect 51396 42109 51408 42143
rect 51389 42103 51408 42109
rect 51466 42143 51524 42149
rect 51466 42109 51478 42143
rect 51512 42140 51524 42143
rect 51641 42143 51699 42149
rect 51512 42112 51580 42140
rect 51512 42109 51524 42112
rect 51466 42103 51524 42109
rect 51389 42100 51395 42103
rect 51552 42072 51580 42112
rect 51641 42109 51653 42143
rect 51687 42140 51699 42143
rect 52086 42140 52092 42152
rect 51687 42112 52092 42140
rect 51687 42109 51699 42112
rect 51641 42103 51699 42109
rect 52086 42100 52092 42112
rect 52144 42100 52150 42152
rect 52730 42140 52736 42152
rect 52691 42112 52736 42140
rect 52730 42100 52736 42112
rect 52788 42100 52794 42152
rect 52914 42140 52920 42152
rect 52875 42112 52920 42140
rect 52914 42100 52920 42112
rect 52972 42100 52978 42152
rect 54018 42140 54024 42152
rect 53979 42112 54024 42140
rect 54018 42100 54024 42112
rect 54076 42100 54082 42152
rect 54110 42100 54116 42152
rect 54168 42140 54174 42152
rect 54277 42143 54335 42149
rect 54277 42140 54289 42143
rect 54168 42112 54289 42140
rect 54168 42100 54174 42112
rect 54277 42109 54289 42112
rect 54323 42109 54335 42143
rect 54277 42103 54335 42109
rect 54846 42100 54852 42152
rect 54904 42140 54910 42152
rect 56060 42149 56088 42180
rect 55861 42143 55919 42149
rect 55861 42140 55873 42143
rect 54904 42112 55873 42140
rect 54904 42100 54910 42112
rect 55861 42109 55873 42112
rect 55907 42109 55919 42143
rect 55861 42103 55919 42109
rect 56045 42143 56103 42149
rect 56045 42109 56057 42143
rect 56091 42109 56103 42143
rect 56045 42103 56103 42109
rect 56134 42100 56140 42152
rect 56192 42140 56198 42152
rect 56781 42143 56839 42149
rect 56781 42140 56793 42143
rect 56192 42112 56793 42140
rect 56192 42100 56198 42112
rect 56781 42109 56793 42112
rect 56827 42109 56839 42143
rect 56781 42103 56839 42109
rect 56965 42143 57023 42149
rect 56965 42109 56977 42143
rect 57011 42109 57023 42143
rect 56965 42103 57023 42109
rect 52822 42072 52828 42084
rect 51552 42044 52828 42072
rect 51552 42004 51580 42044
rect 52822 42032 52828 42044
rect 52880 42032 52886 42084
rect 55398 42032 55404 42084
rect 55456 42072 55462 42084
rect 56980 42072 57008 42103
rect 57974 42072 57980 42084
rect 55456 42044 57008 42072
rect 57935 42044 57980 42072
rect 55456 42032 55462 42044
rect 57974 42032 57980 42044
rect 58032 42032 58038 42084
rect 58158 42072 58164 42084
rect 58119 42044 58164 42072
rect 58158 42032 58164 42044
rect 58216 42032 58222 42084
rect 50264 41976 51580 42004
rect 1104 41914 58880 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 58880 41914
rect 1104 41840 58880 41862
rect 51629 41803 51687 41809
rect 51629 41769 51641 41803
rect 51675 41800 51687 41803
rect 52086 41800 52092 41812
rect 51675 41772 52092 41800
rect 51675 41769 51687 41772
rect 51629 41763 51687 41769
rect 52086 41760 52092 41772
rect 52144 41760 52150 41812
rect 52549 41803 52607 41809
rect 52549 41769 52561 41803
rect 52595 41800 52607 41803
rect 55398 41800 55404 41812
rect 52595 41772 55404 41800
rect 52595 41769 52607 41772
rect 52549 41763 52607 41769
rect 55398 41760 55404 41772
rect 55456 41760 55462 41812
rect 55585 41803 55643 41809
rect 55585 41769 55597 41803
rect 55631 41800 55643 41803
rect 57698 41800 57704 41812
rect 55631 41772 57704 41800
rect 55631 41769 55643 41772
rect 55585 41763 55643 41769
rect 57698 41760 57704 41772
rect 57756 41760 57762 41812
rect 57974 41760 57980 41812
rect 58032 41800 58038 41812
rect 58161 41803 58219 41809
rect 58161 41800 58173 41803
rect 58032 41772 58173 41800
rect 58032 41760 58038 41772
rect 58161 41769 58173 41772
rect 58207 41769 58219 41803
rect 58161 41763 58219 41769
rect 53392 41704 54248 41732
rect 53392 41676 53420 41704
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 50062 41624 50068 41676
rect 50120 41664 50126 41676
rect 50341 41667 50399 41673
rect 50341 41664 50353 41667
rect 50120 41636 50353 41664
rect 50120 41624 50126 41636
rect 50341 41633 50353 41636
rect 50387 41633 50399 41667
rect 50341 41627 50399 41633
rect 50525 41667 50583 41673
rect 50525 41633 50537 41667
rect 50571 41633 50583 41667
rect 51442 41664 51448 41676
rect 51403 41636 51448 41664
rect 50525 41627 50583 41633
rect 50540 41596 50568 41627
rect 51442 41624 51448 41636
rect 51500 41624 51506 41676
rect 51626 41624 51632 41676
rect 51684 41664 51690 41676
rect 52733 41667 52791 41673
rect 51684 41636 51729 41664
rect 51684 41624 51690 41636
rect 52733 41633 52745 41667
rect 52779 41664 52791 41667
rect 53190 41664 53196 41676
rect 52779 41636 53196 41664
rect 52779 41633 52791 41636
rect 52733 41627 52791 41633
rect 53190 41624 53196 41636
rect 53248 41624 53254 41676
rect 53374 41664 53380 41676
rect 53287 41636 53380 41664
rect 53374 41624 53380 41636
rect 53432 41624 53438 41676
rect 53469 41667 53527 41673
rect 53469 41633 53481 41667
rect 53515 41633 53527 41667
rect 53469 41627 53527 41633
rect 53745 41667 53803 41673
rect 53745 41633 53757 41667
rect 53791 41664 53803 41667
rect 53926 41664 53932 41676
rect 53791 41636 53932 41664
rect 53791 41633 53803 41636
rect 53745 41627 53803 41633
rect 53484 41596 53512 41627
rect 53926 41624 53932 41636
rect 53984 41664 53990 41676
rect 54220 41673 54248 41704
rect 54205 41667 54263 41673
rect 53984 41636 54156 41664
rect 53984 41624 53990 41636
rect 53834 41596 53840 41608
rect 50540 41568 53328 41596
rect 53484 41568 53840 41596
rect 50341 41531 50399 41537
rect 50341 41497 50353 41531
rect 50387 41528 50399 41531
rect 50387 41500 51074 41528
rect 50387 41497 50399 41500
rect 50341 41491 50399 41497
rect 51046 41460 51074 41500
rect 52454 41488 52460 41540
rect 52512 41528 52518 41540
rect 53193 41531 53251 41537
rect 53193 41528 53205 41531
rect 52512 41500 53205 41528
rect 52512 41488 52518 41500
rect 53193 41497 53205 41500
rect 53239 41497 53251 41531
rect 53300 41528 53328 41568
rect 53834 41556 53840 41568
rect 53892 41556 53898 41608
rect 54128 41596 54156 41636
rect 54205 41633 54217 41667
rect 54251 41633 54263 41667
rect 54846 41664 54852 41676
rect 54807 41636 54852 41664
rect 54205 41627 54263 41633
rect 54846 41624 54852 41636
rect 54904 41624 54910 41676
rect 55033 41667 55091 41673
rect 55033 41633 55045 41667
rect 55079 41633 55091 41667
rect 55033 41627 55091 41633
rect 55769 41667 55827 41673
rect 55769 41633 55781 41667
rect 55815 41664 55827 41667
rect 56873 41667 56931 41673
rect 55815 41636 56272 41664
rect 55815 41633 55827 41636
rect 55769 41627 55827 41633
rect 54297 41599 54355 41605
rect 54297 41596 54309 41599
rect 54128 41568 54309 41596
rect 54297 41565 54309 41568
rect 54343 41596 54355 41599
rect 55048 41596 55076 41627
rect 54343 41568 55076 41596
rect 54343 41565 54355 41568
rect 54297 41559 54355 41565
rect 53653 41531 53711 41537
rect 53653 41528 53665 41531
rect 53300 41500 53665 41528
rect 53193 41491 53251 41497
rect 53653 41497 53665 41500
rect 53699 41528 53711 41531
rect 54018 41528 54024 41540
rect 53699 41500 54024 41528
rect 53699 41497 53711 41500
rect 53653 41491 53711 41497
rect 54018 41488 54024 41500
rect 54076 41488 54082 41540
rect 56134 41528 56140 41540
rect 54128 41500 56140 41528
rect 54128 41460 54156 41500
rect 56134 41488 56140 41500
rect 56192 41488 56198 41540
rect 54846 41460 54852 41472
rect 51046 41432 54156 41460
rect 54807 41432 54852 41460
rect 54846 41420 54852 41432
rect 54904 41420 54910 41472
rect 56244 41460 56272 41636
rect 56873 41633 56885 41667
rect 56919 41664 56931 41667
rect 58250 41664 58256 41676
rect 56919 41636 58256 41664
rect 56919 41633 56931 41636
rect 56873 41627 56931 41633
rect 58250 41624 58256 41636
rect 58308 41624 58314 41676
rect 57514 41596 57520 41608
rect 57475 41568 57520 41596
rect 57514 41556 57520 41568
rect 57572 41556 57578 41608
rect 57701 41599 57759 41605
rect 57701 41565 57713 41599
rect 57747 41565 57759 41599
rect 57701 41559 57759 41565
rect 56410 41488 56416 41540
rect 56468 41528 56474 41540
rect 57716 41528 57744 41559
rect 56468 41500 57744 41528
rect 56468 41488 56474 41500
rect 57054 41460 57060 41472
rect 56244 41432 57060 41460
rect 57054 41420 57060 41432
rect 57112 41460 57118 41472
rect 57606 41460 57612 41472
rect 57112 41432 57612 41460
rect 57112 41420 57118 41432
rect 57606 41420 57612 41432
rect 57664 41420 57670 41472
rect 1104 41370 58880 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 58880 41370
rect 1104 41296 58880 41318
rect 50893 41259 50951 41265
rect 50893 41225 50905 41259
rect 50939 41256 50951 41259
rect 52733 41259 52791 41265
rect 50939 41228 52684 41256
rect 50939 41225 50951 41228
rect 50893 41219 50951 41225
rect 51074 41012 51080 41064
rect 51132 41052 51138 41064
rect 51353 41055 51411 41061
rect 51353 41052 51365 41055
rect 51132 41024 51365 41052
rect 51132 41012 51138 41024
rect 51353 41021 51365 41024
rect 51399 41052 51411 41055
rect 51442 41052 51448 41064
rect 51399 41024 51448 41052
rect 51399 41021 51411 41024
rect 51353 41015 51411 41021
rect 51442 41012 51448 41024
rect 51500 41012 51506 41064
rect 50614 40944 50620 40996
rect 50672 40984 50678 40996
rect 51598 40987 51656 40993
rect 51598 40984 51610 40987
rect 50672 40956 51610 40984
rect 50672 40944 50678 40956
rect 51598 40953 51610 40956
rect 51644 40953 51656 40987
rect 52656 40984 52684 41228
rect 52733 41225 52745 41259
rect 52779 41256 52791 41259
rect 53374 41256 53380 41268
rect 52779 41228 53380 41256
rect 52779 41225 52791 41228
rect 52733 41219 52791 41225
rect 53374 41216 53380 41228
rect 53432 41216 53438 41268
rect 53834 41216 53840 41268
rect 53892 41256 53898 41268
rect 55953 41259 56011 41265
rect 55953 41256 55965 41259
rect 53892 41228 55965 41256
rect 53892 41216 53898 41228
rect 55953 41225 55965 41228
rect 55999 41225 56011 41259
rect 55953 41219 56011 41225
rect 54110 41012 54116 41064
rect 54168 41052 54174 41064
rect 54573 41055 54631 41061
rect 54573 41052 54585 41055
rect 54168 41024 54585 41052
rect 54168 41012 54174 41024
rect 54573 41021 54585 41024
rect 54619 41052 54631 41055
rect 54662 41052 54668 41064
rect 54619 41024 54668 41052
rect 54619 41021 54631 41024
rect 54573 41015 54631 41021
rect 54662 41012 54668 41024
rect 54720 41012 54726 41064
rect 54846 41061 54852 41064
rect 54840 41015 54852 41061
rect 54904 41052 54910 41064
rect 55968 41052 55996 41219
rect 56413 41055 56471 41061
rect 56413 41052 56425 41055
rect 54904 41024 54940 41052
rect 55968 41024 56425 41052
rect 54846 41012 54852 41015
rect 54904 41012 54910 41024
rect 56413 41021 56425 41024
rect 56459 41021 56471 41055
rect 57514 41052 57520 41064
rect 56413 41015 56471 41021
rect 56520 41024 57520 41052
rect 56520 40984 56548 41024
rect 57514 41012 57520 41024
rect 57572 41012 57578 41064
rect 57238 40984 57244 40996
rect 52656 40956 56548 40984
rect 57199 40956 57244 40984
rect 51598 40947 51656 40953
rect 57238 40944 57244 40956
rect 57296 40944 57302 40996
rect 57422 40984 57428 40996
rect 57383 40956 57428 40984
rect 57422 40944 57428 40956
rect 57480 40944 57486 40996
rect 57974 40984 57980 40996
rect 57935 40956 57980 40984
rect 57974 40944 57980 40956
rect 58032 40944 58038 40996
rect 53834 40876 53840 40928
rect 53892 40916 53898 40928
rect 54018 40916 54024 40928
rect 53892 40888 54024 40916
rect 53892 40876 53898 40888
rect 54018 40876 54024 40888
rect 54076 40916 54082 40928
rect 56505 40919 56563 40925
rect 56505 40916 56517 40919
rect 54076 40888 56517 40916
rect 54076 40876 54082 40888
rect 56505 40885 56517 40888
rect 56551 40885 56563 40919
rect 56505 40879 56563 40885
rect 57882 40876 57888 40928
rect 57940 40916 57946 40928
rect 58069 40919 58127 40925
rect 58069 40916 58081 40919
rect 57940 40888 58081 40916
rect 57940 40876 57946 40888
rect 58069 40885 58081 40888
rect 58115 40885 58127 40919
rect 58069 40879 58127 40885
rect 1104 40826 58880 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 58880 40826
rect 1104 40752 58880 40774
rect 54481 40715 54539 40721
rect 49712 40684 52040 40712
rect 1394 40576 1400 40588
rect 1355 40548 1400 40576
rect 1394 40536 1400 40548
rect 1452 40536 1458 40588
rect 49712 40585 49740 40684
rect 50433 40647 50491 40653
rect 50433 40613 50445 40647
rect 50479 40644 50491 40647
rect 50614 40644 50620 40656
rect 50479 40616 50620 40644
rect 50479 40613 50491 40616
rect 50433 40607 50491 40613
rect 50614 40604 50620 40616
rect 50672 40604 50678 40656
rect 51902 40644 51908 40656
rect 51644 40616 51908 40644
rect 51644 40585 51672 40616
rect 51902 40604 51908 40616
rect 51960 40604 51966 40656
rect 52012 40644 52040 40684
rect 54481 40681 54493 40715
rect 54527 40712 54539 40715
rect 56410 40712 56416 40724
rect 54527 40684 56416 40712
rect 54527 40681 54539 40684
rect 54481 40675 54539 40681
rect 56410 40672 56416 40684
rect 56468 40672 56474 40724
rect 57974 40672 57980 40724
rect 58032 40712 58038 40724
rect 58161 40715 58219 40721
rect 58161 40712 58173 40715
rect 58032 40684 58173 40712
rect 58032 40672 58038 40684
rect 58161 40681 58173 40684
rect 58207 40681 58219 40715
rect 58161 40675 58219 40681
rect 55214 40644 55220 40656
rect 52012 40616 55220 40644
rect 55214 40604 55220 40616
rect 55272 40604 55278 40656
rect 49697 40579 49755 40585
rect 49697 40545 49709 40579
rect 49743 40545 49755 40579
rect 49697 40539 49755 40545
rect 50341 40579 50399 40585
rect 50341 40545 50353 40579
rect 50387 40545 50399 40579
rect 50341 40539 50399 40545
rect 50525 40579 50583 40585
rect 50525 40545 50537 40579
rect 50571 40576 50583 40579
rect 51629 40579 51687 40585
rect 50571 40548 50660 40576
rect 50571 40545 50583 40548
rect 50525 40539 50583 40545
rect 50356 40440 50384 40539
rect 50632 40520 50660 40548
rect 51629 40545 51641 40579
rect 51675 40545 51687 40579
rect 51629 40539 51687 40545
rect 51997 40579 52055 40585
rect 51997 40545 52009 40579
rect 52043 40576 52055 40579
rect 52454 40576 52460 40588
rect 52043 40548 52460 40576
rect 52043 40545 52055 40548
rect 51997 40539 52055 40545
rect 50614 40468 50620 40520
rect 50672 40468 50678 40520
rect 51445 40511 51503 40517
rect 51445 40477 51457 40511
rect 51491 40508 51503 40511
rect 51810 40508 51816 40520
rect 51491 40480 51816 40508
rect 51491 40477 51503 40480
rect 51445 40471 51503 40477
rect 51810 40468 51816 40480
rect 51868 40508 51874 40520
rect 52012 40508 52040 40539
rect 52454 40536 52460 40548
rect 52512 40536 52518 40588
rect 53009 40579 53067 40585
rect 53009 40545 53021 40579
rect 53055 40545 53067 40579
rect 53466 40576 53472 40588
rect 53427 40548 53472 40576
rect 53009 40539 53067 40545
rect 51868 40480 52040 40508
rect 51868 40468 51874 40480
rect 51721 40443 51779 40449
rect 51721 40440 51733 40443
rect 50356 40412 51733 40440
rect 51721 40409 51733 40412
rect 51767 40409 51779 40443
rect 53024 40440 53052 40539
rect 53466 40536 53472 40548
rect 53524 40536 53530 40588
rect 53834 40576 53840 40588
rect 53795 40548 53840 40576
rect 53834 40536 53840 40548
rect 53892 40536 53898 40588
rect 54665 40579 54723 40585
rect 54665 40545 54677 40579
rect 54711 40545 54723 40579
rect 55122 40576 55128 40588
rect 55083 40548 55128 40576
rect 54665 40539 54723 40545
rect 53558 40508 53564 40520
rect 53519 40480 53564 40508
rect 53558 40468 53564 40480
rect 53616 40468 53622 40520
rect 53745 40511 53803 40517
rect 53745 40477 53757 40511
rect 53791 40508 53803 40511
rect 53926 40508 53932 40520
rect 53791 40480 53932 40508
rect 53791 40477 53803 40480
rect 53745 40471 53803 40477
rect 53926 40468 53932 40480
rect 53984 40508 53990 40520
rect 54294 40508 54300 40520
rect 53984 40480 54300 40508
rect 53984 40468 53990 40480
rect 54294 40468 54300 40480
rect 54352 40468 54358 40520
rect 54680 40508 54708 40539
rect 55122 40536 55128 40548
rect 55180 40536 55186 40588
rect 55309 40579 55367 40585
rect 55309 40545 55321 40579
rect 55355 40576 55367 40579
rect 55490 40576 55496 40588
rect 55355 40548 55496 40576
rect 55355 40545 55367 40548
rect 55309 40539 55367 40545
rect 55490 40536 55496 40548
rect 55548 40536 55554 40588
rect 56594 40536 56600 40588
rect 56652 40576 56658 40588
rect 56689 40579 56747 40585
rect 56689 40576 56701 40579
rect 56652 40548 56701 40576
rect 56652 40536 56658 40548
rect 56689 40545 56701 40548
rect 56735 40545 56747 40579
rect 56689 40539 56747 40545
rect 57054 40508 57060 40520
rect 54680 40480 57060 40508
rect 57054 40468 57060 40480
rect 57112 40468 57118 40520
rect 57146 40468 57152 40520
rect 57204 40508 57210 40520
rect 57517 40511 57575 40517
rect 57517 40508 57529 40511
rect 57204 40480 57529 40508
rect 57204 40468 57210 40480
rect 57517 40477 57529 40480
rect 57563 40477 57575 40511
rect 57517 40471 57575 40477
rect 57606 40468 57612 40520
rect 57664 40508 57670 40520
rect 57701 40511 57759 40517
rect 57701 40508 57713 40511
rect 57664 40480 57713 40508
rect 57664 40468 57670 40480
rect 57701 40477 57713 40480
rect 57747 40477 57759 40511
rect 57701 40471 57759 40477
rect 54018 40440 54024 40452
rect 53024 40412 54024 40440
rect 51721 40403 51779 40409
rect 54018 40400 54024 40412
rect 54076 40400 54082 40452
rect 55030 40400 55036 40452
rect 55088 40440 55094 40452
rect 55582 40440 55588 40452
rect 55088 40412 55588 40440
rect 55088 40400 55094 40412
rect 55582 40400 55588 40412
rect 55640 40440 55646 40452
rect 56781 40443 56839 40449
rect 56781 40440 56793 40443
rect 55640 40412 56793 40440
rect 55640 40400 55646 40412
rect 56781 40409 56793 40412
rect 56827 40409 56839 40443
rect 56781 40403 56839 40409
rect 53098 40372 53104 40384
rect 53059 40344 53104 40372
rect 53098 40332 53104 40344
rect 53156 40332 53162 40384
rect 55125 40375 55183 40381
rect 55125 40341 55137 40375
rect 55171 40372 55183 40375
rect 55398 40372 55404 40384
rect 55171 40344 55404 40372
rect 55171 40341 55183 40344
rect 55125 40335 55183 40341
rect 55398 40332 55404 40344
rect 55456 40332 55462 40384
rect 1104 40282 58880 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 58880 40282
rect 1104 40208 58880 40230
rect 51902 40128 51908 40180
rect 51960 40168 51966 40180
rect 52181 40171 52239 40177
rect 52181 40168 52193 40171
rect 51960 40140 52193 40168
rect 51960 40128 51966 40140
rect 52181 40137 52193 40140
rect 52227 40137 52239 40171
rect 52181 40131 52239 40137
rect 53852 40140 57192 40168
rect 50249 40103 50307 40109
rect 50249 40069 50261 40103
rect 50295 40100 50307 40103
rect 53852 40100 53880 40140
rect 54018 40100 54024 40112
rect 50295 40072 53880 40100
rect 53979 40072 54024 40100
rect 50295 40069 50307 40072
rect 50249 40063 50307 40069
rect 54018 40060 54024 40072
rect 54076 40060 54082 40112
rect 52549 40035 52607 40041
rect 52549 40032 52561 40035
rect 50448 40004 52561 40032
rect 1394 39964 1400 39976
rect 1355 39936 1400 39964
rect 1394 39924 1400 39936
rect 1452 39924 1458 39976
rect 50062 39924 50068 39976
rect 50120 39964 50126 39976
rect 50448 39973 50476 40004
rect 52549 40001 52561 40004
rect 52595 40032 52607 40035
rect 52595 40004 54616 40032
rect 52595 40001 52607 40004
rect 52549 39995 52607 40001
rect 50249 39967 50307 39973
rect 50249 39964 50261 39967
rect 50120 39936 50261 39964
rect 50120 39924 50126 39936
rect 50249 39933 50261 39936
rect 50295 39933 50307 39967
rect 50249 39927 50307 39933
rect 50433 39967 50491 39973
rect 50433 39933 50445 39967
rect 50479 39933 50491 39967
rect 50433 39927 50491 39933
rect 51077 39967 51135 39973
rect 51077 39933 51089 39967
rect 51123 39964 51135 39967
rect 51166 39964 51172 39976
rect 51123 39936 51172 39964
rect 51123 39933 51135 39936
rect 51077 39927 51135 39933
rect 50264 39896 50292 39927
rect 51166 39924 51172 39936
rect 51224 39924 51230 39976
rect 51534 39964 51540 39976
rect 51495 39936 51540 39964
rect 51534 39924 51540 39936
rect 51592 39924 51598 39976
rect 51721 39967 51779 39973
rect 51721 39933 51733 39967
rect 51767 39964 51779 39967
rect 51810 39964 51816 39976
rect 51767 39936 51816 39964
rect 51767 39933 51779 39936
rect 51721 39927 51779 39933
rect 51810 39924 51816 39936
rect 51868 39924 51874 39976
rect 52362 39964 52368 39976
rect 52323 39936 52368 39964
rect 52362 39924 52368 39936
rect 52420 39924 52426 39976
rect 52641 39967 52699 39973
rect 52641 39933 52653 39967
rect 52687 39964 52699 39967
rect 53742 39964 53748 39976
rect 52687 39936 53748 39964
rect 52687 39933 52699 39936
rect 52641 39927 52699 39933
rect 53742 39924 53748 39936
rect 53800 39924 53806 39976
rect 53834 39924 53840 39976
rect 53892 39964 53898 39976
rect 54205 39967 54263 39973
rect 54205 39964 54217 39967
rect 53892 39936 54217 39964
rect 53892 39924 53898 39936
rect 54205 39933 54217 39936
rect 54251 39933 54263 39967
rect 54205 39927 54263 39933
rect 54294 39924 54300 39976
rect 54352 39964 54358 39976
rect 54478 39964 54484 39976
rect 54352 39936 54397 39964
rect 54439 39936 54484 39964
rect 54352 39924 54358 39936
rect 54478 39924 54484 39936
rect 54536 39924 54542 39976
rect 54588 39973 54616 40004
rect 54846 39992 54852 40044
rect 54904 40032 54910 40044
rect 57164 40041 57192 40140
rect 57238 40128 57244 40180
rect 57296 40168 57302 40180
rect 57517 40171 57575 40177
rect 57517 40168 57529 40171
rect 57296 40140 57529 40168
rect 57296 40128 57302 40140
rect 57517 40137 57529 40140
rect 57563 40137 57575 40171
rect 57517 40131 57575 40137
rect 55309 40035 55367 40041
rect 55309 40032 55321 40035
rect 54904 40004 55321 40032
rect 54904 39992 54910 40004
rect 55309 40001 55321 40004
rect 55355 40001 55367 40035
rect 55309 39995 55367 40001
rect 57149 40035 57207 40041
rect 57149 40001 57161 40035
rect 57195 40001 57207 40035
rect 57149 39995 57207 40001
rect 54573 39967 54631 39973
rect 54573 39933 54585 39967
rect 54619 39964 54631 39967
rect 55030 39964 55036 39976
rect 54619 39936 55036 39964
rect 54619 39933 54631 39936
rect 54573 39927 54631 39933
rect 55030 39924 55036 39936
rect 55088 39924 55094 39976
rect 55398 39924 55404 39976
rect 55456 39964 55462 39976
rect 55565 39967 55623 39973
rect 55565 39964 55577 39967
rect 55456 39936 55577 39964
rect 55456 39924 55462 39936
rect 55565 39933 55577 39936
rect 55611 39933 55623 39967
rect 55565 39927 55623 39933
rect 57333 39967 57391 39973
rect 57333 39933 57345 39967
rect 57379 39933 57391 39967
rect 57333 39927 57391 39933
rect 50706 39896 50712 39908
rect 50264 39868 50712 39896
rect 50706 39856 50712 39868
rect 50764 39856 50770 39908
rect 57348 39896 57376 39927
rect 50908 39868 57376 39896
rect 50908 39837 50936 39868
rect 50893 39831 50951 39837
rect 50893 39797 50905 39831
rect 50939 39797 50951 39831
rect 50893 39791 50951 39797
rect 51721 39831 51779 39837
rect 51721 39797 51733 39831
rect 51767 39828 51779 39831
rect 53558 39828 53564 39840
rect 51767 39800 53564 39828
rect 51767 39797 51779 39800
rect 51721 39791 51779 39797
rect 53558 39788 53564 39800
rect 53616 39788 53622 39840
rect 53742 39788 53748 39840
rect 53800 39828 53806 39840
rect 54478 39828 54484 39840
rect 53800 39800 54484 39828
rect 53800 39788 53806 39800
rect 54478 39788 54484 39800
rect 54536 39828 54542 39840
rect 55490 39828 55496 39840
rect 54536 39800 55496 39828
rect 54536 39788 54542 39800
rect 55490 39788 55496 39800
rect 55548 39788 55554 39840
rect 56594 39788 56600 39840
rect 56652 39828 56658 39840
rect 56689 39831 56747 39837
rect 56689 39828 56701 39831
rect 56652 39800 56701 39828
rect 56652 39788 56658 39800
rect 56689 39797 56701 39800
rect 56735 39797 56747 39831
rect 56689 39791 56747 39797
rect 1104 39738 58880 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 58880 39738
rect 1104 39664 58880 39686
rect 51813 39627 51871 39633
rect 51813 39593 51825 39627
rect 51859 39624 51871 39627
rect 52362 39624 52368 39636
rect 51859 39596 52368 39624
rect 51859 39593 51871 39596
rect 51813 39587 51871 39593
rect 52362 39584 52368 39596
rect 52420 39624 52426 39636
rect 53006 39624 53012 39636
rect 52420 39596 53012 39624
rect 52420 39584 52426 39596
rect 53006 39584 53012 39596
rect 53064 39584 53070 39636
rect 53834 39584 53840 39636
rect 53892 39624 53898 39636
rect 54846 39624 54852 39636
rect 53892 39596 54852 39624
rect 53892 39584 53898 39596
rect 54846 39584 54852 39596
rect 54904 39584 54910 39636
rect 55490 39584 55496 39636
rect 55548 39624 55554 39636
rect 55677 39627 55735 39633
rect 55677 39624 55689 39627
rect 55548 39596 55689 39624
rect 55548 39584 55554 39596
rect 55677 39593 55689 39596
rect 55723 39593 55735 39627
rect 55677 39587 55735 39593
rect 51534 39516 51540 39568
rect 51592 39556 51598 39568
rect 52273 39559 52331 39565
rect 51592 39528 51856 39556
rect 51592 39516 51598 39528
rect 51828 39497 51856 39528
rect 52273 39525 52285 39559
rect 52319 39556 52331 39559
rect 53990 39559 54048 39565
rect 53990 39556 54002 39559
rect 52319 39528 54002 39556
rect 52319 39525 52331 39528
rect 52273 39519 52331 39525
rect 53990 39525 54002 39528
rect 54036 39525 54048 39559
rect 55858 39556 55864 39568
rect 53990 39519 54048 39525
rect 54128 39528 55864 39556
rect 51629 39491 51687 39497
rect 51629 39457 51641 39491
rect 51675 39457 51687 39491
rect 51629 39451 51687 39457
rect 51813 39491 51871 39497
rect 51813 39457 51825 39491
rect 51859 39488 51871 39491
rect 52546 39488 52552 39500
rect 51859 39460 52552 39488
rect 51859 39457 51871 39460
rect 51813 39451 51871 39457
rect 51644 39420 51672 39451
rect 52546 39448 52552 39460
rect 52604 39448 52610 39500
rect 52641 39491 52699 39497
rect 52641 39457 52653 39491
rect 52687 39457 52699 39491
rect 52641 39451 52699 39457
rect 52362 39420 52368 39432
rect 51644 39392 52368 39420
rect 52362 39380 52368 39392
rect 52420 39420 52426 39432
rect 52656 39420 52684 39451
rect 52730 39448 52736 39500
rect 52788 39488 52794 39500
rect 52917 39491 52975 39497
rect 52788 39460 52833 39488
rect 52788 39448 52794 39460
rect 52917 39457 52929 39491
rect 52963 39488 52975 39491
rect 53006 39488 53012 39500
rect 52963 39460 53012 39488
rect 52963 39457 52975 39460
rect 52917 39451 52975 39457
rect 53006 39448 53012 39460
rect 53064 39448 53070 39500
rect 54128 39488 54156 39528
rect 55858 39516 55864 39528
rect 55916 39516 55922 39568
rect 53116 39460 54156 39488
rect 55585 39491 55643 39497
rect 52420 39392 52684 39420
rect 52420 39380 52426 39392
rect 51902 39312 51908 39364
rect 51960 39352 51966 39364
rect 53116 39352 53144 39460
rect 55585 39457 55597 39491
rect 55631 39457 55643 39491
rect 55585 39451 55643 39457
rect 56781 39491 56839 39497
rect 56781 39457 56793 39491
rect 56827 39488 56839 39491
rect 58069 39491 58127 39497
rect 58069 39488 58081 39491
rect 56827 39460 58081 39488
rect 56827 39457 56839 39460
rect 56781 39451 56839 39457
rect 58069 39457 58081 39460
rect 58115 39457 58127 39491
rect 58069 39451 58127 39457
rect 53742 39420 53748 39432
rect 53703 39392 53748 39420
rect 53742 39380 53748 39392
rect 53800 39380 53806 39432
rect 51960 39324 53144 39352
rect 51960 39312 51966 39324
rect 55030 39312 55036 39364
rect 55088 39352 55094 39364
rect 55125 39355 55183 39361
rect 55125 39352 55137 39355
rect 55088 39324 55137 39352
rect 55088 39312 55094 39324
rect 55125 39321 55137 39324
rect 55171 39352 55183 39355
rect 55600 39352 55628 39451
rect 56686 39380 56692 39432
rect 56744 39420 56750 39432
rect 57425 39423 57483 39429
rect 57425 39420 57437 39423
rect 56744 39392 57437 39420
rect 56744 39380 56750 39392
rect 57425 39389 57437 39392
rect 57471 39389 57483 39423
rect 57425 39383 57483 39389
rect 57514 39380 57520 39432
rect 57572 39420 57578 39432
rect 57609 39423 57667 39429
rect 57609 39420 57621 39423
rect 57572 39392 57621 39420
rect 57572 39380 57578 39392
rect 57609 39389 57621 39392
rect 57655 39389 57667 39423
rect 57609 39383 57667 39389
rect 56962 39352 56968 39364
rect 55171 39324 55628 39352
rect 56923 39324 56968 39352
rect 55171 39321 55183 39324
rect 55125 39315 55183 39321
rect 56962 39312 56968 39324
rect 57020 39312 57026 39364
rect 50525 39287 50583 39293
rect 50525 39253 50537 39287
rect 50571 39284 50583 39287
rect 57146 39284 57152 39296
rect 50571 39256 57152 39284
rect 50571 39253 50583 39256
rect 50525 39247 50583 39253
rect 57146 39244 57152 39256
rect 57204 39244 57210 39296
rect 1104 39194 58880 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 58880 39194
rect 1104 39120 58880 39142
rect 51166 39040 51172 39092
rect 51224 39080 51230 39092
rect 52089 39083 52147 39089
rect 52089 39080 52101 39083
rect 51224 39052 52101 39080
rect 51224 39040 51230 39052
rect 52089 39049 52101 39052
rect 52135 39049 52147 39083
rect 52089 39043 52147 39049
rect 52362 39040 52368 39092
rect 52420 39080 52426 39092
rect 52549 39083 52607 39089
rect 52549 39080 52561 39083
rect 52420 39052 52561 39080
rect 52420 39040 52426 39052
rect 52549 39049 52561 39052
rect 52595 39049 52607 39083
rect 52549 39043 52607 39049
rect 52638 39040 52644 39092
rect 52696 39080 52702 39092
rect 54849 39083 54907 39089
rect 54849 39080 54861 39083
rect 52696 39052 54861 39080
rect 52696 39040 52702 39052
rect 54849 39049 54861 39052
rect 54895 39049 54907 39083
rect 54849 39043 54907 39049
rect 55309 39083 55367 39089
rect 55309 39049 55321 39083
rect 55355 39080 55367 39083
rect 55582 39080 55588 39092
rect 55355 39052 55588 39080
rect 55355 39049 55367 39052
rect 55309 39043 55367 39049
rect 55582 39040 55588 39052
rect 55640 39040 55646 39092
rect 55214 39012 55220 39024
rect 50632 38984 55220 39012
rect 1394 38876 1400 38888
rect 1355 38848 1400 38876
rect 1394 38836 1400 38848
rect 1452 38836 1458 38888
rect 50632 38885 50660 38984
rect 55214 38972 55220 38984
rect 55272 38972 55278 39024
rect 50706 38904 50712 38956
rect 50764 38944 50770 38956
rect 52546 38944 52552 38956
rect 50764 38916 52552 38944
rect 50764 38904 50770 38916
rect 52546 38904 52552 38916
rect 52604 38904 52610 38956
rect 52638 38904 52644 38956
rect 52696 38944 52702 38956
rect 52825 38947 52883 38953
rect 52825 38944 52837 38947
rect 52696 38916 52837 38944
rect 52696 38904 52702 38916
rect 52825 38913 52837 38916
rect 52871 38913 52883 38947
rect 52825 38907 52883 38913
rect 52917 38947 52975 38953
rect 52917 38913 52929 38947
rect 52963 38944 52975 38947
rect 53190 38944 53196 38956
rect 52963 38916 53196 38944
rect 52963 38913 52975 38916
rect 52917 38907 52975 38913
rect 53190 38904 53196 38916
rect 53248 38904 53254 38956
rect 53282 38904 53288 38956
rect 53340 38944 53346 38956
rect 56689 38947 56747 38953
rect 56689 38944 56701 38947
rect 53340 38916 56701 38944
rect 53340 38904 53346 38916
rect 56689 38913 56701 38916
rect 56735 38913 56747 38947
rect 56689 38907 56747 38913
rect 50617 38879 50675 38885
rect 50617 38845 50629 38879
rect 50663 38845 50675 38879
rect 50617 38839 50675 38845
rect 51166 38836 51172 38888
rect 51224 38876 51230 38888
rect 51445 38879 51503 38885
rect 51445 38876 51457 38879
rect 51224 38848 51457 38876
rect 51224 38836 51230 38848
rect 51445 38845 51457 38848
rect 51491 38845 51503 38879
rect 51902 38876 51908 38888
rect 51863 38848 51908 38876
rect 51445 38839 51503 38845
rect 51902 38836 51908 38848
rect 51960 38836 51966 38888
rect 52454 38836 52460 38888
rect 52512 38876 52518 38888
rect 52733 38879 52791 38885
rect 52733 38876 52745 38879
rect 52512 38848 52745 38876
rect 52512 38836 52518 38848
rect 52733 38845 52745 38848
rect 52779 38845 52791 38879
rect 52733 38839 52791 38845
rect 53006 38836 53012 38888
rect 53064 38876 53070 38888
rect 53064 38848 53109 38876
rect 53064 38836 53070 38848
rect 53558 38836 53564 38888
rect 53616 38876 53622 38888
rect 54021 38879 54079 38885
rect 54021 38876 54033 38879
rect 53616 38848 54033 38876
rect 53616 38836 53622 38848
rect 54021 38845 54033 38848
rect 54067 38845 54079 38879
rect 55030 38876 55036 38888
rect 54991 38848 55036 38876
rect 54021 38839 54079 38845
rect 55030 38836 55036 38848
rect 55088 38836 55094 38888
rect 55125 38879 55183 38885
rect 55125 38845 55137 38879
rect 55171 38845 55183 38879
rect 55125 38839 55183 38845
rect 55401 38879 55459 38885
rect 55401 38845 55413 38879
rect 55447 38876 55459 38879
rect 55490 38876 55496 38888
rect 55447 38848 55496 38876
rect 55447 38845 55459 38848
rect 55401 38839 55459 38845
rect 55140 38808 55168 38839
rect 55490 38836 55496 38848
rect 55548 38836 55554 38888
rect 56226 38836 56232 38888
rect 56284 38876 56290 38888
rect 56413 38879 56471 38885
rect 56413 38876 56425 38879
rect 56284 38848 56425 38876
rect 56284 38836 56290 38848
rect 56413 38845 56425 38848
rect 56459 38845 56471 38879
rect 56413 38839 56471 38845
rect 56594 38808 56600 38820
rect 51276 38780 54984 38808
rect 55140 38780 56600 38808
rect 51276 38749 51304 38780
rect 51261 38743 51319 38749
rect 51261 38709 51273 38743
rect 51307 38709 51319 38743
rect 51261 38703 51319 38709
rect 51994 38700 52000 38752
rect 52052 38740 52058 38752
rect 53190 38740 53196 38752
rect 52052 38712 53196 38740
rect 52052 38700 52058 38712
rect 53190 38700 53196 38712
rect 53248 38700 53254 38752
rect 54110 38740 54116 38752
rect 54071 38712 54116 38740
rect 54110 38700 54116 38712
rect 54168 38700 54174 38752
rect 54956 38740 54984 38780
rect 56594 38768 56600 38780
rect 56652 38768 56658 38820
rect 57698 38768 57704 38820
rect 57756 38808 57762 38820
rect 57977 38811 58035 38817
rect 57977 38808 57989 38811
rect 57756 38780 57989 38808
rect 57756 38768 57762 38780
rect 57977 38777 57989 38780
rect 58023 38777 58035 38811
rect 57977 38771 58035 38777
rect 57514 38740 57520 38752
rect 54956 38712 57520 38740
rect 57514 38700 57520 38712
rect 57572 38700 57578 38752
rect 57882 38700 57888 38752
rect 57940 38740 57946 38752
rect 58069 38743 58127 38749
rect 58069 38740 58081 38743
rect 57940 38712 58081 38740
rect 57940 38700 57946 38712
rect 58069 38709 58081 38712
rect 58115 38709 58127 38743
rect 58069 38703 58127 38709
rect 1104 38650 58880 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 58880 38650
rect 1104 38576 58880 38598
rect 50433 38539 50491 38545
rect 50433 38505 50445 38539
rect 50479 38536 50491 38539
rect 50706 38536 50712 38548
rect 50479 38508 50712 38536
rect 50479 38505 50491 38508
rect 50433 38499 50491 38505
rect 50706 38496 50712 38508
rect 50764 38496 50770 38548
rect 52733 38539 52791 38545
rect 52733 38505 52745 38539
rect 52779 38536 52791 38539
rect 52822 38536 52828 38548
rect 52779 38508 52828 38536
rect 52779 38505 52791 38508
rect 52733 38499 52791 38505
rect 52822 38496 52828 38508
rect 52880 38496 52886 38548
rect 53101 38539 53159 38545
rect 53101 38536 53113 38539
rect 52932 38508 53113 38536
rect 51905 38471 51963 38477
rect 51905 38468 51917 38471
rect 51644 38440 51917 38468
rect 49694 38360 49700 38412
rect 49752 38400 49758 38412
rect 51644 38409 51672 38440
rect 51905 38437 51917 38440
rect 51951 38468 51963 38471
rect 52546 38468 52552 38480
rect 51951 38440 52552 38468
rect 51951 38437 51963 38440
rect 51905 38431 51963 38437
rect 52546 38428 52552 38440
rect 52604 38428 52610 38480
rect 50341 38403 50399 38409
rect 50341 38400 50353 38403
rect 49752 38372 50353 38400
rect 49752 38360 49758 38372
rect 50341 38369 50353 38372
rect 50387 38369 50399 38403
rect 50341 38363 50399 38369
rect 50525 38403 50583 38409
rect 50525 38369 50537 38403
rect 50571 38400 50583 38403
rect 51629 38403 51687 38409
rect 50571 38372 51074 38400
rect 50571 38369 50583 38372
rect 50525 38363 50583 38369
rect 51046 38264 51074 38372
rect 51629 38369 51641 38403
rect 51675 38369 51687 38403
rect 51994 38400 52000 38412
rect 51955 38372 52000 38400
rect 51629 38363 51687 38369
rect 51994 38360 52000 38372
rect 52052 38360 52058 38412
rect 52638 38360 52644 38412
rect 52696 38400 52702 38412
rect 52932 38400 52960 38508
rect 53101 38505 53113 38508
rect 53147 38505 53159 38539
rect 53101 38499 53159 38505
rect 53285 38539 53343 38545
rect 53285 38505 53297 38539
rect 53331 38536 53343 38539
rect 54110 38536 54116 38548
rect 53331 38508 54116 38536
rect 53331 38505 53343 38508
rect 53285 38499 53343 38505
rect 54110 38496 54116 38508
rect 54168 38496 54174 38548
rect 54202 38496 54208 38548
rect 54260 38536 54266 38548
rect 56686 38536 56692 38548
rect 54260 38508 56692 38536
rect 54260 38496 54266 38508
rect 56686 38496 56692 38508
rect 56744 38496 56750 38548
rect 57241 38539 57299 38545
rect 57241 38505 57253 38539
rect 57287 38536 57299 38539
rect 57606 38536 57612 38548
rect 57287 38508 57612 38536
rect 57287 38505 57299 38508
rect 57241 38499 57299 38505
rect 57606 38496 57612 38508
rect 57664 38496 57670 38548
rect 53190 38468 53196 38480
rect 53024 38440 53196 38468
rect 53024 38409 53052 38440
rect 53190 38428 53196 38440
rect 53248 38468 53254 38480
rect 54297 38471 54355 38477
rect 54297 38468 54309 38471
rect 53248 38440 54309 38468
rect 53248 38428 53254 38440
rect 54297 38437 54309 38440
rect 54343 38437 54355 38471
rect 54297 38431 54355 38437
rect 54496 38440 55352 38468
rect 52696 38372 52960 38400
rect 53009 38403 53067 38409
rect 52696 38360 52702 38372
rect 53009 38369 53021 38403
rect 53055 38369 53067 38403
rect 53009 38363 53067 38369
rect 54018 38360 54024 38412
rect 54076 38400 54082 38412
rect 54496 38409 54524 38440
rect 54481 38403 54539 38409
rect 54481 38400 54493 38403
rect 54076 38372 54493 38400
rect 54076 38360 54082 38372
rect 54481 38369 54493 38372
rect 54527 38369 54539 38403
rect 54481 38363 54539 38369
rect 54573 38403 54631 38409
rect 54573 38369 54585 38403
rect 54619 38400 54631 38403
rect 54754 38400 54760 38412
rect 54619 38372 54760 38400
rect 54619 38369 54631 38372
rect 54573 38363 54631 38369
rect 54754 38360 54760 38372
rect 54812 38360 54818 38412
rect 55324 38409 55352 38440
rect 54849 38403 54907 38409
rect 54849 38369 54861 38403
rect 54895 38369 54907 38403
rect 54849 38363 54907 38369
rect 55309 38403 55367 38409
rect 55309 38369 55321 38403
rect 55355 38369 55367 38403
rect 55309 38363 55367 38369
rect 51445 38335 51503 38341
rect 51445 38301 51457 38335
rect 51491 38332 51503 38335
rect 52012 38332 52040 38360
rect 51491 38304 52040 38332
rect 52917 38335 52975 38341
rect 51491 38301 51503 38304
rect 51445 38295 51503 38301
rect 52917 38301 52929 38335
rect 52963 38332 52975 38335
rect 53098 38332 53104 38344
rect 52963 38304 53104 38332
rect 52963 38301 52975 38304
rect 52917 38295 52975 38301
rect 53098 38292 53104 38304
rect 53156 38292 53162 38344
rect 53374 38332 53380 38344
rect 53335 38304 53380 38332
rect 53374 38292 53380 38304
rect 53432 38292 53438 38344
rect 54864 38332 54892 38363
rect 57054 38360 57060 38412
rect 57112 38400 57118 38412
rect 57425 38403 57483 38409
rect 57425 38400 57437 38403
rect 57112 38372 57437 38400
rect 57112 38360 57118 38372
rect 57425 38369 57437 38372
rect 57471 38369 57483 38403
rect 57974 38400 57980 38412
rect 57935 38372 57980 38400
rect 57425 38363 57483 38369
rect 57974 38360 57980 38372
rect 58032 38360 58038 38412
rect 58158 38400 58164 38412
rect 58119 38372 58164 38400
rect 58158 38360 58164 38372
rect 58216 38360 58222 38412
rect 55582 38332 55588 38344
rect 54864 38304 55588 38332
rect 55582 38292 55588 38304
rect 55640 38292 55646 38344
rect 56962 38264 56968 38276
rect 51046 38236 52960 38264
rect 50062 38156 50068 38208
rect 50120 38196 50126 38208
rect 51721 38199 51779 38205
rect 51721 38196 51733 38199
rect 50120 38168 51733 38196
rect 50120 38156 50126 38168
rect 51721 38165 51733 38168
rect 51767 38165 51779 38199
rect 52932 38196 52960 38236
rect 54772 38236 56968 38264
rect 54772 38205 54800 38236
rect 56962 38224 56968 38236
rect 57020 38224 57026 38276
rect 54757 38199 54815 38205
rect 54757 38196 54769 38199
rect 52932 38168 54769 38196
rect 51721 38159 51779 38165
rect 54757 38165 54769 38168
rect 54803 38165 54815 38199
rect 54757 38159 54815 38165
rect 55401 38199 55459 38205
rect 55401 38165 55413 38199
rect 55447 38196 55459 38199
rect 55582 38196 55588 38208
rect 55447 38168 55588 38196
rect 55447 38165 55459 38168
rect 55401 38159 55459 38165
rect 55582 38156 55588 38168
rect 55640 38156 55646 38208
rect 1104 38106 58880 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 58880 38106
rect 1104 38032 58880 38054
rect 49605 37995 49663 38001
rect 49605 37961 49617 37995
rect 49651 37992 49663 37995
rect 53006 37992 53012 38004
rect 49651 37964 52868 37992
rect 52967 37964 53012 37992
rect 49651 37961 49663 37964
rect 49605 37955 49663 37961
rect 52089 37927 52147 37933
rect 52089 37893 52101 37927
rect 52135 37893 52147 37927
rect 52840 37924 52868 37964
rect 53006 37952 53012 37964
rect 53064 37952 53070 38004
rect 53466 37952 53472 38004
rect 53524 37992 53530 38004
rect 54481 37995 54539 38001
rect 54481 37992 54493 37995
rect 53524 37964 54493 37992
rect 53524 37952 53530 37964
rect 54481 37961 54493 37964
rect 54527 37961 54539 37995
rect 57974 37992 57980 38004
rect 54481 37955 54539 37961
rect 55048 37964 57560 37992
rect 57935 37964 57980 37992
rect 55048 37924 55076 37964
rect 56962 37924 56968 37936
rect 52840 37896 55076 37924
rect 56923 37896 56968 37924
rect 52089 37887 52147 37893
rect 52104 37856 52132 37887
rect 56962 37884 56968 37896
rect 57020 37884 57026 37936
rect 54018 37856 54024 37868
rect 52104 37828 54024 37856
rect 54018 37816 54024 37828
rect 54076 37816 54082 37868
rect 54754 37856 54760 37868
rect 54220 37828 54760 37856
rect 1394 37788 1400 37800
rect 1355 37760 1400 37788
rect 1394 37748 1400 37760
rect 1452 37748 1458 37800
rect 50062 37788 50068 37800
rect 50023 37760 50068 37788
rect 50062 37748 50068 37760
rect 50120 37748 50126 37800
rect 50249 37791 50307 37797
rect 50249 37757 50261 37791
rect 50295 37788 50307 37791
rect 50614 37788 50620 37800
rect 50295 37760 50620 37788
rect 50295 37757 50307 37760
rect 50249 37751 50307 37757
rect 50614 37748 50620 37760
rect 50672 37748 50678 37800
rect 50709 37791 50767 37797
rect 50709 37757 50721 37791
rect 50755 37788 50767 37791
rect 51350 37788 51356 37800
rect 50755 37760 51356 37788
rect 50755 37757 50767 37760
rect 50709 37751 50767 37757
rect 51350 37748 51356 37760
rect 51408 37748 51414 37800
rect 52917 37791 52975 37797
rect 52917 37757 52929 37791
rect 52963 37788 52975 37791
rect 53466 37788 53472 37800
rect 52963 37760 53472 37788
rect 52963 37757 52975 37760
rect 52917 37751 52975 37757
rect 53466 37748 53472 37760
rect 53524 37748 53530 37800
rect 50157 37723 50215 37729
rect 50157 37689 50169 37723
rect 50203 37720 50215 37723
rect 50954 37723 51012 37729
rect 50954 37720 50966 37723
rect 50203 37692 50966 37720
rect 50203 37689 50215 37692
rect 50157 37683 50215 37689
rect 50954 37689 50966 37692
rect 51000 37689 51012 37723
rect 54036 37720 54064 37816
rect 54220 37797 54248 37828
rect 54754 37816 54760 37828
rect 54812 37856 54818 37868
rect 57532 37865 57560 37964
rect 57974 37952 57980 37964
rect 58032 37952 58038 38004
rect 57517 37859 57575 37865
rect 54812 37828 55168 37856
rect 54812 37816 54818 37828
rect 54205 37791 54263 37797
rect 54205 37757 54217 37791
rect 54251 37757 54263 37791
rect 54662 37788 54668 37800
rect 54205 37751 54263 37757
rect 54404 37760 54668 37788
rect 54404 37720 54432 37760
rect 54662 37748 54668 37760
rect 54720 37748 54726 37800
rect 54846 37748 54852 37800
rect 54904 37788 54910 37800
rect 55033 37791 55091 37797
rect 55033 37788 55045 37791
rect 54904 37760 55045 37788
rect 54904 37748 54910 37760
rect 55033 37757 55045 37760
rect 55079 37757 55091 37791
rect 55140 37788 55168 37828
rect 57517 37825 57529 37859
rect 57563 37825 57575 37859
rect 57517 37819 57575 37825
rect 56873 37791 56931 37797
rect 55140 37760 56456 37788
rect 55033 37751 55091 37757
rect 50954 37683 51012 37689
rect 51046 37692 52224 37720
rect 54036 37692 54432 37720
rect 54573 37723 54631 37729
rect 49050 37612 49056 37664
rect 49108 37652 49114 37664
rect 51046 37652 51074 37692
rect 49108 37624 51074 37652
rect 52196 37652 52224 37692
rect 54573 37689 54585 37723
rect 54619 37720 54631 37723
rect 54938 37720 54944 37732
rect 54619 37692 54944 37720
rect 54619 37689 54631 37692
rect 54573 37683 54631 37689
rect 54938 37680 54944 37692
rect 54996 37680 55002 37732
rect 55300 37723 55358 37729
rect 55300 37689 55312 37723
rect 55346 37720 55358 37723
rect 55490 37720 55496 37732
rect 55346 37692 55496 37720
rect 55346 37689 55358 37692
rect 55300 37683 55358 37689
rect 55490 37680 55496 37692
rect 55548 37680 55554 37732
rect 55214 37652 55220 37664
rect 52196 37624 55220 37652
rect 49108 37612 49114 37624
rect 55214 37612 55220 37624
rect 55272 37612 55278 37664
rect 56428 37661 56456 37760
rect 56873 37757 56885 37791
rect 56919 37757 56931 37791
rect 56873 37751 56931 37757
rect 56413 37655 56471 37661
rect 56413 37621 56425 37655
rect 56459 37652 56471 37655
rect 56888 37652 56916 37751
rect 57606 37748 57612 37800
rect 57664 37788 57670 37800
rect 57701 37791 57759 37797
rect 57701 37788 57713 37791
rect 57664 37760 57713 37788
rect 57664 37748 57670 37760
rect 57701 37757 57713 37760
rect 57747 37757 57759 37791
rect 57701 37751 57759 37757
rect 56459 37624 56916 37652
rect 56459 37621 56471 37624
rect 56413 37615 56471 37621
rect 1104 37562 58880 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 58880 37562
rect 1104 37488 58880 37510
rect 50341 37451 50399 37457
rect 50341 37417 50353 37451
rect 50387 37448 50399 37451
rect 54938 37448 54944 37460
rect 50387 37420 51074 37448
rect 50387 37417 50399 37420
rect 50341 37411 50399 37417
rect 51046 37380 51074 37420
rect 54312 37420 54800 37448
rect 54899 37420 54944 37448
rect 51046 37352 53880 37380
rect 49050 37312 49056 37324
rect 49011 37284 49056 37312
rect 49050 37272 49056 37284
rect 49108 37272 49114 37324
rect 49694 37312 49700 37324
rect 49655 37284 49700 37312
rect 49694 37272 49700 37284
rect 49752 37272 49758 37324
rect 49881 37315 49939 37321
rect 49881 37281 49893 37315
rect 49927 37312 49939 37315
rect 50525 37315 50583 37321
rect 49927 37284 50476 37312
rect 49927 37281 49939 37284
rect 49881 37275 49939 37281
rect 49786 37244 49792 37256
rect 49747 37216 49792 37244
rect 49786 37204 49792 37216
rect 49844 37204 49850 37256
rect 50448 37244 50476 37284
rect 50525 37281 50537 37315
rect 50571 37312 50583 37315
rect 51166 37312 51172 37324
rect 50571 37284 51172 37312
rect 50571 37281 50583 37284
rect 50525 37275 50583 37281
rect 51166 37272 51172 37284
rect 51224 37272 51230 37324
rect 51902 37312 51908 37324
rect 51863 37284 51908 37312
rect 51902 37272 51908 37284
rect 51960 37272 51966 37324
rect 52086 37312 52092 37324
rect 52047 37284 52092 37312
rect 52086 37272 52092 37284
rect 52144 37272 52150 37324
rect 52454 37272 52460 37324
rect 52512 37312 52518 37324
rect 52805 37315 52863 37321
rect 52805 37312 52817 37315
rect 52512 37284 52817 37312
rect 52512 37272 52518 37284
rect 52805 37281 52817 37284
rect 52851 37281 52863 37315
rect 53852 37312 53880 37352
rect 54312 37312 54340 37420
rect 54662 37380 54668 37392
rect 54623 37352 54668 37380
rect 54662 37340 54668 37352
rect 54720 37340 54726 37392
rect 54772 37380 54800 37420
rect 54938 37408 54944 37420
rect 54996 37408 55002 37460
rect 55490 37448 55496 37460
rect 55451 37420 55496 37448
rect 55490 37408 55496 37420
rect 55548 37408 55554 37460
rect 57698 37448 57704 37460
rect 57659 37420 57704 37448
rect 57698 37408 57704 37420
rect 57756 37408 57762 37460
rect 54772 37352 57284 37380
rect 53852 37284 54340 37312
rect 54389 37315 54447 37321
rect 52805 37275 52863 37281
rect 54389 37281 54401 37315
rect 54435 37281 54447 37315
rect 54570 37312 54576 37324
rect 54531 37284 54576 37312
rect 54389 37275 54447 37281
rect 52362 37244 52368 37256
rect 50448 37216 52368 37244
rect 52362 37204 52368 37216
rect 52420 37204 52426 37256
rect 52549 37247 52607 37253
rect 52549 37244 52561 37247
rect 52472 37216 52561 37244
rect 51994 37176 52000 37188
rect 51955 37148 52000 37176
rect 51994 37136 52000 37148
rect 52052 37136 52058 37188
rect 51350 37068 51356 37120
rect 51408 37108 51414 37120
rect 52472 37108 52500 37216
rect 52549 37213 52561 37216
rect 52595 37213 52607 37247
rect 52549 37207 52607 37213
rect 53834 37204 53840 37256
rect 53892 37244 53898 37256
rect 54404 37244 54432 37275
rect 54570 37272 54576 37284
rect 54628 37272 54634 37324
rect 54754 37272 54760 37324
rect 54812 37312 54818 37324
rect 54812 37284 54857 37312
rect 54812 37272 54818 37284
rect 55122 37272 55128 37324
rect 55180 37312 55186 37324
rect 55401 37315 55459 37321
rect 55401 37312 55413 37315
rect 55180 37284 55413 37312
rect 55180 37272 55186 37284
rect 55401 37281 55413 37284
rect 55447 37281 55459 37315
rect 55582 37312 55588 37324
rect 55543 37284 55588 37312
rect 55401 37275 55459 37281
rect 55582 37272 55588 37284
rect 55640 37272 55646 37324
rect 57256 37321 57284 37352
rect 57241 37315 57299 37321
rect 57241 37281 57253 37315
rect 57287 37281 57299 37315
rect 57241 37275 57299 37281
rect 57054 37244 57060 37256
rect 53892 37216 54432 37244
rect 57015 37216 57060 37244
rect 53892 37204 53898 37216
rect 57054 37204 57060 37216
rect 57112 37204 57118 37256
rect 51408 37080 52500 37108
rect 53929 37111 53987 37117
rect 51408 37068 51414 37080
rect 53929 37077 53941 37111
rect 53975 37108 53987 37111
rect 54018 37108 54024 37120
rect 53975 37080 54024 37108
rect 53975 37077 53987 37080
rect 53929 37071 53987 37077
rect 54018 37068 54024 37080
rect 54076 37108 54082 37120
rect 54570 37108 54576 37120
rect 54076 37080 54576 37108
rect 54076 37068 54082 37080
rect 54570 37068 54576 37080
rect 54628 37068 54634 37120
rect 1104 37018 58880 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 58880 37018
rect 1104 36944 58880 36966
rect 52273 36907 52331 36913
rect 52273 36873 52285 36907
rect 52319 36904 52331 36907
rect 52454 36904 52460 36916
rect 52319 36876 52460 36904
rect 52319 36873 52331 36876
rect 52273 36867 52331 36873
rect 52454 36864 52460 36876
rect 52512 36864 52518 36916
rect 53834 36864 53840 36916
rect 53892 36904 53898 36916
rect 56137 36907 56195 36913
rect 56137 36904 56149 36907
rect 53892 36876 56149 36904
rect 53892 36864 53898 36876
rect 56137 36873 56149 36876
rect 56183 36873 56195 36907
rect 56137 36867 56195 36873
rect 57241 36907 57299 36913
rect 57241 36873 57253 36907
rect 57287 36904 57299 36907
rect 57606 36904 57612 36916
rect 57287 36876 57612 36904
rect 57287 36873 57299 36876
rect 57241 36867 57299 36873
rect 52086 36796 52092 36848
rect 52144 36836 52150 36848
rect 53742 36836 53748 36848
rect 52144 36808 53748 36836
rect 52144 36796 52150 36808
rect 52545 36768 52573 36808
rect 53742 36796 53748 36808
rect 53800 36796 53806 36848
rect 52518 36740 52573 36768
rect 1394 36700 1400 36712
rect 1355 36672 1400 36700
rect 1394 36660 1400 36672
rect 1452 36660 1458 36712
rect 50065 36703 50123 36709
rect 50065 36669 50077 36703
rect 50111 36669 50123 36703
rect 50065 36663 50123 36669
rect 50080 36632 50108 36663
rect 50154 36660 50160 36712
rect 50212 36700 50218 36712
rect 52518 36709 52546 36740
rect 50321 36703 50379 36709
rect 50321 36700 50333 36703
rect 50212 36672 50333 36700
rect 50212 36660 50218 36672
rect 50321 36669 50333 36672
rect 50367 36669 50379 36703
rect 52518 36703 52587 36709
rect 52518 36672 52541 36703
rect 50321 36663 50379 36669
rect 52529 36669 52541 36672
rect 52575 36669 52587 36703
rect 52529 36663 52587 36669
rect 52641 36703 52699 36709
rect 52641 36669 52653 36703
rect 52687 36669 52699 36703
rect 52641 36663 52699 36669
rect 51350 36632 51356 36644
rect 50080 36604 51356 36632
rect 51350 36592 51356 36604
rect 51408 36592 51414 36644
rect 52669 36576 52697 36663
rect 52730 36660 52736 36712
rect 52788 36709 52794 36712
rect 52788 36700 52796 36709
rect 52917 36703 52975 36709
rect 52788 36672 52833 36700
rect 52788 36663 52796 36672
rect 52917 36669 52929 36703
rect 52963 36700 52975 36703
rect 53006 36700 53012 36712
rect 52963 36672 53012 36700
rect 52963 36669 52975 36672
rect 52917 36663 52975 36669
rect 52788 36660 52794 36663
rect 53006 36660 53012 36672
rect 53064 36660 53070 36712
rect 54018 36700 54024 36712
rect 53979 36672 54024 36700
rect 54018 36660 54024 36672
rect 54076 36660 54082 36712
rect 54294 36660 54300 36712
rect 54352 36700 54358 36712
rect 54757 36703 54815 36709
rect 54757 36700 54769 36703
rect 54352 36672 54769 36700
rect 54352 36660 54358 36672
rect 54757 36669 54769 36672
rect 54803 36700 54815 36703
rect 54846 36700 54852 36712
rect 54803 36672 54852 36700
rect 54803 36669 54815 36672
rect 54757 36663 54815 36669
rect 54846 36660 54852 36672
rect 54904 36660 54910 36712
rect 56152 36700 56180 36867
rect 57606 36864 57612 36876
rect 57664 36864 57670 36916
rect 58158 36768 58164 36780
rect 58119 36740 58164 36768
rect 58158 36728 58164 36740
rect 58216 36728 58222 36780
rect 56597 36703 56655 36709
rect 56597 36700 56609 36703
rect 56152 36672 56609 36700
rect 56597 36669 56609 36672
rect 56643 36669 56655 36703
rect 57422 36700 57428 36712
rect 57383 36672 57428 36700
rect 56597 36663 56655 36669
rect 57422 36660 57428 36672
rect 57480 36660 57486 36712
rect 54662 36592 54668 36644
rect 54720 36632 54726 36644
rect 55002 36635 55060 36641
rect 55002 36632 55014 36635
rect 54720 36604 55014 36632
rect 54720 36592 54726 36604
rect 55002 36601 55014 36604
rect 55048 36601 55060 36635
rect 57974 36632 57980 36644
rect 57935 36604 57980 36632
rect 55002 36595 55060 36601
rect 57974 36592 57980 36604
rect 58032 36592 58038 36644
rect 51074 36524 51080 36576
rect 51132 36564 51138 36576
rect 51445 36567 51503 36573
rect 51445 36564 51457 36567
rect 51132 36536 51457 36564
rect 51132 36524 51138 36536
rect 51445 36533 51457 36536
rect 51491 36533 51503 36567
rect 51445 36527 51503 36533
rect 52638 36524 52644 36576
rect 52696 36524 52702 36576
rect 54110 36564 54116 36576
rect 54071 36536 54116 36564
rect 54110 36524 54116 36536
rect 54168 36524 54174 36576
rect 54846 36524 54852 36576
rect 54904 36564 54910 36576
rect 56689 36567 56747 36573
rect 56689 36564 56701 36567
rect 54904 36536 56701 36564
rect 54904 36524 54910 36536
rect 56689 36533 56701 36536
rect 56735 36533 56747 36567
rect 56689 36527 56747 36533
rect 1104 36474 58880 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 58880 36474
rect 1104 36400 58880 36422
rect 52457 36363 52515 36369
rect 52457 36329 52469 36363
rect 52503 36360 52515 36363
rect 52546 36360 52552 36372
rect 52503 36332 52552 36360
rect 52503 36329 52515 36332
rect 52457 36323 52515 36329
rect 52546 36320 52552 36332
rect 52604 36320 52610 36372
rect 52638 36320 52644 36372
rect 52696 36360 52702 36372
rect 53561 36363 53619 36369
rect 53561 36360 53573 36363
rect 52696 36332 53573 36360
rect 52696 36320 52702 36332
rect 53561 36329 53573 36332
rect 53607 36329 53619 36363
rect 54662 36360 54668 36372
rect 54623 36332 54668 36360
rect 53561 36323 53619 36329
rect 54662 36320 54668 36332
rect 54720 36320 54726 36372
rect 56962 36360 56968 36372
rect 56923 36332 56968 36360
rect 56962 36320 56968 36332
rect 57020 36320 57026 36372
rect 57974 36320 57980 36372
rect 58032 36360 58038 36372
rect 58161 36363 58219 36369
rect 58161 36360 58173 36363
rect 58032 36332 58173 36360
rect 58032 36320 58038 36332
rect 58161 36329 58173 36332
rect 58207 36329 58219 36363
rect 58161 36323 58219 36329
rect 51994 36252 52000 36304
rect 52052 36292 52058 36304
rect 53006 36292 53012 36304
rect 52052 36264 53012 36292
rect 52052 36252 52058 36264
rect 1394 36224 1400 36236
rect 1355 36196 1400 36224
rect 1394 36184 1400 36196
rect 1452 36184 1458 36236
rect 51258 36184 51264 36236
rect 51316 36224 51322 36236
rect 52656 36233 52684 36264
rect 53006 36252 53012 36264
rect 53064 36252 53070 36304
rect 54018 36292 54024 36304
rect 53760 36264 54024 36292
rect 53760 36233 53788 36264
rect 54018 36252 54024 36264
rect 54076 36252 54082 36304
rect 55398 36292 55404 36304
rect 54588 36264 55404 36292
rect 51537 36227 51595 36233
rect 51537 36224 51549 36227
rect 51316 36196 51549 36224
rect 51316 36184 51322 36196
rect 51537 36193 51549 36196
rect 51583 36193 51595 36227
rect 51537 36187 51595 36193
rect 52641 36227 52699 36233
rect 52641 36193 52653 36227
rect 52687 36193 52699 36227
rect 52641 36187 52699 36193
rect 53745 36227 53803 36233
rect 53745 36193 53757 36227
rect 53791 36193 53803 36227
rect 53745 36187 53803 36193
rect 53834 36184 53840 36236
rect 53892 36224 53898 36236
rect 54110 36224 54116 36236
rect 53892 36196 53937 36224
rect 54023 36196 54116 36224
rect 53892 36184 53898 36196
rect 54110 36184 54116 36196
rect 54168 36184 54174 36236
rect 54588 36233 54616 36264
rect 55398 36252 55404 36264
rect 55456 36252 55462 36304
rect 54573 36227 54631 36233
rect 54573 36193 54585 36227
rect 54619 36193 54631 36227
rect 54573 36187 54631 36193
rect 54757 36227 54815 36233
rect 54757 36193 54769 36227
rect 54803 36193 54815 36227
rect 55582 36224 55588 36236
rect 55543 36196 55588 36224
rect 54757 36187 54815 36193
rect 52362 36116 52368 36168
rect 52420 36156 52426 36168
rect 52822 36156 52828 36168
rect 52420 36128 52828 36156
rect 52420 36116 52426 36128
rect 52822 36116 52828 36128
rect 52880 36116 52886 36168
rect 52917 36159 52975 36165
rect 52917 36125 52929 36159
rect 52963 36156 52975 36159
rect 54128 36156 54156 36184
rect 54772 36156 54800 36187
rect 55582 36184 55588 36196
rect 55640 36184 55646 36236
rect 56870 36224 56876 36236
rect 56831 36196 56876 36224
rect 56870 36184 56876 36196
rect 56928 36184 56934 36236
rect 56962 36184 56968 36236
rect 57020 36224 57026 36236
rect 57701 36227 57759 36233
rect 57701 36224 57713 36227
rect 57020 36196 57713 36224
rect 57020 36184 57026 36196
rect 57701 36193 57713 36196
rect 57747 36193 57759 36227
rect 57701 36187 57759 36193
rect 52963 36128 54800 36156
rect 57517 36159 57575 36165
rect 52963 36125 52975 36128
rect 52917 36119 52975 36125
rect 57517 36125 57529 36159
rect 57563 36125 57575 36159
rect 57517 36119 57575 36125
rect 50525 36091 50583 36097
rect 50525 36057 50537 36091
rect 50571 36088 50583 36091
rect 57532 36088 57560 36119
rect 50571 36060 57560 36088
rect 50571 36057 50583 36060
rect 50525 36051 50583 36057
rect 51629 36023 51687 36029
rect 51629 35989 51641 36023
rect 51675 36020 51687 36023
rect 52730 36020 52736 36032
rect 51675 35992 52736 36020
rect 51675 35989 51687 35992
rect 51629 35983 51687 35989
rect 52730 35980 52736 35992
rect 52788 35980 52794 36032
rect 52822 35980 52828 36032
rect 52880 36020 52886 36032
rect 54021 36023 54079 36029
rect 54021 36020 54033 36023
rect 52880 35992 54033 36020
rect 52880 35980 52886 35992
rect 54021 35989 54033 35992
rect 54067 36020 54079 36023
rect 54846 36020 54852 36032
rect 54067 35992 54852 36020
rect 54067 35989 54079 35992
rect 54021 35983 54079 35989
rect 54846 35980 54852 35992
rect 54904 35980 54910 36032
rect 54938 35980 54944 36032
rect 54996 36020 55002 36032
rect 55677 36023 55735 36029
rect 55677 36020 55689 36023
rect 54996 35992 55689 36020
rect 54996 35980 55002 35992
rect 55677 35989 55689 35992
rect 55723 35989 55735 36023
rect 55677 35983 55735 35989
rect 1104 35930 58880 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 58880 35930
rect 1104 35856 58880 35878
rect 55214 35816 55220 35828
rect 49712 35788 55220 35816
rect 49712 35621 49740 35788
rect 55214 35776 55220 35788
rect 55272 35776 55278 35828
rect 56870 35776 56876 35828
rect 56928 35816 56934 35828
rect 57241 35819 57299 35825
rect 57241 35816 57253 35819
rect 56928 35788 57253 35816
rect 56928 35776 56934 35788
rect 57241 35785 57253 35788
rect 57287 35785 57299 35819
rect 57241 35779 57299 35785
rect 50341 35751 50399 35757
rect 50341 35717 50353 35751
rect 50387 35748 50399 35751
rect 50387 35720 57100 35748
rect 50387 35717 50399 35720
rect 50341 35711 50399 35717
rect 51166 35680 51172 35692
rect 50540 35652 51172 35680
rect 50540 35621 50568 35652
rect 51166 35640 51172 35652
rect 51224 35640 51230 35692
rect 56962 35680 56968 35692
rect 53024 35652 56968 35680
rect 49697 35615 49755 35621
rect 49697 35581 49709 35615
rect 49743 35581 49755 35615
rect 49697 35575 49755 35581
rect 50525 35615 50583 35621
rect 50525 35581 50537 35615
rect 50571 35581 50583 35615
rect 50525 35575 50583 35581
rect 50890 35572 50896 35624
rect 50948 35612 50954 35624
rect 50985 35615 51043 35621
rect 50985 35612 50997 35615
rect 50948 35584 50997 35612
rect 50948 35572 50954 35584
rect 50985 35581 50997 35584
rect 51031 35581 51043 35615
rect 51718 35612 51724 35624
rect 51679 35584 51724 35612
rect 50985 35575 51043 35581
rect 51718 35572 51724 35584
rect 51776 35572 51782 35624
rect 51905 35615 51963 35621
rect 51905 35581 51917 35615
rect 51951 35612 51963 35615
rect 52086 35612 52092 35624
rect 51951 35584 52092 35612
rect 51951 35581 51963 35584
rect 51905 35575 51963 35581
rect 50614 35504 50620 35556
rect 50672 35544 50678 35556
rect 51920 35544 51948 35575
rect 52086 35572 52092 35584
rect 52144 35572 52150 35624
rect 53024 35612 53052 35652
rect 56962 35640 56968 35652
rect 57020 35640 57026 35692
rect 57072 35689 57100 35720
rect 57057 35683 57115 35689
rect 57057 35649 57069 35683
rect 57103 35649 57115 35683
rect 57057 35643 57115 35649
rect 52932 35584 53052 35612
rect 50672 35516 51948 35544
rect 50672 35504 50678 35516
rect 51077 35479 51135 35485
rect 51077 35445 51089 35479
rect 51123 35476 51135 35479
rect 51258 35476 51264 35488
rect 51123 35448 51264 35476
rect 51123 35445 51135 35448
rect 51077 35439 51135 35445
rect 51258 35436 51264 35448
rect 51316 35436 51322 35488
rect 51810 35476 51816 35488
rect 51771 35448 51816 35476
rect 51810 35436 51816 35448
rect 51868 35436 51874 35488
rect 52932 35485 52960 35584
rect 53098 35572 53104 35624
rect 53156 35612 53162 35624
rect 53156 35584 53201 35612
rect 53156 35572 53162 35584
rect 53926 35572 53932 35624
rect 53984 35612 53990 35624
rect 56873 35615 56931 35621
rect 56873 35612 56885 35615
rect 53984 35584 56885 35612
rect 53984 35572 53990 35584
rect 56873 35581 56885 35584
rect 56919 35581 56931 35615
rect 56873 35575 56931 35581
rect 57977 35615 58035 35621
rect 57977 35581 57989 35615
rect 58023 35612 58035 35615
rect 58066 35612 58072 35624
rect 58023 35584 58072 35612
rect 58023 35581 58035 35584
rect 57977 35575 58035 35581
rect 58066 35572 58072 35584
rect 58124 35612 58130 35624
rect 58342 35612 58348 35624
rect 58124 35584 58348 35612
rect 58124 35572 58130 35584
rect 58342 35572 58348 35584
rect 58400 35572 58406 35624
rect 53006 35504 53012 35556
rect 53064 35544 53070 35556
rect 54481 35547 54539 35553
rect 54481 35544 54493 35547
rect 53064 35516 54493 35544
rect 53064 35504 53070 35516
rect 54481 35513 54493 35516
rect 54527 35544 54539 35547
rect 55217 35547 55275 35553
rect 55217 35544 55229 35547
rect 54527 35516 55229 35544
rect 54527 35513 54539 35516
rect 54481 35507 54539 35513
rect 55217 35513 55229 35516
rect 55263 35513 55275 35547
rect 55398 35544 55404 35556
rect 55359 35516 55404 35544
rect 55217 35507 55275 35513
rect 55398 35504 55404 35516
rect 55456 35504 55462 35556
rect 56226 35544 56232 35556
rect 56187 35516 56232 35544
rect 56226 35504 56232 35516
rect 56284 35544 56290 35556
rect 56686 35544 56692 35556
rect 56284 35516 56692 35544
rect 56284 35504 56290 35516
rect 56686 35504 56692 35516
rect 56744 35504 56750 35556
rect 52917 35479 52975 35485
rect 52917 35445 52929 35479
rect 52963 35445 52975 35479
rect 52917 35439 52975 35445
rect 53098 35436 53104 35488
rect 53156 35476 53162 35488
rect 54386 35476 54392 35488
rect 53156 35448 54392 35476
rect 53156 35436 53162 35448
rect 54386 35436 54392 35448
rect 54444 35436 54450 35488
rect 54573 35479 54631 35485
rect 54573 35445 54585 35479
rect 54619 35476 54631 35479
rect 55122 35476 55128 35488
rect 54619 35448 55128 35476
rect 54619 35445 54631 35448
rect 54573 35439 54631 35445
rect 55122 35436 55128 35448
rect 55180 35436 55186 35488
rect 56318 35476 56324 35488
rect 56279 35448 56324 35476
rect 56318 35436 56324 35448
rect 56376 35436 56382 35488
rect 56594 35436 56600 35488
rect 56652 35476 56658 35488
rect 57422 35476 57428 35488
rect 56652 35448 57428 35476
rect 56652 35436 56658 35448
rect 57422 35436 57428 35448
rect 57480 35476 57486 35488
rect 57882 35476 57888 35488
rect 57480 35448 57888 35476
rect 57480 35436 57486 35448
rect 57882 35436 57888 35448
rect 57940 35476 57946 35488
rect 58161 35479 58219 35485
rect 58161 35476 58173 35479
rect 57940 35448 58173 35476
rect 57940 35436 57946 35448
rect 58161 35445 58173 35448
rect 58207 35445 58219 35479
rect 58161 35439 58219 35445
rect 1104 35386 58880 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 58880 35386
rect 1104 35312 58880 35334
rect 53926 35272 53932 35284
rect 51736 35244 53932 35272
rect 49789 35207 49847 35213
rect 49789 35173 49801 35207
rect 49835 35204 49847 35207
rect 51736 35204 51764 35244
rect 53926 35232 53932 35244
rect 53984 35232 53990 35284
rect 56962 35272 56968 35284
rect 56923 35244 56968 35272
rect 56962 35232 56968 35244
rect 57020 35232 57026 35284
rect 49835 35176 51764 35204
rect 49835 35173 49847 35176
rect 49789 35167 49847 35173
rect 51810 35164 51816 35216
rect 51868 35204 51874 35216
rect 52058 35207 52116 35213
rect 52058 35204 52070 35207
rect 51868 35176 52070 35204
rect 51868 35164 51874 35176
rect 52058 35173 52070 35176
rect 52104 35173 52116 35207
rect 56318 35204 56324 35216
rect 52058 35167 52116 35173
rect 52196 35176 56324 35204
rect 1394 35136 1400 35148
rect 1355 35108 1400 35136
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 49694 35136 49700 35148
rect 49655 35108 49700 35136
rect 49694 35096 49700 35108
rect 49752 35096 49758 35148
rect 49878 35136 49884 35148
rect 49839 35108 49884 35136
rect 49878 35096 49884 35108
rect 49936 35096 49942 35148
rect 50525 35139 50583 35145
rect 50525 35105 50537 35139
rect 50571 35136 50583 35139
rect 51166 35136 51172 35148
rect 50571 35108 51172 35136
rect 50571 35105 50583 35108
rect 50525 35099 50583 35105
rect 51166 35096 51172 35108
rect 51224 35096 51230 35148
rect 52196 35136 52224 35176
rect 56318 35164 56324 35176
rect 56376 35164 56382 35216
rect 51736 35108 52224 35136
rect 53653 35139 53711 35145
rect 49712 35068 49740 35096
rect 50062 35068 50068 35080
rect 49712 35040 50068 35068
rect 50062 35028 50068 35040
rect 50120 35068 50126 35080
rect 51736 35068 51764 35108
rect 53653 35105 53665 35139
rect 53699 35136 53711 35139
rect 54386 35136 54392 35148
rect 53699 35108 54392 35136
rect 53699 35105 53711 35108
rect 53653 35099 53711 35105
rect 50120 35040 51764 35068
rect 51813 35071 51871 35077
rect 50120 35028 50126 35040
rect 51813 35037 51825 35071
rect 51859 35037 51871 35071
rect 51813 35031 51871 35037
rect 50338 35000 50344 35012
rect 50299 34972 50344 35000
rect 50338 34960 50344 34972
rect 50396 34960 50402 35012
rect 51442 34960 51448 35012
rect 51500 35000 51506 35012
rect 51828 35000 51856 35031
rect 53190 35000 53196 35012
rect 51500 34972 51856 35000
rect 53103 34972 53196 35000
rect 51500 34960 51506 34972
rect 53190 34960 53196 34972
rect 53248 35000 53254 35012
rect 53668 35000 53696 35099
rect 54386 35096 54392 35108
rect 54444 35096 54450 35148
rect 54564 35139 54622 35145
rect 54564 35105 54576 35139
rect 54610 35136 54622 35139
rect 55030 35136 55036 35148
rect 54610 35108 55036 35136
rect 54610 35105 54622 35108
rect 54564 35099 54622 35105
rect 55030 35096 55036 35108
rect 55088 35096 55094 35148
rect 56873 35139 56931 35145
rect 56873 35105 56885 35139
rect 56919 35136 56931 35139
rect 58161 35139 58219 35145
rect 58161 35136 58173 35139
rect 56919 35108 58173 35136
rect 56919 35105 56931 35108
rect 56873 35099 56931 35105
rect 58161 35105 58173 35108
rect 58207 35105 58219 35139
rect 58161 35099 58219 35105
rect 53834 35028 53840 35080
rect 53892 35068 53898 35080
rect 54294 35068 54300 35080
rect 53892 35040 54300 35068
rect 53892 35028 53898 35040
rect 54294 35028 54300 35040
rect 54352 35028 54358 35080
rect 57517 35071 57575 35077
rect 57517 35037 57529 35071
rect 57563 35037 57575 35071
rect 57517 35031 57575 35037
rect 57701 35071 57759 35077
rect 57701 35037 57713 35071
rect 57747 35068 57759 35071
rect 58250 35068 58256 35080
rect 57747 35040 58256 35068
rect 57747 35037 57759 35040
rect 57701 35031 57759 35037
rect 57532 35000 57560 35031
rect 58250 35028 58256 35040
rect 58308 35028 58314 35080
rect 53248 34972 53696 35000
rect 55232 34972 57560 35000
rect 53248 34960 53254 34972
rect 50154 34892 50160 34944
rect 50212 34932 50218 34944
rect 53006 34932 53012 34944
rect 50212 34904 53012 34932
rect 50212 34892 50218 34904
rect 53006 34892 53012 34904
rect 53064 34892 53070 34944
rect 53745 34935 53803 34941
rect 53745 34901 53757 34935
rect 53791 34932 53803 34935
rect 54202 34932 54208 34944
rect 53791 34904 54208 34932
rect 53791 34901 53803 34904
rect 53745 34895 53803 34901
rect 54202 34892 54208 34904
rect 54260 34892 54266 34944
rect 54294 34892 54300 34944
rect 54352 34932 54358 34944
rect 55232 34932 55260 34972
rect 54352 34904 55260 34932
rect 54352 34892 54358 34904
rect 55582 34892 55588 34944
rect 55640 34932 55646 34944
rect 55677 34935 55735 34941
rect 55677 34932 55689 34935
rect 55640 34904 55689 34932
rect 55640 34892 55646 34904
rect 55677 34901 55689 34904
rect 55723 34901 55735 34935
rect 55677 34895 55735 34901
rect 1104 34842 58880 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 58880 34842
rect 1104 34768 58880 34790
rect 50154 34688 50160 34740
rect 50212 34728 50218 34740
rect 50341 34731 50399 34737
rect 50341 34728 50353 34731
rect 50212 34700 50353 34728
rect 50212 34688 50218 34700
rect 50341 34697 50353 34700
rect 50387 34697 50399 34731
rect 50341 34691 50399 34697
rect 50890 34688 50896 34740
rect 50948 34728 50954 34740
rect 51261 34731 51319 34737
rect 51261 34728 51273 34731
rect 50948 34700 51273 34728
rect 50948 34688 50954 34700
rect 51261 34697 51273 34700
rect 51307 34697 51319 34731
rect 51261 34691 51319 34697
rect 51718 34688 51724 34740
rect 51776 34728 51782 34740
rect 51997 34731 52055 34737
rect 51997 34728 52009 34731
rect 51776 34700 52009 34728
rect 51776 34688 51782 34700
rect 51997 34697 52009 34700
rect 52043 34697 52055 34731
rect 51997 34691 52055 34697
rect 52086 34688 52092 34740
rect 52144 34728 52150 34740
rect 52917 34731 52975 34737
rect 52917 34728 52929 34731
rect 52144 34700 52929 34728
rect 52144 34688 52150 34700
rect 52917 34697 52929 34700
rect 52963 34697 52975 34731
rect 54294 34728 54300 34740
rect 52917 34691 52975 34697
rect 54128 34700 54300 34728
rect 49697 34663 49755 34669
rect 49697 34629 49709 34663
rect 49743 34660 49755 34663
rect 54128 34660 54156 34700
rect 54294 34688 54300 34700
rect 54352 34688 54358 34740
rect 55030 34728 55036 34740
rect 54991 34700 55036 34728
rect 55030 34688 55036 34700
rect 55088 34688 55094 34740
rect 55122 34688 55128 34740
rect 55180 34728 55186 34740
rect 58069 34731 58127 34737
rect 58069 34728 58081 34731
rect 55180 34700 58081 34728
rect 55180 34688 55186 34700
rect 58069 34697 58081 34700
rect 58115 34697 58127 34731
rect 58069 34691 58127 34697
rect 54938 34660 54944 34672
rect 49743 34632 54156 34660
rect 54404 34632 54944 34660
rect 49743 34629 49755 34632
rect 49697 34623 49755 34629
rect 51721 34595 51779 34601
rect 51721 34561 51733 34595
rect 51767 34592 51779 34595
rect 51767 34564 52316 34592
rect 51767 34561 51779 34564
rect 51721 34555 51779 34561
rect 50157 34527 50215 34533
rect 50157 34493 50169 34527
rect 50203 34524 50215 34527
rect 50982 34524 50988 34536
rect 50203 34496 50988 34524
rect 50203 34493 50215 34496
rect 50157 34487 50215 34493
rect 50982 34484 50988 34496
rect 51040 34484 51046 34536
rect 51902 34524 51908 34536
rect 51863 34496 51908 34524
rect 51902 34484 51908 34496
rect 51960 34484 51966 34536
rect 52288 34533 52316 34564
rect 52273 34527 52331 34533
rect 52273 34493 52285 34527
rect 52319 34524 52331 34527
rect 53558 34524 53564 34536
rect 52319 34496 53564 34524
rect 52319 34493 52331 34496
rect 52273 34487 52331 34493
rect 53558 34484 53564 34496
rect 53616 34524 53622 34536
rect 54021 34527 54079 34533
rect 54021 34524 54033 34527
rect 53616 34496 54033 34524
rect 53616 34484 53622 34496
rect 54021 34493 54033 34496
rect 54067 34493 54079 34527
rect 54202 34524 54208 34536
rect 54163 34496 54208 34524
rect 54021 34487 54079 34493
rect 54202 34484 54208 34496
rect 54260 34484 54266 34536
rect 54297 34527 54355 34533
rect 54297 34493 54309 34527
rect 54343 34524 54355 34527
rect 54404 34524 54432 34632
rect 54938 34620 54944 34632
rect 54996 34620 55002 34672
rect 56410 34660 56416 34672
rect 56371 34632 56416 34660
rect 56410 34620 56416 34632
rect 56468 34620 56474 34672
rect 54481 34595 54539 34601
rect 54481 34561 54493 34595
rect 54527 34592 54539 34595
rect 54662 34592 54668 34604
rect 54527 34564 54668 34592
rect 54527 34561 54539 34564
rect 54481 34555 54539 34561
rect 54662 34552 54668 34564
rect 54720 34552 54726 34604
rect 54846 34552 54852 34604
rect 54904 34592 54910 34604
rect 57054 34592 57060 34604
rect 54904 34564 55260 34592
rect 57015 34564 57060 34592
rect 54904 34552 54910 34564
rect 54570 34524 54576 34536
rect 54343 34496 54432 34524
rect 54531 34496 54576 34524
rect 54343 34493 54355 34496
rect 54297 34487 54355 34493
rect 54570 34484 54576 34496
rect 54628 34484 54634 34536
rect 55232 34533 55260 34564
rect 57054 34552 57060 34564
rect 57112 34552 57118 34604
rect 55033 34527 55091 34533
rect 55033 34524 55045 34527
rect 55017 34493 55045 34524
rect 55079 34493 55091 34527
rect 55017 34487 55091 34493
rect 55229 34527 55287 34533
rect 55229 34493 55241 34527
rect 55275 34493 55287 34527
rect 56870 34524 56876 34536
rect 56831 34496 56876 34524
rect 55229 34487 55287 34493
rect 50798 34416 50804 34468
rect 50856 34456 50862 34468
rect 50893 34459 50951 34465
rect 50893 34456 50905 34459
rect 50856 34428 50905 34456
rect 50856 34416 50862 34428
rect 50893 34425 50905 34428
rect 50939 34425 50951 34459
rect 50893 34419 50951 34425
rect 51074 34416 51080 34468
rect 51132 34456 51138 34468
rect 51920 34456 51948 34484
rect 52181 34459 52239 34465
rect 52181 34456 52193 34459
rect 51132 34428 51177 34456
rect 51920 34428 52193 34456
rect 51132 34416 51138 34428
rect 52181 34425 52193 34428
rect 52227 34425 52239 34459
rect 52181 34419 52239 34425
rect 52362 34416 52368 34468
rect 52420 34456 52426 34468
rect 52825 34459 52883 34465
rect 52825 34456 52837 34459
rect 52420 34428 52837 34456
rect 52420 34416 52426 34428
rect 52825 34425 52837 34428
rect 52871 34425 52883 34459
rect 54220 34456 54248 34484
rect 54846 34456 54852 34468
rect 54220 34428 54852 34456
rect 52825 34419 52883 34425
rect 54846 34416 54852 34428
rect 54904 34416 54910 34468
rect 55017 34456 55045 34487
rect 56870 34484 56876 34496
rect 56928 34484 56934 34536
rect 57517 34527 57575 34533
rect 57517 34524 57529 34527
rect 57164 34496 57529 34524
rect 55398 34456 55404 34468
rect 55017 34428 55404 34456
rect 55398 34416 55404 34428
rect 55456 34456 55462 34468
rect 55950 34456 55956 34468
rect 55456 34428 55956 34456
rect 55456 34416 55462 34428
rect 55950 34416 55956 34428
rect 56008 34416 56014 34468
rect 56229 34459 56287 34465
rect 56229 34425 56241 34459
rect 56275 34456 56287 34459
rect 57164 34456 57192 34496
rect 57517 34493 57529 34496
rect 57563 34493 57575 34527
rect 57974 34524 57980 34536
rect 57935 34496 57980 34524
rect 57517 34487 57575 34493
rect 57974 34484 57980 34496
rect 58032 34484 58038 34536
rect 56275 34428 57192 34456
rect 56275 34425 56287 34428
rect 56229 34419 56287 34425
rect 50706 34348 50712 34400
rect 50764 34388 50770 34400
rect 52730 34388 52736 34400
rect 50764 34360 52736 34388
rect 50764 34348 50770 34360
rect 52730 34348 52736 34360
rect 52788 34348 52794 34400
rect 52914 34348 52920 34400
rect 52972 34388 52978 34400
rect 57146 34388 57152 34400
rect 52972 34360 57152 34388
rect 52972 34348 52978 34360
rect 57146 34348 57152 34360
rect 57204 34348 57210 34400
rect 1104 34298 58880 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 58880 34298
rect 1104 34224 58880 34246
rect 50433 34187 50491 34193
rect 50433 34153 50445 34187
rect 50479 34184 50491 34187
rect 50614 34184 50620 34196
rect 50479 34156 50620 34184
rect 50479 34153 50491 34156
rect 50433 34147 50491 34153
rect 50614 34144 50620 34156
rect 50672 34144 50678 34196
rect 51902 34184 51908 34196
rect 51863 34156 51908 34184
rect 51902 34144 51908 34156
rect 51960 34144 51966 34196
rect 52730 34144 52736 34196
rect 52788 34184 52794 34196
rect 52788 34156 56180 34184
rect 52788 34144 52794 34156
rect 55214 34116 55220 34128
rect 49712 34088 55220 34116
rect 1394 34048 1400 34060
rect 1355 34020 1400 34048
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 49712 34057 49740 34088
rect 55214 34076 55220 34088
rect 55272 34076 55278 34128
rect 49697 34051 49755 34057
rect 49697 34017 49709 34051
rect 49743 34017 49755 34051
rect 49697 34011 49755 34017
rect 50062 34008 50068 34060
rect 50120 34048 50126 34060
rect 50341 34051 50399 34057
rect 50341 34048 50353 34051
rect 50120 34020 50353 34048
rect 50120 34008 50126 34020
rect 50341 34017 50353 34020
rect 50387 34017 50399 34051
rect 50341 34011 50399 34017
rect 50525 34051 50583 34057
rect 50525 34017 50537 34051
rect 50571 34048 50583 34051
rect 52089 34051 52147 34057
rect 50571 34020 51074 34048
rect 50571 34017 50583 34020
rect 50525 34011 50583 34017
rect 51046 33844 51074 34020
rect 52089 34017 52101 34051
rect 52135 34048 52147 34051
rect 52178 34048 52184 34060
rect 52135 34020 52184 34048
rect 52135 34017 52147 34020
rect 52089 34011 52147 34017
rect 52178 34008 52184 34020
rect 52236 34008 52242 34060
rect 53010 34051 53068 34057
rect 53010 34048 53022 34051
rect 52932 34020 53022 34048
rect 52365 33983 52423 33989
rect 52365 33949 52377 33983
rect 52411 33980 52423 33983
rect 52454 33980 52460 33992
rect 52411 33952 52460 33980
rect 52411 33949 52423 33952
rect 52365 33943 52423 33949
rect 52454 33940 52460 33952
rect 52512 33980 52518 33992
rect 52932 33980 52960 34020
rect 53010 34017 53022 34020
rect 53056 34017 53068 34051
rect 53010 34011 53068 34017
rect 53101 34051 53159 34057
rect 53101 34017 53113 34051
rect 53147 34017 53159 34051
rect 53374 34048 53380 34060
rect 53335 34020 53380 34048
rect 53101 34011 53159 34017
rect 52512 33952 52960 33980
rect 53116 33980 53144 34011
rect 53374 34008 53380 34020
rect 53432 34008 53438 34060
rect 54656 34051 54714 34057
rect 54656 34017 54668 34051
rect 54702 34048 54714 34051
rect 56042 34048 56048 34060
rect 54702 34020 56048 34048
rect 54702 34017 54714 34020
rect 54656 34011 54714 34017
rect 56042 34008 56048 34020
rect 56100 34008 56106 34060
rect 56152 34048 56180 34156
rect 56686 34144 56692 34196
rect 56744 34184 56750 34196
rect 56873 34187 56931 34193
rect 56873 34184 56885 34187
rect 56744 34156 56885 34184
rect 56744 34144 56750 34156
rect 56873 34153 56885 34156
rect 56919 34153 56931 34187
rect 56873 34147 56931 34153
rect 56778 34116 56784 34128
rect 56739 34088 56784 34116
rect 56778 34076 56784 34088
rect 56836 34076 56842 34128
rect 57517 34051 57575 34057
rect 57517 34048 57529 34051
rect 56152 34020 57529 34048
rect 57517 34017 57529 34020
rect 57563 34017 57575 34051
rect 57517 34011 57575 34017
rect 53116 33952 53788 33980
rect 52512 33940 52518 33952
rect 52825 33915 52883 33921
rect 52825 33881 52837 33915
rect 52871 33912 52883 33915
rect 53006 33912 53012 33924
rect 52871 33884 53012 33912
rect 52871 33881 52883 33884
rect 52825 33875 52883 33881
rect 53006 33872 53012 33884
rect 53064 33872 53070 33924
rect 52273 33847 52331 33853
rect 52273 33844 52285 33847
rect 51046 33816 52285 33844
rect 52273 33813 52285 33816
rect 52319 33844 52331 33847
rect 53116 33844 53144 33952
rect 53282 33844 53288 33856
rect 52319 33816 53144 33844
rect 53243 33816 53288 33844
rect 52319 33813 52331 33816
rect 52273 33807 52331 33813
rect 53282 33804 53288 33816
rect 53340 33804 53346 33856
rect 53760 33844 53788 33952
rect 53834 33940 53840 33992
rect 53892 33980 53898 33992
rect 54389 33983 54447 33989
rect 54389 33980 54401 33983
rect 53892 33952 54401 33980
rect 53892 33940 53898 33952
rect 54389 33949 54401 33952
rect 54435 33949 54447 33983
rect 54389 33943 54447 33949
rect 57606 33940 57612 33992
rect 57664 33980 57670 33992
rect 57701 33983 57759 33989
rect 57701 33980 57713 33983
rect 57664 33952 57713 33980
rect 57664 33940 57670 33952
rect 57701 33949 57713 33952
rect 57747 33949 57759 33983
rect 57701 33943 57759 33949
rect 57974 33940 57980 33992
rect 58032 33940 58038 33992
rect 55398 33872 55404 33924
rect 55456 33912 55462 33924
rect 55769 33915 55827 33921
rect 55769 33912 55781 33915
rect 55456 33884 55781 33912
rect 55456 33872 55462 33884
rect 55769 33881 55781 33884
rect 55815 33912 55827 33915
rect 57992 33912 58020 33940
rect 55815 33884 58020 33912
rect 55815 33881 55827 33884
rect 55769 33875 55827 33881
rect 55122 33844 55128 33856
rect 53760 33816 55128 33844
rect 55122 33804 55128 33816
rect 55180 33804 55186 33856
rect 57974 33844 57980 33856
rect 57935 33816 57980 33844
rect 57974 33804 57980 33816
rect 58032 33804 58038 33856
rect 1104 33754 58880 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 58880 33754
rect 1104 33680 58880 33702
rect 49789 33643 49847 33649
rect 49789 33609 49801 33643
rect 49835 33640 49847 33643
rect 50706 33640 50712 33652
rect 49835 33612 50712 33640
rect 49835 33609 49847 33612
rect 49789 33603 49847 33609
rect 50706 33600 50712 33612
rect 50764 33600 50770 33652
rect 51997 33643 52055 33649
rect 51997 33609 52009 33643
rect 52043 33640 52055 33643
rect 52454 33640 52460 33652
rect 52043 33612 52460 33640
rect 52043 33609 52055 33612
rect 51997 33603 52055 33609
rect 52454 33600 52460 33612
rect 52512 33640 52518 33652
rect 55493 33643 55551 33649
rect 52512 33612 55444 33640
rect 52512 33600 52518 33612
rect 50249 33575 50307 33581
rect 50249 33541 50261 33575
rect 50295 33572 50307 33575
rect 52914 33572 52920 33584
rect 50295 33544 52920 33572
rect 50295 33541 50307 33544
rect 50249 33535 50307 33541
rect 52914 33532 52920 33544
rect 52972 33532 52978 33584
rect 53101 33575 53159 33581
rect 53101 33541 53113 33575
rect 53147 33572 53159 33575
rect 54386 33572 54392 33584
rect 53147 33544 54392 33572
rect 53147 33541 53159 33544
rect 53101 33535 53159 33541
rect 54386 33532 54392 33544
rect 54444 33532 54450 33584
rect 54481 33575 54539 33581
rect 54481 33541 54493 33575
rect 54527 33572 54539 33575
rect 55416 33572 55444 33612
rect 55493 33609 55505 33643
rect 55539 33640 55551 33643
rect 55582 33640 55588 33652
rect 55539 33612 55588 33640
rect 55539 33609 55551 33612
rect 55493 33603 55551 33609
rect 55582 33600 55588 33612
rect 55640 33600 55646 33652
rect 56042 33640 56048 33652
rect 56003 33612 56048 33640
rect 56042 33600 56048 33612
rect 56100 33600 56106 33652
rect 58158 33572 58164 33584
rect 54527 33544 54699 33572
rect 55416 33544 56272 33572
rect 58119 33544 58164 33572
rect 54527 33541 54539 33544
rect 54481 33535 54539 33541
rect 50890 33464 50896 33516
rect 50948 33504 50954 33516
rect 53374 33504 53380 33516
rect 50948 33476 51028 33504
rect 50948 33464 50954 33476
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 50062 33396 50068 33448
rect 50120 33436 50126 33448
rect 50249 33439 50307 33445
rect 50249 33436 50261 33439
rect 50120 33408 50261 33436
rect 50120 33396 50126 33408
rect 50249 33405 50261 33408
rect 50295 33405 50307 33439
rect 50249 33399 50307 33405
rect 50433 33439 50491 33445
rect 50433 33405 50445 33439
rect 50479 33436 50491 33439
rect 50706 33436 50712 33448
rect 50479 33408 50712 33436
rect 50479 33405 50491 33408
rect 50433 33399 50491 33405
rect 50706 33396 50712 33408
rect 50764 33396 50770 33448
rect 51000 33445 51028 33476
rect 51920 33476 53380 33504
rect 51920 33445 51948 33476
rect 52840 33448 52868 33476
rect 53374 33464 53380 33476
rect 53432 33504 53438 33516
rect 54671 33504 54699 33544
rect 54754 33504 54760 33516
rect 53432 33476 54524 33504
rect 54671 33476 54760 33504
rect 53432 33464 53438 33476
rect 50985 33439 51043 33445
rect 50985 33405 50997 33439
rect 51031 33405 51043 33439
rect 50985 33399 51043 33405
rect 51905 33439 51963 33445
rect 51905 33405 51917 33439
rect 51951 33405 51963 33439
rect 52546 33436 52552 33448
rect 52507 33408 52552 33436
rect 51905 33399 51963 33405
rect 52546 33396 52552 33408
rect 52604 33396 52610 33448
rect 52822 33436 52828 33448
rect 52735 33408 52828 33436
rect 52822 33396 52828 33408
rect 52880 33396 52886 33448
rect 52917 33439 52975 33445
rect 52917 33405 52929 33439
rect 52963 33436 52975 33439
rect 53282 33436 53288 33448
rect 52963 33408 53288 33436
rect 52963 33405 52975 33408
rect 52917 33399 52975 33405
rect 53282 33396 53288 33408
rect 53340 33396 53346 33448
rect 53466 33396 53472 33448
rect 53524 33436 53530 33448
rect 54386 33445 54392 33448
rect 54205 33439 54263 33445
rect 54205 33436 54217 33439
rect 53524 33408 54217 33436
rect 53524 33396 53530 33408
rect 54205 33405 54217 33408
rect 54251 33405 54263 33439
rect 54205 33399 54263 33405
rect 54343 33439 54392 33445
rect 54343 33405 54355 33439
rect 54389 33405 54392 33439
rect 54343 33399 54392 33405
rect 54386 33396 54392 33399
rect 54444 33396 54450 33448
rect 54496 33436 54524 33476
rect 54754 33464 54760 33476
rect 54812 33464 54818 33516
rect 55141 33476 55352 33504
rect 54573 33439 54631 33445
rect 54573 33436 54585 33439
rect 54496 33408 54585 33436
rect 54573 33405 54585 33408
rect 54619 33405 54631 33439
rect 54573 33399 54631 33405
rect 54662 33396 54668 33448
rect 54720 33436 54726 33448
rect 55141 33436 55169 33476
rect 55324 33445 55352 33476
rect 54720 33408 55169 33436
rect 55217 33439 55275 33445
rect 54720 33396 54726 33408
rect 55217 33405 55229 33439
rect 55263 33405 55275 33439
rect 55217 33399 55275 33405
rect 55309 33439 55367 33445
rect 55309 33405 55321 33439
rect 55355 33405 55367 33439
rect 55309 33399 55367 33405
rect 52733 33371 52791 33377
rect 52733 33337 52745 33371
rect 52779 33337 52791 33371
rect 52733 33331 52791 33337
rect 54021 33371 54079 33377
rect 54021 33337 54033 33371
rect 54067 33368 54079 33371
rect 55232 33368 55260 33399
rect 55490 33396 55496 33448
rect 55548 33436 55554 33448
rect 55585 33439 55643 33445
rect 55585 33436 55597 33439
rect 55548 33408 55597 33436
rect 55548 33396 55554 33408
rect 55585 33405 55597 33408
rect 55631 33405 55643 33439
rect 56042 33436 56048 33448
rect 56003 33408 56048 33436
rect 55585 33399 55643 33405
rect 56042 33396 56048 33408
rect 56100 33396 56106 33448
rect 56244 33445 56272 33544
rect 58158 33532 58164 33544
rect 58216 33532 58222 33584
rect 56229 33439 56287 33445
rect 56229 33405 56241 33439
rect 56275 33405 56287 33439
rect 57974 33436 57980 33448
rect 57935 33408 57980 33436
rect 56229 33399 56287 33405
rect 57974 33396 57980 33408
rect 58032 33396 58038 33448
rect 54067 33340 55260 33368
rect 57241 33371 57299 33377
rect 54067 33337 54079 33340
rect 54021 33331 54079 33337
rect 57241 33337 57253 33371
rect 57287 33368 57299 33371
rect 57514 33368 57520 33380
rect 57287 33340 57520 33368
rect 57287 33337 57299 33340
rect 57241 33331 57299 33337
rect 51077 33303 51135 33309
rect 51077 33269 51089 33303
rect 51123 33300 51135 33303
rect 51350 33300 51356 33312
rect 51123 33272 51356 33300
rect 51123 33269 51135 33272
rect 51077 33263 51135 33269
rect 51350 33260 51356 33272
rect 51408 33300 51414 33312
rect 52270 33300 52276 33312
rect 51408 33272 52276 33300
rect 51408 33260 51414 33272
rect 52270 33260 52276 33272
rect 52328 33260 52334 33312
rect 52748 33300 52776 33331
rect 57514 33328 57520 33340
rect 57572 33328 57578 33380
rect 53190 33300 53196 33312
rect 52748 33272 53196 33300
rect 53190 33260 53196 33272
rect 53248 33260 53254 33312
rect 55030 33300 55036 33312
rect 54991 33272 55036 33300
rect 55030 33260 55036 33272
rect 55088 33260 55094 33312
rect 57330 33300 57336 33312
rect 57291 33272 57336 33300
rect 57330 33260 57336 33272
rect 57388 33260 57394 33312
rect 1104 33210 58880 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 58880 33210
rect 1104 33136 58880 33158
rect 52638 33096 52644 33108
rect 50540 33068 52644 33096
rect 49694 32960 49700 32972
rect 49655 32932 49700 32960
rect 49694 32920 49700 32932
rect 49752 32920 49758 32972
rect 50540 32969 50568 33068
rect 52638 33056 52644 33068
rect 52696 33056 52702 33108
rect 52822 33096 52828 33108
rect 52783 33068 52828 33096
rect 52822 33056 52828 33068
rect 52880 33056 52886 33108
rect 53558 33096 53564 33108
rect 53519 33068 53564 33096
rect 53558 33056 53564 33068
rect 53616 33056 53622 33108
rect 54294 33056 54300 33108
rect 54352 33096 54358 33108
rect 55122 33096 55128 33108
rect 54352 33068 55128 33096
rect 54352 33056 54358 33068
rect 55122 33056 55128 33068
rect 55180 33096 55186 33108
rect 55180 33068 55536 33096
rect 55180 33056 55186 33068
rect 52362 32988 52368 33040
rect 52420 33028 52426 33040
rect 53469 33031 53527 33037
rect 53469 33028 53481 33031
rect 52420 33000 53481 33028
rect 52420 32988 52426 33000
rect 53469 32997 53481 33000
rect 53515 32997 53527 33031
rect 53469 32991 53527 32997
rect 54110 32988 54116 33040
rect 54168 33028 54174 33040
rect 54168 33000 55260 33028
rect 54168 32988 54174 33000
rect 50525 32963 50583 32969
rect 50525 32929 50537 32963
rect 50571 32929 50583 32963
rect 50525 32923 50583 32929
rect 51534 32920 51540 32972
rect 51592 32960 51598 32972
rect 51701 32963 51759 32969
rect 51701 32960 51713 32963
rect 51592 32932 51713 32960
rect 51592 32920 51598 32932
rect 51701 32929 51713 32932
rect 51747 32929 51759 32963
rect 53650 32960 53656 32972
rect 53611 32932 53656 32960
rect 51701 32923 51759 32929
rect 53650 32920 53656 32932
rect 53708 32920 53714 32972
rect 54294 32960 54300 32972
rect 54255 32932 54300 32960
rect 54294 32920 54300 32932
rect 54352 32920 54358 32972
rect 55232 32969 55260 33000
rect 55508 32969 55536 33068
rect 55125 32963 55183 32969
rect 55125 32929 55137 32963
rect 55171 32929 55183 32963
rect 55125 32923 55183 32929
rect 55217 32963 55275 32969
rect 55217 32929 55229 32963
rect 55263 32929 55275 32963
rect 55217 32923 55275 32929
rect 55493 32963 55551 32969
rect 55493 32929 55505 32963
rect 55539 32929 55551 32963
rect 57146 32960 57152 32972
rect 57107 32932 57152 32960
rect 55493 32923 55551 32929
rect 51445 32895 51503 32901
rect 51445 32892 51457 32895
rect 51046 32864 51457 32892
rect 49510 32784 49516 32836
rect 49568 32824 49574 32836
rect 51046 32824 51074 32864
rect 51445 32861 51457 32864
rect 51491 32861 51503 32895
rect 51445 32855 51503 32861
rect 54389 32895 54447 32901
rect 54389 32861 54401 32895
rect 54435 32892 54447 32895
rect 55140 32892 55168 32923
rect 57146 32920 57152 32932
rect 57204 32920 57210 32972
rect 57330 32892 57336 32904
rect 54435 32864 55168 32892
rect 57291 32864 57336 32892
rect 54435 32861 54447 32864
rect 54389 32855 54447 32861
rect 49568 32796 51074 32824
rect 49568 32784 49574 32796
rect 52546 32784 52552 32836
rect 52604 32824 52610 32836
rect 53285 32827 53343 32833
rect 53285 32824 53297 32827
rect 52604 32796 53297 32824
rect 52604 32784 52610 32796
rect 53285 32793 53297 32796
rect 53331 32824 53343 32827
rect 54018 32824 54024 32836
rect 53331 32796 54024 32824
rect 53331 32793 53343 32796
rect 53285 32787 53343 32793
rect 54018 32784 54024 32796
rect 54076 32824 54082 32836
rect 54478 32824 54484 32836
rect 54076 32796 54484 32824
rect 54076 32784 54082 32796
rect 54478 32784 54484 32796
rect 54536 32784 54542 32836
rect 54754 32784 54760 32836
rect 54812 32824 54818 32836
rect 54941 32827 54999 32833
rect 54941 32824 54953 32827
rect 54812 32796 54953 32824
rect 54812 32784 54818 32796
rect 54941 32793 54953 32796
rect 54987 32793 54999 32827
rect 55140 32824 55168 32864
rect 57330 32852 57336 32864
rect 57388 32852 57394 32904
rect 55490 32824 55496 32836
rect 55140 32796 55496 32824
rect 54941 32787 54999 32793
rect 55490 32784 55496 32796
rect 55548 32784 55554 32836
rect 57514 32824 57520 32836
rect 57475 32796 57520 32824
rect 57514 32784 57520 32796
rect 57572 32784 57578 32836
rect 50341 32759 50399 32765
rect 50341 32725 50353 32759
rect 50387 32756 50399 32759
rect 52730 32756 52736 32768
rect 50387 32728 52736 32756
rect 50387 32725 50399 32728
rect 50341 32719 50399 32725
rect 52730 32716 52736 32728
rect 52788 32716 52794 32768
rect 53837 32759 53895 32765
rect 53837 32725 53849 32759
rect 53883 32756 53895 32759
rect 54294 32756 54300 32768
rect 53883 32728 54300 32756
rect 53883 32725 53895 32728
rect 53837 32719 53895 32725
rect 54294 32716 54300 32728
rect 54352 32716 54358 32768
rect 54846 32716 54852 32768
rect 54904 32756 54910 32768
rect 55401 32759 55459 32765
rect 55401 32756 55413 32759
rect 54904 32728 55413 32756
rect 54904 32716 54910 32728
rect 55401 32725 55413 32728
rect 55447 32756 55459 32759
rect 56594 32756 56600 32768
rect 55447 32728 56600 32756
rect 55447 32725 55459 32728
rect 55401 32719 55459 32725
rect 56594 32716 56600 32728
rect 56652 32716 56658 32768
rect 1104 32666 58880 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 58880 32666
rect 1104 32592 58880 32614
rect 51534 32552 51540 32564
rect 51495 32524 51540 32552
rect 51534 32512 51540 32524
rect 51592 32512 51598 32564
rect 52730 32512 52736 32564
rect 52788 32552 52794 32564
rect 52788 32524 57744 32552
rect 52788 32512 52794 32524
rect 50985 32487 51043 32493
rect 50985 32453 50997 32487
rect 51031 32484 51043 32487
rect 52178 32484 52184 32496
rect 51031 32456 52184 32484
rect 51031 32453 51043 32456
rect 50985 32447 51043 32453
rect 52178 32444 52184 32456
rect 52236 32444 52242 32496
rect 52825 32487 52883 32493
rect 52825 32453 52837 32487
rect 52871 32484 52883 32487
rect 54938 32484 54944 32496
rect 52871 32456 54944 32484
rect 52871 32453 52883 32456
rect 52825 32447 52883 32453
rect 54938 32444 54944 32456
rect 54996 32444 55002 32496
rect 56594 32444 56600 32496
rect 56652 32484 56658 32496
rect 56689 32487 56747 32493
rect 56689 32484 56701 32487
rect 56652 32456 56701 32484
rect 56652 32444 56658 32456
rect 56689 32453 56701 32456
rect 56735 32453 56747 32487
rect 56689 32447 56747 32453
rect 53006 32416 53012 32428
rect 51828 32388 53012 32416
rect 1394 32348 1400 32360
rect 1355 32320 1400 32348
rect 1394 32308 1400 32320
rect 1452 32308 1458 32360
rect 51828 32357 51856 32388
rect 53006 32376 53012 32388
rect 53064 32416 53070 32428
rect 53650 32416 53656 32428
rect 53064 32388 53656 32416
rect 53064 32376 53070 32388
rect 53650 32376 53656 32388
rect 53708 32376 53714 32428
rect 53742 32376 53748 32428
rect 53800 32416 53806 32428
rect 54021 32419 54079 32425
rect 54021 32416 54033 32419
rect 53800 32388 54033 32416
rect 53800 32376 53806 32388
rect 54021 32385 54033 32388
rect 54067 32385 54079 32419
rect 54294 32416 54300 32428
rect 54255 32388 54300 32416
rect 54021 32379 54079 32385
rect 54294 32376 54300 32388
rect 54352 32376 54358 32428
rect 54481 32419 54539 32425
rect 54481 32385 54493 32419
rect 54527 32416 54539 32419
rect 55030 32416 55036 32428
rect 54527 32388 55036 32416
rect 54527 32385 54539 32388
rect 54481 32379 54539 32385
rect 55030 32376 55036 32388
rect 55088 32376 55094 32428
rect 57716 32425 57744 32524
rect 57701 32419 57759 32425
rect 57701 32385 57713 32419
rect 57747 32385 57759 32419
rect 57701 32379 57759 32385
rect 50893 32351 50951 32357
rect 50893 32317 50905 32351
rect 50939 32317 50951 32351
rect 50893 32311 50951 32317
rect 51077 32351 51135 32357
rect 51077 32317 51089 32351
rect 51123 32348 51135 32351
rect 51813 32351 51871 32357
rect 51813 32348 51825 32351
rect 51123 32320 51825 32348
rect 51123 32317 51135 32320
rect 51077 32311 51135 32317
rect 51813 32317 51825 32320
rect 51859 32317 51871 32351
rect 51813 32311 51871 32317
rect 51905 32351 51963 32357
rect 51905 32317 51917 32351
rect 51951 32317 51963 32351
rect 51905 32311 51963 32317
rect 50908 32280 50936 32311
rect 51718 32280 51724 32292
rect 50908 32252 51724 32280
rect 51718 32240 51724 32252
rect 51776 32280 51782 32292
rect 51920 32280 51948 32311
rect 51994 32308 52000 32360
rect 52052 32348 52058 32360
rect 52178 32348 52184 32360
rect 52052 32320 52097 32348
rect 52139 32320 52184 32348
rect 52052 32308 52058 32320
rect 52178 32308 52184 32320
rect 52236 32308 52242 32360
rect 52825 32351 52883 32357
rect 52825 32317 52837 32351
rect 52871 32348 52883 32351
rect 52917 32351 52975 32357
rect 52917 32348 52929 32351
rect 52871 32320 52929 32348
rect 52871 32317 52883 32320
rect 52825 32311 52883 32317
rect 52917 32317 52929 32320
rect 52963 32317 52975 32351
rect 52917 32311 52975 32317
rect 53282 32308 53288 32360
rect 53340 32348 53346 32360
rect 54205 32351 54263 32357
rect 54205 32348 54217 32351
rect 53340 32320 54217 32348
rect 53340 32308 53346 32320
rect 54205 32317 54217 32320
rect 54251 32317 54263 32351
rect 54205 32311 54263 32317
rect 54389 32351 54447 32357
rect 54389 32317 54401 32351
rect 54435 32317 54447 32351
rect 54389 32311 54447 32317
rect 55309 32351 55367 32357
rect 55309 32317 55321 32351
rect 55355 32348 55367 32351
rect 55950 32348 55956 32360
rect 55355 32320 55956 32348
rect 55355 32317 55367 32320
rect 55309 32311 55367 32317
rect 51776 32252 51948 32280
rect 51776 32240 51782 32252
rect 52270 32240 52276 32292
rect 52328 32280 52334 32292
rect 54404 32280 54432 32311
rect 55950 32308 55956 32320
rect 56008 32308 56014 32360
rect 57517 32351 57575 32357
rect 57517 32317 57529 32351
rect 57563 32317 57575 32351
rect 57517 32311 57575 32317
rect 52328 32252 54432 32280
rect 52328 32240 52334 32252
rect 55398 32240 55404 32292
rect 55456 32280 55462 32292
rect 55554 32283 55612 32289
rect 55554 32280 55566 32283
rect 55456 32252 55566 32280
rect 55456 32240 55462 32252
rect 55554 32249 55566 32252
rect 55600 32249 55612 32283
rect 55554 32243 55612 32249
rect 50706 32172 50712 32224
rect 50764 32212 50770 32224
rect 53009 32215 53067 32221
rect 53009 32212 53021 32215
rect 50764 32184 53021 32212
rect 50764 32172 50770 32184
rect 53009 32181 53021 32184
rect 53055 32212 53067 32215
rect 54110 32212 54116 32224
rect 53055 32184 54116 32212
rect 53055 32181 53067 32184
rect 53009 32175 53067 32181
rect 54110 32172 54116 32184
rect 54168 32172 54174 32224
rect 54294 32172 54300 32224
rect 54352 32212 54358 32224
rect 57532 32212 57560 32311
rect 54352 32184 57560 32212
rect 54352 32172 54358 32184
rect 57974 32172 57980 32224
rect 58032 32212 58038 32224
rect 58161 32215 58219 32221
rect 58161 32212 58173 32215
rect 58032 32184 58173 32212
rect 58032 32172 58038 32184
rect 58161 32181 58173 32184
rect 58207 32181 58219 32215
rect 58161 32175 58219 32181
rect 1104 32122 58880 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 58880 32122
rect 1104 32048 58880 32070
rect 51718 32008 51724 32020
rect 51679 31980 51724 32008
rect 51718 31968 51724 31980
rect 51776 31968 51782 32020
rect 54113 32011 54171 32017
rect 51920 31980 52132 32008
rect 51920 31940 51948 31980
rect 50540 31912 51948 31940
rect 52104 31940 52132 31980
rect 54113 31977 54125 32011
rect 54159 32008 54171 32011
rect 54478 32008 54484 32020
rect 54159 31980 54484 32008
rect 54159 31977 54171 31980
rect 54113 31971 54171 31977
rect 54478 31968 54484 31980
rect 54536 32008 54542 32020
rect 54536 31980 55076 32008
rect 54536 31968 54542 31980
rect 54294 31940 54300 31952
rect 52104 31912 54300 31940
rect 48314 31832 48320 31884
rect 48372 31872 48378 31884
rect 50540 31881 50568 31912
rect 54294 31900 54300 31912
rect 54352 31900 54358 31952
rect 55048 31949 55076 31980
rect 55033 31943 55091 31949
rect 55033 31909 55045 31943
rect 55079 31909 55091 31943
rect 55033 31903 55091 31909
rect 55122 31900 55128 31952
rect 55180 31940 55186 31952
rect 57974 31940 57980 31952
rect 55180 31912 55225 31940
rect 57935 31912 57980 31940
rect 55180 31900 55186 31912
rect 57974 31900 57980 31912
rect 58032 31900 58038 31952
rect 58158 31940 58164 31952
rect 58119 31912 58164 31940
rect 58158 31900 58164 31912
rect 58216 31900 58222 31952
rect 49881 31875 49939 31881
rect 49881 31872 49893 31875
rect 48372 31844 49893 31872
rect 48372 31832 48378 31844
rect 49881 31841 49893 31844
rect 49927 31841 49939 31875
rect 49881 31835 49939 31841
rect 50525 31875 50583 31881
rect 50525 31841 50537 31875
rect 50571 31841 50583 31875
rect 51810 31872 51816 31884
rect 50525 31835 50583 31841
rect 51046 31844 51816 31872
rect 51046 31804 51074 31844
rect 51810 31832 51816 31844
rect 51868 31832 51874 31884
rect 51997 31875 52055 31881
rect 51997 31841 52009 31875
rect 52043 31872 52055 31875
rect 52362 31872 52368 31884
rect 52043 31844 52368 31872
rect 52043 31841 52055 31844
rect 51997 31835 52055 31841
rect 52362 31832 52368 31844
rect 52420 31832 52426 31884
rect 52454 31832 52460 31884
rect 52512 31872 52518 31884
rect 52989 31875 53047 31881
rect 52989 31872 53001 31875
rect 52512 31844 53001 31872
rect 52512 31832 52518 31844
rect 52989 31841 53001 31844
rect 53035 31841 53047 31875
rect 52989 31835 53047 31841
rect 54570 31832 54576 31884
rect 54628 31872 54634 31884
rect 54849 31875 54907 31881
rect 54849 31872 54861 31875
rect 54628 31844 54861 31872
rect 54628 31832 54634 31844
rect 54849 31841 54861 31844
rect 54895 31841 54907 31875
rect 54849 31835 54907 31841
rect 54938 31832 54944 31884
rect 54996 31872 55002 31884
rect 55217 31875 55275 31881
rect 55217 31872 55229 31875
rect 54996 31844 55229 31872
rect 54996 31832 55002 31844
rect 55217 31841 55229 31844
rect 55263 31841 55275 31875
rect 55217 31835 55275 31841
rect 57241 31875 57299 31881
rect 57241 31841 57253 31875
rect 57287 31872 57299 31875
rect 58066 31872 58072 31884
rect 57287 31844 58072 31872
rect 57287 31841 57299 31844
rect 57241 31835 57299 31841
rect 58066 31832 58072 31844
rect 58124 31832 58130 31884
rect 51902 31804 51908 31816
rect 49712 31776 51074 31804
rect 51863 31776 51908 31804
rect 49712 31745 49740 31776
rect 51902 31764 51908 31776
rect 51960 31764 51966 31816
rect 52089 31807 52147 31813
rect 52089 31773 52101 31807
rect 52135 31773 52147 31807
rect 52089 31767 52147 31773
rect 52181 31807 52239 31813
rect 52181 31773 52193 31807
rect 52227 31804 52239 31807
rect 52227 31776 52684 31804
rect 52227 31773 52239 31776
rect 52181 31767 52239 31773
rect 49697 31739 49755 31745
rect 49697 31705 49709 31739
rect 49743 31736 49755 31739
rect 52104 31736 52132 31767
rect 52546 31736 52552 31748
rect 49743 31708 49777 31736
rect 52104 31708 52552 31736
rect 49743 31705 49755 31708
rect 49697 31699 49755 31705
rect 52546 31696 52552 31708
rect 52604 31696 52610 31748
rect 52178 31628 52184 31680
rect 52236 31668 52242 31680
rect 52454 31668 52460 31680
rect 52236 31640 52460 31668
rect 52236 31628 52242 31640
rect 52454 31628 52460 31640
rect 52512 31628 52518 31680
rect 52656 31668 52684 31776
rect 52730 31764 52736 31816
rect 52788 31804 52794 31816
rect 57422 31804 57428 31816
rect 52788 31776 52833 31804
rect 57383 31776 57428 31804
rect 52788 31764 52794 31776
rect 57422 31764 57428 31776
rect 57480 31764 57486 31816
rect 54570 31696 54576 31748
rect 54628 31736 54634 31748
rect 56410 31736 56416 31748
rect 54628 31708 56416 31736
rect 54628 31696 54634 31708
rect 56410 31696 56416 31708
rect 56468 31696 56474 31748
rect 54386 31668 54392 31680
rect 52656 31640 54392 31668
rect 54386 31628 54392 31640
rect 54444 31628 54450 31680
rect 54662 31628 54668 31680
rect 54720 31668 54726 31680
rect 55401 31671 55459 31677
rect 55401 31668 55413 31671
rect 54720 31640 55413 31668
rect 54720 31628 54726 31640
rect 55401 31637 55413 31640
rect 55447 31637 55459 31671
rect 55401 31631 55459 31637
rect 1104 31578 58880 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 58880 31578
rect 1104 31504 58880 31526
rect 50801 31467 50859 31473
rect 50801 31433 50813 31467
rect 50847 31464 50859 31467
rect 51258 31464 51264 31476
rect 50847 31436 51264 31464
rect 50847 31433 50859 31436
rect 50801 31427 50859 31433
rect 51258 31424 51264 31436
rect 51316 31424 51322 31476
rect 51442 31464 51448 31476
rect 51355 31436 51448 31464
rect 51442 31424 51448 31436
rect 51500 31464 51506 31476
rect 52730 31464 52736 31476
rect 51500 31436 52736 31464
rect 51500 31424 51506 31436
rect 52730 31424 52736 31436
rect 52788 31424 52794 31476
rect 54386 31464 54392 31476
rect 54347 31436 54392 31464
rect 54386 31424 54392 31436
rect 54444 31424 54450 31476
rect 54754 31464 54760 31476
rect 54715 31436 54760 31464
rect 54754 31424 54760 31436
rect 54812 31424 54818 31476
rect 57330 31464 57336 31476
rect 55140 31436 57336 31464
rect 49329 31399 49387 31405
rect 49329 31365 49341 31399
rect 49375 31396 49387 31399
rect 51460 31396 51488 31424
rect 49375 31368 51488 31396
rect 49375 31365 49387 31368
rect 49329 31359 49387 31365
rect 51534 31356 51540 31408
rect 51592 31396 51598 31408
rect 51994 31396 52000 31408
rect 51592 31368 52000 31396
rect 51592 31356 51598 31368
rect 51994 31356 52000 31368
rect 52052 31356 52058 31408
rect 52917 31399 52975 31405
rect 52917 31365 52929 31399
rect 52963 31396 52975 31399
rect 55140 31396 55168 31436
rect 57330 31424 57336 31436
rect 57388 31424 57394 31476
rect 58066 31464 58072 31476
rect 58027 31436 58072 31464
rect 58066 31424 58072 31436
rect 58124 31424 58130 31476
rect 52963 31368 55168 31396
rect 52963 31365 52975 31368
rect 52917 31359 52975 31365
rect 49988 31300 54524 31328
rect 1394 31260 1400 31272
rect 1355 31232 1400 31260
rect 1394 31220 1400 31232
rect 1452 31220 1458 31272
rect 48866 31220 48872 31272
rect 48924 31260 48930 31272
rect 49988 31269 50016 31300
rect 49513 31263 49571 31269
rect 49513 31260 49525 31263
rect 48924 31232 49525 31260
rect 48924 31220 48930 31232
rect 49513 31229 49525 31232
rect 49559 31229 49571 31263
rect 49513 31223 49571 31229
rect 49973 31263 50031 31269
rect 49973 31229 49985 31263
rect 50019 31229 50031 31263
rect 49973 31223 50031 31229
rect 51994 31220 52000 31272
rect 52052 31260 52058 31272
rect 52273 31263 52331 31269
rect 52273 31260 52285 31263
rect 52052 31232 52285 31260
rect 52052 31220 52058 31232
rect 52273 31229 52285 31232
rect 52319 31229 52331 31263
rect 52273 31223 52331 31229
rect 52362 31220 52368 31272
rect 52420 31260 52426 31272
rect 52457 31263 52515 31269
rect 52457 31260 52469 31263
rect 52420 31232 52469 31260
rect 52420 31220 52426 31232
rect 52457 31229 52469 31232
rect 52503 31229 52515 31263
rect 52457 31223 52515 31229
rect 53101 31263 53159 31269
rect 53101 31229 53113 31263
rect 53147 31229 53159 31263
rect 53101 31223 53159 31229
rect 51166 31152 51172 31204
rect 51224 31192 51230 31204
rect 51353 31195 51411 31201
rect 51353 31192 51365 31195
rect 51224 31164 51365 31192
rect 51224 31152 51230 31164
rect 51353 31161 51365 31164
rect 51399 31192 51411 31195
rect 51399 31164 51672 31192
rect 51399 31161 51411 31164
rect 51353 31155 51411 31161
rect 51445 31127 51503 31133
rect 51445 31093 51457 31127
rect 51491 31124 51503 31127
rect 51534 31124 51540 31136
rect 51491 31096 51540 31124
rect 51491 31093 51503 31096
rect 51445 31087 51503 31093
rect 51534 31084 51540 31096
rect 51592 31084 51598 31136
rect 51644 31124 51672 31164
rect 51718 31152 51724 31204
rect 51776 31192 51782 31204
rect 53116 31192 53144 31223
rect 51776 31164 53144 31192
rect 54496 31192 54524 31300
rect 54573 31263 54631 31269
rect 54573 31229 54585 31263
rect 54619 31260 54631 31263
rect 54662 31260 54668 31272
rect 54619 31232 54668 31260
rect 54619 31229 54631 31232
rect 54573 31223 54631 31229
rect 54662 31220 54668 31232
rect 54720 31220 54726 31272
rect 54846 31260 54852 31272
rect 54807 31232 54852 31260
rect 54846 31220 54852 31232
rect 54904 31220 54910 31272
rect 54938 31220 54944 31272
rect 54996 31260 55002 31272
rect 55309 31263 55367 31269
rect 55309 31260 55321 31263
rect 54996 31232 55321 31260
rect 54996 31220 55002 31232
rect 55309 31229 55321 31232
rect 55355 31260 55367 31263
rect 55950 31260 55956 31272
rect 55355 31232 55956 31260
rect 55355 31229 55367 31232
rect 55309 31223 55367 31229
rect 55950 31220 55956 31232
rect 56008 31220 56014 31272
rect 57422 31260 57428 31272
rect 57383 31232 57428 31260
rect 57422 31220 57428 31232
rect 57480 31220 57486 31272
rect 57609 31263 57667 31269
rect 57609 31229 57621 31263
rect 57655 31229 57667 31263
rect 57609 31223 57667 31229
rect 55214 31192 55220 31204
rect 54496 31164 55220 31192
rect 51776 31152 51782 31164
rect 55214 31152 55220 31164
rect 55272 31152 55278 31204
rect 55576 31195 55634 31201
rect 55576 31161 55588 31195
rect 55622 31192 55634 31195
rect 55674 31192 55680 31204
rect 55622 31164 55680 31192
rect 55622 31161 55634 31164
rect 55576 31155 55634 31161
rect 55674 31152 55680 31164
rect 55732 31152 55738 31204
rect 57624 31192 57652 31223
rect 55784 31164 57652 31192
rect 52086 31124 52092 31136
rect 51644 31096 52092 31124
rect 52086 31084 52092 31096
rect 52144 31084 52150 31136
rect 52457 31127 52515 31133
rect 52457 31093 52469 31127
rect 52503 31124 52515 31127
rect 52822 31124 52828 31136
rect 52503 31096 52828 31124
rect 52503 31093 52515 31096
rect 52457 31087 52515 31093
rect 52822 31084 52828 31096
rect 52880 31084 52886 31136
rect 52914 31084 52920 31136
rect 52972 31124 52978 31136
rect 55784 31124 55812 31164
rect 52972 31096 55812 31124
rect 52972 31084 52978 31096
rect 56410 31084 56416 31136
rect 56468 31124 56474 31136
rect 56689 31127 56747 31133
rect 56689 31124 56701 31127
rect 56468 31096 56701 31124
rect 56468 31084 56474 31096
rect 56689 31093 56701 31096
rect 56735 31093 56747 31127
rect 56689 31087 56747 31093
rect 1104 31034 58880 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 58880 31034
rect 1104 30960 58880 30982
rect 50433 30923 50491 30929
rect 50433 30889 50445 30923
rect 50479 30920 50491 30923
rect 50706 30920 50712 30932
rect 50479 30892 50712 30920
rect 50479 30889 50491 30892
rect 50433 30883 50491 30889
rect 50706 30880 50712 30892
rect 50764 30880 50770 30932
rect 52178 30920 52184 30932
rect 52139 30892 52184 30920
rect 52178 30880 52184 30892
rect 52236 30880 52242 30932
rect 52362 30880 52368 30932
rect 52420 30920 52426 30932
rect 54297 30923 54355 30929
rect 54297 30920 54309 30923
rect 52420 30892 54309 30920
rect 52420 30880 52426 30892
rect 54297 30889 54309 30892
rect 54343 30889 54355 30923
rect 55398 30920 55404 30932
rect 55359 30892 55404 30920
rect 54297 30883 54355 30889
rect 55398 30880 55404 30892
rect 55456 30880 55462 30932
rect 49050 30812 49056 30864
rect 49108 30852 49114 30864
rect 49108 30824 50384 30852
rect 49108 30812 49114 30824
rect 1394 30784 1400 30796
rect 1355 30756 1400 30784
rect 1394 30744 1400 30756
rect 1452 30744 1458 30796
rect 50356 30793 50384 30824
rect 51994 30812 52000 30864
rect 52052 30852 52058 30864
rect 52052 30824 52546 30852
rect 52052 30812 52058 30824
rect 49697 30787 49755 30793
rect 49697 30753 49709 30787
rect 49743 30753 49755 30787
rect 49697 30747 49755 30753
rect 50341 30787 50399 30793
rect 50341 30753 50353 30787
rect 50387 30753 50399 30787
rect 50522 30784 50528 30796
rect 50483 30756 50528 30784
rect 50341 30747 50399 30753
rect 49712 30648 49740 30747
rect 50522 30744 50528 30756
rect 50580 30744 50586 30796
rect 50614 30744 50620 30796
rect 50672 30784 50678 30796
rect 51718 30784 51724 30796
rect 50672 30756 51724 30784
rect 50672 30744 50678 30756
rect 51718 30744 51724 30756
rect 51776 30744 51782 30796
rect 52362 30744 52368 30796
rect 52420 30793 52426 30796
rect 52518 30793 52546 30824
rect 52420 30787 52469 30793
rect 52420 30753 52423 30787
rect 52457 30753 52469 30787
rect 52518 30787 52588 30793
rect 52518 30756 52542 30787
rect 52420 30747 52469 30753
rect 52530 30753 52542 30756
rect 52576 30753 52588 30787
rect 52530 30747 52588 30753
rect 52420 30744 52426 30747
rect 52638 30744 52644 30796
rect 52696 30784 52702 30796
rect 52822 30784 52828 30796
rect 52696 30756 52741 30784
rect 52783 30756 52828 30784
rect 52696 30744 52702 30756
rect 52822 30744 52828 30756
rect 52880 30784 52886 30796
rect 53561 30787 53619 30793
rect 53561 30784 53573 30787
rect 52880 30756 53573 30784
rect 52880 30744 52886 30756
rect 53561 30753 53573 30756
rect 53607 30753 53619 30787
rect 53561 30747 53619 30753
rect 53650 30744 53656 30796
rect 53708 30784 53714 30796
rect 53745 30787 53803 30793
rect 53745 30784 53757 30787
rect 53708 30756 53757 30784
rect 53708 30744 53714 30756
rect 53745 30753 53757 30756
rect 53791 30753 53803 30787
rect 53745 30747 53803 30753
rect 53760 30716 53788 30747
rect 53834 30744 53840 30796
rect 53892 30784 53898 30796
rect 54478 30784 54484 30796
rect 53892 30756 53937 30784
rect 54439 30756 54484 30784
rect 53892 30744 53898 30756
rect 54478 30744 54484 30756
rect 54536 30744 54542 30796
rect 54570 30744 54576 30796
rect 54628 30784 54634 30796
rect 54628 30756 54673 30784
rect 54628 30744 54634 30756
rect 54754 30744 54760 30796
rect 54812 30784 54818 30796
rect 54849 30787 54907 30793
rect 54849 30784 54861 30787
rect 54812 30756 54861 30784
rect 54812 30744 54818 30756
rect 54849 30753 54861 30756
rect 54895 30753 54907 30787
rect 55306 30784 55312 30796
rect 55267 30756 55312 30784
rect 54849 30747 54907 30753
rect 55306 30744 55312 30756
rect 55364 30744 55370 30796
rect 55490 30784 55496 30796
rect 55451 30756 55496 30784
rect 55490 30744 55496 30756
rect 55548 30744 55554 30796
rect 57238 30784 57244 30796
rect 57199 30756 57244 30784
rect 57238 30744 57244 30756
rect 57296 30744 57302 30796
rect 57974 30784 57980 30796
rect 57935 30756 57980 30784
rect 57974 30744 57980 30756
rect 58032 30744 58038 30796
rect 55324 30716 55352 30744
rect 56042 30716 56048 30728
rect 53760 30688 54800 30716
rect 55324 30688 56048 30716
rect 51442 30648 51448 30660
rect 49712 30620 51448 30648
rect 51442 30608 51448 30620
rect 51500 30608 51506 30660
rect 51537 30651 51595 30657
rect 51537 30617 51549 30651
rect 51583 30648 51595 30651
rect 52914 30648 52920 30660
rect 51583 30620 52920 30648
rect 51583 30617 51595 30620
rect 51537 30611 51595 30617
rect 52914 30608 52920 30620
rect 52972 30608 52978 30660
rect 53377 30651 53435 30657
rect 53377 30617 53389 30651
rect 53423 30648 53435 30651
rect 54202 30648 54208 30660
rect 53423 30620 54208 30648
rect 53423 30617 53435 30620
rect 53377 30611 53435 30617
rect 54202 30608 54208 30620
rect 54260 30608 54266 30660
rect 54772 30657 54800 30688
rect 56042 30676 56048 30688
rect 56100 30676 56106 30728
rect 54757 30651 54815 30657
rect 54757 30617 54769 30651
rect 54803 30648 54815 30651
rect 56502 30648 56508 30660
rect 54803 30620 56508 30648
rect 54803 30617 54815 30620
rect 54757 30611 54815 30617
rect 56502 30608 56508 30620
rect 56560 30608 56566 30660
rect 57422 30648 57428 30660
rect 57383 30620 57428 30648
rect 57422 30608 57428 30620
rect 57480 30608 57486 30660
rect 58158 30648 58164 30660
rect 58119 30620 58164 30648
rect 58158 30608 58164 30620
rect 58216 30608 58222 30660
rect 51258 30540 51264 30592
rect 51316 30580 51322 30592
rect 57514 30580 57520 30592
rect 51316 30552 57520 30580
rect 51316 30540 51322 30552
rect 57514 30540 57520 30552
rect 57572 30540 57578 30592
rect 1104 30490 58880 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 58880 30490
rect 1104 30416 58880 30438
rect 49050 30336 49056 30388
rect 49108 30376 49114 30388
rect 49108 30348 51074 30376
rect 49108 30336 49114 30348
rect 48774 30200 48780 30252
rect 48832 30240 48838 30252
rect 49510 30240 49516 30252
rect 48832 30212 49516 30240
rect 48832 30200 48838 30212
rect 49510 30200 49516 30212
rect 49568 30200 49574 30252
rect 51046 30240 51074 30348
rect 51534 30336 51540 30388
rect 51592 30376 51598 30388
rect 52638 30376 52644 30388
rect 51592 30348 52644 30376
rect 51592 30336 51598 30348
rect 52638 30336 52644 30348
rect 52696 30336 52702 30388
rect 52917 30379 52975 30385
rect 52917 30345 52929 30379
rect 52963 30345 52975 30379
rect 52917 30339 52975 30345
rect 53101 30379 53159 30385
rect 53101 30345 53113 30379
rect 53147 30376 53159 30379
rect 53466 30376 53472 30388
rect 53147 30348 53472 30376
rect 53147 30345 53159 30348
rect 53101 30339 53159 30345
rect 51997 30311 52055 30317
rect 51997 30277 52009 30311
rect 52043 30308 52055 30311
rect 52270 30308 52276 30320
rect 52043 30280 52276 30308
rect 52043 30277 52055 30280
rect 51997 30271 52055 30277
rect 52270 30268 52276 30280
rect 52328 30268 52334 30320
rect 52362 30268 52368 30320
rect 52420 30308 52426 30320
rect 52932 30308 52960 30339
rect 53466 30336 53472 30348
rect 53524 30336 53530 30388
rect 54754 30336 54760 30388
rect 54812 30376 54818 30388
rect 55122 30376 55128 30388
rect 54812 30348 55128 30376
rect 54812 30336 54818 30348
rect 55122 30336 55128 30348
rect 55180 30336 55186 30388
rect 55674 30376 55680 30388
rect 55635 30348 55680 30376
rect 55674 30336 55680 30348
rect 55732 30336 55738 30388
rect 57974 30376 57980 30388
rect 57935 30348 57980 30376
rect 57974 30336 57980 30348
rect 58032 30336 58038 30388
rect 56781 30311 56839 30317
rect 56781 30308 56793 30311
rect 52420 30280 52960 30308
rect 53208 30280 56793 30308
rect 52420 30268 52426 30280
rect 53208 30240 53236 30280
rect 56781 30277 56793 30280
rect 56827 30277 56839 30311
rect 56781 30271 56839 30277
rect 54018 30240 54024 30252
rect 51046 30212 53236 30240
rect 53979 30212 54024 30240
rect 54018 30200 54024 30212
rect 54076 30240 54082 30252
rect 54573 30243 54631 30249
rect 54573 30240 54585 30243
rect 54076 30212 54585 30240
rect 54076 30200 54082 30212
rect 54573 30209 54585 30212
rect 54619 30209 54631 30243
rect 54573 30203 54631 30209
rect 55122 30200 55128 30252
rect 55180 30240 55186 30252
rect 57514 30240 57520 30252
rect 55180 30212 55904 30240
rect 57475 30212 57520 30240
rect 55180 30200 55186 30212
rect 47854 30132 47860 30184
rect 47912 30172 47918 30184
rect 49053 30175 49111 30181
rect 49053 30172 49065 30175
rect 47912 30144 49065 30172
rect 47912 30132 47918 30144
rect 49053 30141 49065 30144
rect 49099 30141 49111 30175
rect 49053 30135 49111 30141
rect 51905 30175 51963 30181
rect 51905 30141 51917 30175
rect 51951 30172 51963 30175
rect 52362 30172 52368 30184
rect 51951 30144 52368 30172
rect 51951 30141 51963 30144
rect 51905 30135 51963 30141
rect 52362 30132 52368 30144
rect 52420 30132 52426 30184
rect 52454 30132 52460 30184
rect 52512 30172 52518 30184
rect 52549 30175 52607 30181
rect 52549 30172 52561 30175
rect 52512 30144 52561 30172
rect 52512 30132 52518 30144
rect 52549 30141 52561 30144
rect 52595 30141 52607 30175
rect 54036 30172 54064 30200
rect 54202 30172 54208 30184
rect 52549 30135 52607 30141
rect 52932 30144 54064 30172
rect 54163 30144 54208 30172
rect 1854 30104 1860 30116
rect 1815 30076 1860 30104
rect 1854 30064 1860 30076
rect 1912 30064 1918 30116
rect 49418 30064 49424 30116
rect 49476 30104 49482 30116
rect 49758 30107 49816 30113
rect 49758 30104 49770 30107
rect 49476 30076 49770 30104
rect 49476 30064 49482 30076
rect 49758 30073 49770 30076
rect 49804 30073 49816 30107
rect 49758 30067 49816 30073
rect 49878 30064 49884 30116
rect 49936 30104 49942 30116
rect 52932 30113 52960 30144
rect 54202 30132 54208 30144
rect 54260 30172 54266 30184
rect 54435 30175 54493 30181
rect 54435 30172 54447 30175
rect 54260 30144 54447 30172
rect 54260 30132 54266 30144
rect 54435 30141 54447 30144
rect 54481 30141 54493 30175
rect 54435 30135 54493 30141
rect 54662 30132 54668 30184
rect 54720 30172 54726 30184
rect 55033 30175 55091 30181
rect 55033 30172 55045 30175
rect 54720 30144 55045 30172
rect 54720 30132 54726 30144
rect 55033 30141 55045 30144
rect 55079 30141 55091 30175
rect 55033 30135 55091 30141
rect 55306 30132 55312 30184
rect 55364 30172 55370 30184
rect 55876 30181 55904 30212
rect 57514 30200 57520 30212
rect 57572 30200 57578 30252
rect 55677 30175 55735 30181
rect 55677 30172 55689 30175
rect 55364 30144 55689 30172
rect 55364 30132 55370 30144
rect 55677 30141 55689 30144
rect 55723 30141 55735 30175
rect 55677 30135 55735 30141
rect 55861 30175 55919 30181
rect 55861 30141 55873 30175
rect 55907 30141 55919 30175
rect 55861 30135 55919 30141
rect 57701 30175 57759 30181
rect 57701 30141 57713 30175
rect 57747 30141 57759 30175
rect 57701 30135 57759 30141
rect 52917 30107 52975 30113
rect 49936 30076 51074 30104
rect 49936 30064 49942 30076
rect 1946 30036 1952 30048
rect 1907 30008 1952 30036
rect 1946 29996 1952 30008
rect 2004 29996 2010 30048
rect 48866 30036 48872 30048
rect 48827 30008 48872 30036
rect 48866 29996 48872 30008
rect 48924 29996 48930 30048
rect 48958 29996 48964 30048
rect 49016 30036 49022 30048
rect 50154 30036 50160 30048
rect 49016 30008 50160 30036
rect 49016 29996 49022 30008
rect 50154 29996 50160 30008
rect 50212 30036 50218 30048
rect 50614 30036 50620 30048
rect 50212 30008 50620 30036
rect 50212 29996 50218 30008
rect 50614 29996 50620 30008
rect 50672 29996 50678 30048
rect 50890 30036 50896 30048
rect 50851 30008 50896 30036
rect 50890 29996 50896 30008
rect 50948 29996 50954 30048
rect 51046 30036 51074 30076
rect 52917 30073 52929 30107
rect 52963 30073 52975 30107
rect 56597 30107 56655 30113
rect 52917 30067 52975 30073
rect 54036 30076 54524 30104
rect 54036 30036 54064 30076
rect 51046 30008 54064 30036
rect 54110 29996 54116 30048
rect 54168 30036 54174 30048
rect 54389 30039 54447 30045
rect 54389 30036 54401 30039
rect 54168 30008 54401 30036
rect 54168 29996 54174 30008
rect 54389 30005 54401 30008
rect 54435 30005 54447 30039
rect 54496 30036 54524 30076
rect 56597 30073 56609 30107
rect 56643 30104 56655 30107
rect 56778 30104 56784 30116
rect 56643 30076 56784 30104
rect 56643 30073 56655 30076
rect 56597 30067 56655 30073
rect 56778 30064 56784 30076
rect 56836 30064 56842 30116
rect 56870 30064 56876 30116
rect 56928 30104 56934 30116
rect 57716 30104 57744 30135
rect 56928 30076 57744 30104
rect 56928 30064 56934 30076
rect 57514 30036 57520 30048
rect 54496 30008 57520 30036
rect 54389 29999 54447 30005
rect 57514 29996 57520 30008
rect 57572 29996 57578 30048
rect 1104 29946 58880 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 58880 29946
rect 1104 29872 58880 29894
rect 48685 29835 48743 29841
rect 48685 29801 48697 29835
rect 48731 29801 48743 29835
rect 49418 29832 49424 29844
rect 49379 29804 49424 29832
rect 48685 29795 48743 29801
rect 48700 29764 48728 29795
rect 49418 29792 49424 29804
rect 49476 29792 49482 29844
rect 57977 29835 58035 29841
rect 49896 29804 57100 29832
rect 49896 29764 49924 29804
rect 50433 29767 50491 29773
rect 50433 29764 50445 29767
rect 48700 29736 49924 29764
rect 50172 29736 50445 29764
rect 1857 29699 1915 29705
rect 1857 29665 1869 29699
rect 1903 29696 1915 29699
rect 2130 29696 2136 29708
rect 1903 29668 2136 29696
rect 1903 29665 1915 29668
rect 1857 29659 1915 29665
rect 2130 29656 2136 29668
rect 2188 29656 2194 29708
rect 48869 29699 48927 29705
rect 48869 29665 48881 29699
rect 48915 29696 48927 29699
rect 48958 29696 48964 29708
rect 48915 29668 48964 29696
rect 48915 29665 48927 29668
rect 48869 29659 48927 29665
rect 48958 29656 48964 29668
rect 49016 29656 49022 29708
rect 50172 29705 50200 29736
rect 50433 29733 50445 29736
rect 50479 29764 50491 29767
rect 51258 29764 51264 29776
rect 50479 29736 51264 29764
rect 50479 29733 50491 29736
rect 50433 29727 50491 29733
rect 51258 29724 51264 29736
rect 51316 29724 51322 29776
rect 51994 29724 52000 29776
rect 52052 29764 52058 29776
rect 52641 29767 52699 29773
rect 52641 29764 52653 29767
rect 52052 29736 52653 29764
rect 52052 29724 52058 29736
rect 52641 29733 52653 29736
rect 52687 29733 52699 29767
rect 52641 29727 52699 29733
rect 52822 29724 52828 29776
rect 52880 29764 52886 29776
rect 53282 29764 53288 29776
rect 52880 29736 53288 29764
rect 52880 29724 52886 29736
rect 53282 29724 53288 29736
rect 53340 29724 53346 29776
rect 54205 29767 54263 29773
rect 54205 29733 54217 29767
rect 54251 29764 54263 29767
rect 54938 29764 54944 29776
rect 54251 29736 54944 29764
rect 54251 29733 54263 29736
rect 54205 29727 54263 29733
rect 54938 29724 54944 29736
rect 54996 29724 55002 29776
rect 49329 29699 49387 29705
rect 49329 29665 49341 29699
rect 49375 29665 49387 29699
rect 49329 29659 49387 29665
rect 49513 29699 49571 29705
rect 49513 29665 49525 29699
rect 49559 29696 49571 29699
rect 50157 29699 50215 29705
rect 49559 29668 50108 29696
rect 49559 29665 49571 29668
rect 49513 29659 49571 29665
rect 49344 29560 49372 29659
rect 49970 29628 49976 29640
rect 49931 29600 49976 29628
rect 49970 29588 49976 29600
rect 50028 29588 50034 29640
rect 50080 29628 50108 29668
rect 50157 29665 50169 29699
rect 50203 29665 50215 29699
rect 50157 29659 50215 29665
rect 50890 29656 50896 29708
rect 50948 29696 50954 29708
rect 51445 29699 51503 29705
rect 51445 29696 51457 29699
rect 50948 29668 51457 29696
rect 50948 29656 50954 29668
rect 51445 29665 51457 29668
rect 51491 29665 51503 29699
rect 52362 29696 52368 29708
rect 52323 29668 52368 29696
rect 51445 29659 51503 29665
rect 52362 29656 52368 29668
rect 52420 29656 52426 29708
rect 52454 29656 52460 29708
rect 52512 29696 52518 29708
rect 52733 29699 52791 29705
rect 52733 29696 52745 29699
rect 52512 29668 52745 29696
rect 52512 29656 52518 29668
rect 52733 29665 52745 29668
rect 52779 29665 52791 29699
rect 52733 29659 52791 29665
rect 53193 29699 53251 29705
rect 53193 29665 53205 29699
rect 53239 29665 53251 29699
rect 53193 29659 53251 29665
rect 50080 29600 50384 29628
rect 50249 29563 50307 29569
rect 50249 29560 50261 29563
rect 49344 29532 50261 29560
rect 50249 29529 50261 29532
rect 50295 29529 50307 29563
rect 50356 29560 50384 29600
rect 50430 29588 50436 29640
rect 50488 29628 50494 29640
rect 50525 29631 50583 29637
rect 50525 29628 50537 29631
rect 50488 29600 50537 29628
rect 50488 29588 50494 29600
rect 50525 29597 50537 29600
rect 50571 29597 50583 29631
rect 52270 29628 52276 29640
rect 52231 29600 52276 29628
rect 50525 29591 50583 29597
rect 52270 29588 52276 29600
rect 52328 29628 52334 29640
rect 53208 29628 53236 29659
rect 54018 29656 54024 29708
rect 54076 29696 54082 29708
rect 54553 29699 54611 29705
rect 54553 29696 54565 29699
rect 54076 29668 54565 29696
rect 54076 29656 54082 29668
rect 54553 29665 54565 29668
rect 54599 29665 54611 29699
rect 54553 29659 54611 29665
rect 54846 29656 54852 29708
rect 54904 29696 54910 29708
rect 57072 29705 57100 29804
rect 57977 29801 57989 29835
rect 58023 29832 58035 29835
rect 58250 29832 58256 29844
rect 58023 29804 58256 29832
rect 58023 29801 58035 29804
rect 57977 29795 58035 29801
rect 58250 29792 58256 29804
rect 58308 29792 58314 29844
rect 57057 29699 57115 29705
rect 54904 29668 55720 29696
rect 54904 29656 54910 29668
rect 54202 29628 54208 29640
rect 52328 29600 53236 29628
rect 54115 29600 54208 29628
rect 52328 29588 52334 29600
rect 54202 29588 54208 29600
rect 54260 29628 54266 29640
rect 54297 29631 54355 29637
rect 54297 29628 54309 29631
rect 54260 29600 54309 29628
rect 54260 29588 54266 29600
rect 54297 29597 54309 29600
rect 54343 29597 54355 29631
rect 54297 29591 54355 29597
rect 53742 29560 53748 29572
rect 50356 29532 53748 29560
rect 50249 29523 50307 29529
rect 53742 29520 53748 29532
rect 53800 29520 53806 29572
rect 55692 29569 55720 29668
rect 57057 29665 57069 29699
rect 57103 29665 57115 29699
rect 57057 29659 57115 29665
rect 57882 29656 57888 29708
rect 57940 29696 57946 29708
rect 58161 29699 58219 29705
rect 58161 29696 58173 29699
rect 57940 29668 58173 29696
rect 57940 29656 57946 29668
rect 58161 29665 58173 29668
rect 58207 29665 58219 29699
rect 58161 29659 58219 29665
rect 55950 29588 55956 29640
rect 56008 29628 56014 29640
rect 56873 29631 56931 29637
rect 56873 29628 56885 29631
rect 56008 29600 56885 29628
rect 56008 29588 56014 29600
rect 56873 29597 56885 29600
rect 56919 29597 56931 29631
rect 56873 29591 56931 29597
rect 55677 29563 55735 29569
rect 55677 29529 55689 29563
rect 55723 29529 55735 29563
rect 57238 29560 57244 29572
rect 57199 29532 57244 29560
rect 55677 29523 55735 29529
rect 57238 29520 57244 29532
rect 57296 29520 57302 29572
rect 1394 29452 1400 29504
rect 1452 29492 1458 29504
rect 1949 29495 2007 29501
rect 1949 29492 1961 29495
rect 1452 29464 1961 29492
rect 1452 29452 1458 29464
rect 1949 29461 1961 29464
rect 1995 29461 2007 29495
rect 2682 29492 2688 29504
rect 2643 29464 2688 29492
rect 1949 29455 2007 29461
rect 2682 29452 2688 29464
rect 2740 29452 2746 29504
rect 51534 29492 51540 29504
rect 51495 29464 51540 29492
rect 51534 29452 51540 29464
rect 51592 29452 51598 29504
rect 1104 29402 58880 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 58880 29402
rect 1104 29328 58880 29350
rect 1854 29248 1860 29300
rect 1912 29288 1918 29300
rect 1949 29291 2007 29297
rect 1949 29288 1961 29291
rect 1912 29260 1961 29288
rect 1912 29248 1918 29260
rect 1949 29257 1961 29260
rect 1995 29257 2007 29291
rect 1949 29251 2007 29257
rect 47673 29291 47731 29297
rect 47673 29257 47685 29291
rect 47719 29288 47731 29291
rect 48314 29288 48320 29300
rect 47719 29260 48320 29288
rect 47719 29257 47731 29260
rect 47673 29251 47731 29257
rect 48314 29248 48320 29260
rect 48372 29248 48378 29300
rect 48961 29291 49019 29297
rect 48961 29257 48973 29291
rect 49007 29288 49019 29291
rect 49878 29288 49884 29300
rect 49007 29260 49884 29288
rect 49007 29257 49019 29260
rect 48961 29251 49019 29257
rect 49878 29248 49884 29260
rect 49936 29248 49942 29300
rect 49970 29248 49976 29300
rect 50028 29288 50034 29300
rect 50065 29291 50123 29297
rect 50065 29288 50077 29291
rect 50028 29260 50077 29288
rect 50028 29248 50034 29260
rect 50065 29257 50077 29260
rect 50111 29288 50123 29291
rect 50430 29288 50436 29300
rect 50111 29260 50436 29288
rect 50111 29257 50123 29260
rect 50065 29251 50123 29257
rect 50430 29248 50436 29260
rect 50488 29248 50494 29300
rect 51534 29288 51540 29300
rect 51368 29260 51540 29288
rect 50525 29223 50583 29229
rect 50525 29189 50537 29223
rect 50571 29220 50583 29223
rect 50614 29220 50620 29232
rect 50571 29192 50620 29220
rect 50571 29189 50583 29192
rect 50525 29183 50583 29189
rect 50614 29180 50620 29192
rect 50672 29180 50678 29232
rect 1581 29155 1639 29161
rect 1581 29121 1593 29155
rect 1627 29152 1639 29155
rect 2682 29152 2688 29164
rect 1627 29124 2688 29152
rect 1627 29121 1639 29124
rect 1581 29115 1639 29121
rect 2682 29112 2688 29124
rect 2740 29112 2746 29164
rect 49510 29152 49516 29164
rect 49471 29124 49516 29152
rect 49510 29112 49516 29124
rect 49568 29112 49574 29164
rect 50706 29152 50712 29164
rect 50264 29124 50712 29152
rect 1762 29084 1768 29096
rect 1723 29056 1768 29084
rect 1762 29044 1768 29056
rect 1820 29044 1826 29096
rect 47854 29084 47860 29096
rect 47815 29056 47860 29084
rect 47854 29044 47860 29056
rect 47912 29044 47918 29096
rect 49050 29044 49056 29096
rect 49108 29084 49114 29096
rect 50264 29093 50292 29124
rect 50706 29112 50712 29124
rect 50764 29152 50770 29164
rect 51368 29152 51396 29260
rect 51534 29248 51540 29260
rect 51592 29248 51598 29300
rect 54018 29288 54024 29300
rect 53979 29260 54024 29288
rect 54018 29248 54024 29260
rect 54076 29248 54082 29300
rect 55769 29291 55827 29297
rect 55769 29257 55781 29291
rect 55815 29288 55827 29291
rect 56870 29288 56876 29300
rect 55815 29260 56876 29288
rect 55815 29257 55827 29260
rect 55769 29251 55827 29257
rect 56870 29248 56876 29260
rect 56928 29248 56934 29300
rect 57241 29291 57299 29297
rect 57241 29257 57253 29291
rect 57287 29288 57299 29291
rect 57606 29288 57612 29300
rect 57287 29260 57612 29288
rect 57287 29257 57299 29260
rect 57241 29251 57299 29257
rect 57606 29248 57612 29260
rect 57664 29248 57670 29300
rect 51442 29180 51448 29232
rect 51500 29220 51506 29232
rect 55490 29220 55496 29232
rect 51500 29192 55496 29220
rect 51500 29180 51506 29192
rect 55490 29180 55496 29192
rect 55548 29180 55554 29232
rect 56502 29220 56508 29232
rect 56463 29192 56508 29220
rect 56502 29180 56508 29192
rect 56560 29180 56566 29232
rect 50764 29124 51580 29152
rect 50764 29112 50770 29124
rect 49421 29087 49479 29093
rect 49421 29084 49433 29087
rect 49108 29056 49433 29084
rect 49108 29044 49114 29056
rect 49421 29053 49433 29056
rect 49467 29053 49479 29087
rect 49421 29047 49479 29053
rect 49605 29087 49663 29093
rect 49605 29053 49617 29087
rect 49651 29053 49663 29087
rect 49605 29047 49663 29053
rect 50249 29087 50307 29093
rect 50249 29053 50261 29087
rect 50295 29053 50307 29087
rect 50249 29047 50307 29053
rect 50341 29087 50399 29093
rect 50341 29053 50353 29087
rect 50387 29053 50399 29087
rect 50341 29047 50399 29053
rect 50617 29087 50675 29093
rect 50617 29053 50629 29087
rect 50663 29084 50675 29087
rect 50890 29084 50896 29096
rect 50663 29056 50896 29084
rect 50663 29053 50675 29056
rect 50617 29047 50675 29053
rect 49620 29016 49648 29047
rect 50356 29016 50384 29047
rect 50890 29044 50896 29056
rect 50948 29044 50954 29096
rect 51442 29084 51448 29096
rect 51046 29056 51448 29084
rect 51046 29016 51074 29056
rect 51442 29044 51448 29056
rect 51500 29044 51506 29096
rect 51552 29093 51580 29124
rect 52362 29112 52368 29164
rect 52420 29152 52426 29164
rect 52457 29155 52515 29161
rect 52457 29152 52469 29155
rect 52420 29124 52469 29152
rect 52420 29112 52426 29124
rect 52457 29121 52469 29124
rect 52503 29121 52515 29155
rect 52457 29115 52515 29121
rect 52733 29155 52791 29161
rect 52733 29121 52745 29155
rect 52779 29121 52791 29155
rect 52733 29115 52791 29121
rect 51537 29087 51595 29093
rect 51537 29053 51549 29087
rect 51583 29053 51595 29087
rect 51718 29084 51724 29096
rect 51679 29056 51724 29084
rect 51537 29047 51595 29053
rect 51718 29044 51724 29056
rect 51776 29044 51782 29096
rect 51813 29087 51871 29093
rect 51813 29053 51825 29087
rect 51859 29084 51871 29087
rect 51994 29084 52000 29096
rect 51859 29056 52000 29084
rect 51859 29053 51871 29056
rect 51813 29047 51871 29053
rect 49620 28988 51074 29016
rect 51166 28976 51172 29028
rect 51224 29016 51230 29028
rect 51828 29016 51856 29047
rect 51994 29044 52000 29056
rect 52052 29044 52058 29096
rect 52273 29087 52331 29093
rect 52273 29053 52285 29087
rect 52319 29084 52331 29087
rect 52638 29084 52644 29096
rect 52319 29056 52644 29084
rect 52319 29053 52331 29056
rect 52273 29047 52331 29053
rect 52638 29044 52644 29056
rect 52696 29044 52702 29096
rect 51224 28988 51856 29016
rect 51224 28976 51230 28988
rect 51902 28976 51908 29028
rect 51960 29016 51966 29028
rect 52748 29016 52776 29115
rect 53742 29112 53748 29164
rect 53800 29152 53806 29164
rect 53800 29124 54248 29152
rect 53800 29112 53806 29124
rect 52825 29087 52883 29093
rect 52825 29053 52837 29087
rect 52871 29084 52883 29087
rect 53466 29084 53472 29096
rect 52871 29056 53472 29084
rect 52871 29053 52883 29056
rect 52825 29047 52883 29053
rect 53466 29044 53472 29056
rect 53524 29044 53530 29096
rect 54021 29087 54079 29093
rect 54021 29053 54033 29087
rect 54067 29084 54079 29087
rect 54110 29084 54116 29096
rect 54067 29056 54116 29084
rect 54067 29053 54079 29056
rect 54021 29047 54079 29053
rect 54110 29044 54116 29056
rect 54168 29044 54174 29096
rect 54220 29093 54248 29124
rect 54205 29087 54263 29093
rect 54205 29053 54217 29087
rect 54251 29053 54263 29087
rect 54938 29084 54944 29096
rect 54899 29056 54944 29084
rect 54205 29047 54263 29053
rect 54938 29044 54944 29056
rect 54996 29044 55002 29096
rect 55122 29084 55128 29096
rect 55083 29056 55128 29084
rect 55122 29044 55128 29056
rect 55180 29044 55186 29096
rect 55953 29087 56011 29093
rect 55953 29053 55965 29087
rect 55999 29084 56011 29087
rect 56226 29084 56232 29096
rect 55999 29056 56232 29084
rect 55999 29053 56011 29056
rect 55953 29047 56011 29053
rect 56226 29044 56232 29056
rect 56284 29044 56290 29096
rect 56410 29084 56416 29096
rect 56371 29056 56416 29084
rect 56410 29044 56416 29056
rect 56468 29044 56474 29096
rect 57425 29087 57483 29093
rect 57425 29053 57437 29087
rect 57471 29084 57483 29087
rect 57882 29084 57888 29096
rect 57471 29056 57888 29084
rect 57471 29053 57483 29056
rect 57425 29047 57483 29053
rect 57882 29044 57888 29056
rect 57940 29044 57946 29096
rect 51960 28988 52776 29016
rect 55033 29019 55091 29025
rect 51960 28976 51966 28988
rect 55033 28985 55045 29019
rect 55079 29016 55091 29019
rect 55214 29016 55220 29028
rect 55079 28988 55220 29016
rect 55079 28985 55091 28988
rect 55033 28979 55091 28985
rect 55214 28976 55220 28988
rect 55272 28976 55278 29028
rect 57974 29016 57980 29028
rect 57935 28988 57980 29016
rect 57974 28976 57980 28988
rect 58032 28976 58038 29028
rect 58158 29016 58164 29028
rect 58119 28988 58164 29016
rect 58158 28976 58164 28988
rect 58216 28976 58222 29028
rect 49234 28908 49240 28960
rect 49292 28948 49298 28960
rect 50982 28948 50988 28960
rect 49292 28920 50988 28948
rect 49292 28908 49298 28920
rect 50982 28908 50988 28920
rect 51040 28908 51046 28960
rect 51261 28951 51319 28957
rect 51261 28917 51273 28951
rect 51307 28948 51319 28951
rect 51718 28948 51724 28960
rect 51307 28920 51724 28948
rect 51307 28917 51319 28920
rect 51261 28911 51319 28917
rect 51718 28908 51724 28920
rect 51776 28908 51782 28960
rect 1104 28858 58880 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 50326 28858
rect 50378 28806 50390 28858
rect 50442 28806 50454 28858
rect 50506 28806 50518 28858
rect 50570 28806 58880 28858
rect 1104 28784 58880 28806
rect 47765 28747 47823 28753
rect 47765 28713 47777 28747
rect 47811 28744 47823 28747
rect 47854 28744 47860 28756
rect 47811 28716 47860 28744
rect 47811 28713 47823 28716
rect 47765 28707 47823 28713
rect 47854 28704 47860 28716
rect 47912 28704 47918 28756
rect 49418 28744 49424 28756
rect 47964 28716 49424 28744
rect 1765 28611 1823 28617
rect 1765 28577 1777 28611
rect 1811 28608 1823 28611
rect 3970 28608 3976 28620
rect 1811 28580 3976 28608
rect 1811 28577 1823 28580
rect 1765 28571 1823 28577
rect 3970 28568 3976 28580
rect 4028 28568 4034 28620
rect 47964 28617 47992 28716
rect 49418 28704 49424 28716
rect 49476 28704 49482 28756
rect 50433 28747 50491 28753
rect 50433 28713 50445 28747
rect 50479 28744 50491 28747
rect 51442 28744 51448 28756
rect 50479 28716 51448 28744
rect 50479 28713 50491 28716
rect 50433 28707 50491 28713
rect 51442 28704 51448 28716
rect 51500 28704 51506 28756
rect 52454 28744 52460 28756
rect 51552 28716 52224 28744
rect 52415 28716 52460 28744
rect 51552 28676 51580 28716
rect 48424 28648 51580 28676
rect 48424 28617 48452 28648
rect 51626 28636 51632 28688
rect 51684 28676 51690 28688
rect 52196 28676 52224 28716
rect 52454 28704 52460 28716
rect 52512 28704 52518 28756
rect 55122 28704 55128 28756
rect 55180 28744 55186 28756
rect 55217 28747 55275 28753
rect 55217 28744 55229 28747
rect 55180 28716 55229 28744
rect 55180 28704 55186 28716
rect 55217 28713 55229 28716
rect 55263 28713 55275 28747
rect 55217 28707 55275 28713
rect 57974 28704 57980 28756
rect 58032 28744 58038 28756
rect 58161 28747 58219 28753
rect 58161 28744 58173 28747
rect 58032 28716 58173 28744
rect 58032 28704 58038 28716
rect 58161 28713 58173 28716
rect 58207 28713 58219 28747
rect 58161 28707 58219 28713
rect 55306 28676 55312 28688
rect 51684 28648 52132 28676
rect 52196 28648 55312 28676
rect 51684 28636 51690 28648
rect 47305 28611 47363 28617
rect 47305 28577 47317 28611
rect 47351 28577 47363 28611
rect 47305 28571 47363 28577
rect 47949 28611 48007 28617
rect 47949 28577 47961 28611
rect 47995 28577 48007 28611
rect 47949 28571 48007 28577
rect 48409 28611 48467 28617
rect 48409 28577 48421 28611
rect 48455 28577 48467 28611
rect 49050 28608 49056 28620
rect 49011 28580 49056 28608
rect 48409 28571 48467 28577
rect 1949 28543 2007 28549
rect 1949 28509 1961 28543
rect 1995 28540 2007 28543
rect 3142 28540 3148 28552
rect 1995 28512 3148 28540
rect 1995 28509 2007 28512
rect 1949 28503 2007 28509
rect 3142 28500 3148 28512
rect 3200 28500 3206 28552
rect 47320 28540 47348 28571
rect 49050 28568 49056 28580
rect 49108 28568 49114 28620
rect 49234 28608 49240 28620
rect 49195 28580 49240 28608
rect 49234 28568 49240 28580
rect 49292 28568 49298 28620
rect 49694 28608 49700 28620
rect 49655 28580 49700 28608
rect 49694 28568 49700 28580
rect 49752 28568 49758 28620
rect 49881 28611 49939 28617
rect 49881 28577 49893 28611
rect 49927 28608 49939 28611
rect 49970 28608 49976 28620
rect 49927 28580 49976 28608
rect 49927 28577 49939 28580
rect 49881 28571 49939 28577
rect 49970 28568 49976 28580
rect 50028 28568 50034 28620
rect 50341 28611 50399 28617
rect 50341 28577 50353 28611
rect 50387 28608 50399 28611
rect 50614 28608 50620 28620
rect 50387 28580 50620 28608
rect 50387 28577 50399 28580
rect 50341 28571 50399 28577
rect 50614 28568 50620 28580
rect 50672 28568 50678 28620
rect 51718 28608 51724 28620
rect 51679 28580 51724 28608
rect 51718 28568 51724 28580
rect 51776 28568 51782 28620
rect 51902 28608 51908 28620
rect 51863 28580 51908 28608
rect 51902 28568 51908 28580
rect 51960 28568 51966 28620
rect 52104 28617 52132 28648
rect 55306 28636 55312 28648
rect 55364 28636 55370 28688
rect 52089 28611 52147 28617
rect 52089 28577 52101 28611
rect 52135 28577 52147 28611
rect 52089 28571 52147 28577
rect 52178 28568 52184 28620
rect 52236 28608 52242 28620
rect 52273 28611 52331 28617
rect 52273 28608 52285 28611
rect 52236 28580 52285 28608
rect 52236 28568 52242 28580
rect 52273 28577 52285 28580
rect 52319 28577 52331 28611
rect 52273 28571 52331 28577
rect 52454 28568 52460 28620
rect 52512 28608 52518 28620
rect 53541 28611 53599 28617
rect 53541 28608 53553 28611
rect 52512 28580 53553 28608
rect 52512 28568 52518 28580
rect 53541 28577 53553 28580
rect 53587 28577 53599 28611
rect 55125 28611 55183 28617
rect 55125 28608 55137 28611
rect 53541 28571 53599 28577
rect 54680 28580 55137 28608
rect 48866 28540 48872 28552
rect 47320 28512 48872 28540
rect 48866 28500 48872 28512
rect 48924 28500 48930 28552
rect 49789 28543 49847 28549
rect 49789 28509 49801 28543
rect 49835 28540 49847 28543
rect 51920 28540 51948 28568
rect 49835 28512 51948 28540
rect 51997 28543 52055 28549
rect 49835 28509 49847 28512
rect 49789 28503 49847 28509
rect 51997 28509 52009 28543
rect 52043 28540 52055 28543
rect 53190 28540 53196 28552
rect 52043 28512 53196 28540
rect 52043 28509 52055 28512
rect 51997 28503 52055 28509
rect 53190 28500 53196 28512
rect 53248 28500 53254 28552
rect 53285 28543 53343 28549
rect 53285 28509 53297 28543
rect 53331 28509 53343 28543
rect 53285 28503 53343 28509
rect 2130 28472 2136 28484
rect 2091 28444 2136 28472
rect 2130 28432 2136 28444
rect 2188 28432 2194 28484
rect 49053 28475 49111 28481
rect 49053 28441 49065 28475
rect 49099 28472 49111 28475
rect 52178 28472 52184 28484
rect 49099 28444 52184 28472
rect 49099 28441 49111 28444
rect 49053 28435 49111 28441
rect 52178 28432 52184 28444
rect 52236 28432 52242 28484
rect 52914 28432 52920 28484
rect 52972 28472 52978 28484
rect 53300 28472 53328 28503
rect 52972 28444 53328 28472
rect 52972 28432 52978 28444
rect 47121 28407 47179 28413
rect 47121 28373 47133 28407
rect 47167 28404 47179 28407
rect 48774 28404 48780 28416
rect 47167 28376 48780 28404
rect 47167 28373 47179 28376
rect 47121 28367 47179 28373
rect 48774 28364 48780 28376
rect 48832 28364 48838 28416
rect 53300 28404 53328 28444
rect 54202 28404 54208 28416
rect 53300 28376 54208 28404
rect 54202 28364 54208 28376
rect 54260 28364 54266 28416
rect 54294 28364 54300 28416
rect 54352 28404 54358 28416
rect 54680 28413 54708 28580
rect 55125 28577 55137 28580
rect 55171 28577 55183 28611
rect 56870 28608 56876 28620
rect 56831 28580 56876 28608
rect 55125 28571 55183 28577
rect 56870 28568 56876 28580
rect 56928 28568 56934 28620
rect 57054 28608 57060 28620
rect 57015 28580 57060 28608
rect 57054 28568 57060 28580
rect 57112 28568 57118 28620
rect 57514 28608 57520 28620
rect 57475 28580 57520 28608
rect 57514 28568 57520 28580
rect 57572 28568 57578 28620
rect 56594 28500 56600 28552
rect 56652 28540 56658 28552
rect 57701 28543 57759 28549
rect 57701 28540 57713 28543
rect 56652 28512 57713 28540
rect 56652 28500 56658 28512
rect 57701 28509 57713 28512
rect 57747 28509 57759 28543
rect 57701 28503 57759 28509
rect 54665 28407 54723 28413
rect 54665 28404 54677 28407
rect 54352 28376 54677 28404
rect 54352 28364 54358 28376
rect 54665 28373 54677 28376
rect 54711 28373 54723 28407
rect 54665 28367 54723 28373
rect 1104 28314 58880 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 58880 28314
rect 1104 28240 58880 28262
rect 1762 28160 1768 28212
rect 1820 28200 1826 28212
rect 2501 28203 2559 28209
rect 2501 28200 2513 28203
rect 1820 28172 2513 28200
rect 1820 28160 1826 28172
rect 2501 28169 2513 28172
rect 2547 28169 2559 28203
rect 3142 28200 3148 28212
rect 3103 28172 3148 28200
rect 2501 28163 2559 28169
rect 3142 28160 3148 28172
rect 3200 28160 3206 28212
rect 3970 28200 3976 28212
rect 3931 28172 3976 28200
rect 3970 28160 3976 28172
rect 4028 28160 4034 28212
rect 50157 28203 50215 28209
rect 50157 28169 50169 28203
rect 50203 28200 50215 28203
rect 50614 28200 50620 28212
rect 50203 28172 50620 28200
rect 50203 28169 50215 28172
rect 50157 28163 50215 28169
rect 50614 28160 50620 28172
rect 50672 28160 50678 28212
rect 52454 28200 52460 28212
rect 52415 28172 52460 28200
rect 52454 28160 52460 28172
rect 52512 28160 52518 28212
rect 52748 28172 53144 28200
rect 51997 28135 52055 28141
rect 51997 28101 52009 28135
rect 52043 28132 52055 28135
rect 52748 28132 52776 28172
rect 52043 28104 52776 28132
rect 52043 28101 52055 28104
rect 51997 28095 52055 28101
rect 52822 28092 52828 28144
rect 52880 28092 52886 28144
rect 2682 27996 2688 28008
rect 2643 27968 2688 27996
rect 2682 27956 2688 27968
rect 2740 27996 2746 28008
rect 3329 27999 3387 28005
rect 3329 27996 3341 27999
rect 2740 27968 3341 27996
rect 2740 27956 2746 27968
rect 3329 27965 3341 27968
rect 3375 27965 3387 27999
rect 48774 27996 48780 28008
rect 48687 27968 48780 27996
rect 3329 27959 3387 27965
rect 48774 27956 48780 27968
rect 48832 27956 48838 28008
rect 50617 27999 50675 28005
rect 50617 27965 50629 27999
rect 50663 27965 50675 27999
rect 50617 27959 50675 27965
rect 1857 27931 1915 27937
rect 1857 27897 1869 27931
rect 1903 27928 1915 27931
rect 2038 27928 2044 27940
rect 1903 27900 2044 27928
rect 1903 27897 1915 27900
rect 1857 27891 1915 27897
rect 2038 27888 2044 27900
rect 2096 27888 2102 27940
rect 1946 27860 1952 27872
rect 1907 27832 1952 27860
rect 1946 27820 1952 27832
rect 2004 27820 2010 27872
rect 48792 27860 48820 27956
rect 49044 27931 49102 27937
rect 49044 27897 49056 27931
rect 49090 27928 49102 27931
rect 50632 27928 50660 27959
rect 50706 27956 50712 28008
rect 50764 27996 50770 28008
rect 50801 27999 50859 28005
rect 50801 27996 50813 27999
rect 50764 27968 50813 27996
rect 50764 27956 50770 27968
rect 50801 27965 50813 27968
rect 50847 27965 50859 27999
rect 51074 27996 51080 28008
rect 50801 27959 50859 27965
rect 50908 27968 51080 27996
rect 50908 27928 50936 27968
rect 51074 27956 51080 27968
rect 51132 27956 51138 28008
rect 51534 27956 51540 28008
rect 51592 27996 51598 28008
rect 51813 27999 51871 28005
rect 51813 27996 51825 27999
rect 51592 27968 51825 27996
rect 51592 27956 51598 27968
rect 51813 27965 51825 27968
rect 51859 27996 51871 27999
rect 52270 27996 52276 28008
rect 51859 27968 52276 27996
rect 51859 27965 51871 27968
rect 51813 27959 51871 27965
rect 52270 27956 52276 27968
rect 52328 27956 52334 28008
rect 52730 27996 52736 28008
rect 52691 27968 52736 27996
rect 52730 27956 52736 27968
rect 52788 27956 52794 28008
rect 52840 28005 52868 28092
rect 52822 27999 52880 28005
rect 52822 27965 52834 27999
rect 52868 27965 52880 27999
rect 52822 27959 52880 27965
rect 52917 27999 52975 28005
rect 52917 27965 52929 27999
rect 52963 27996 52975 27999
rect 53006 27996 53012 28008
rect 52963 27968 53012 27996
rect 52963 27965 52975 27968
rect 52917 27959 52975 27965
rect 53006 27956 53012 27968
rect 53064 27956 53070 28008
rect 53116 28005 53144 28172
rect 56870 28160 56876 28212
rect 56928 28200 56934 28212
rect 57425 28203 57483 28209
rect 57425 28200 57437 28203
rect 56928 28172 57437 28200
rect 56928 28160 56934 28172
rect 57425 28169 57437 28172
rect 57471 28169 57483 28203
rect 57425 28163 57483 28169
rect 54202 28092 54208 28144
rect 54260 28132 54266 28144
rect 54389 28135 54447 28141
rect 54389 28132 54401 28135
rect 54260 28104 54401 28132
rect 54260 28092 54266 28104
rect 54389 28101 54401 28104
rect 54435 28101 54447 28135
rect 54389 28095 54447 28101
rect 55122 28092 55128 28144
rect 55180 28092 55186 28144
rect 54481 28067 54539 28073
rect 54481 28033 54493 28067
rect 54527 28064 54539 28067
rect 54662 28064 54668 28076
rect 54527 28036 54668 28064
rect 54527 28033 54539 28036
rect 54481 28027 54539 28033
rect 54662 28024 54668 28036
rect 54720 28064 54726 28076
rect 55140 28064 55168 28092
rect 54720 28036 55168 28064
rect 54720 28024 54726 28036
rect 53101 27999 53159 28005
rect 53101 27965 53113 27999
rect 53147 27996 53159 27999
rect 54205 27999 54263 28005
rect 54205 27996 54217 27999
rect 53147 27968 54217 27996
rect 53147 27965 53159 27968
rect 53101 27959 53159 27965
rect 54205 27965 54217 27968
rect 54251 27965 54263 27999
rect 54205 27959 54263 27965
rect 55030 27956 55036 28008
rect 55088 27996 55094 28008
rect 55125 27999 55183 28005
rect 55125 27996 55137 27999
rect 55088 27968 55137 27996
rect 55088 27956 55094 27968
rect 55125 27965 55137 27968
rect 55171 27965 55183 27999
rect 55125 27959 55183 27965
rect 55214 27956 55220 28008
rect 55272 27996 55278 28008
rect 55381 27999 55439 28005
rect 55381 27996 55393 27999
rect 55272 27968 55393 27996
rect 55272 27956 55278 27968
rect 55381 27965 55393 27968
rect 55427 27965 55439 27999
rect 55381 27959 55439 27965
rect 57057 27999 57115 28005
rect 57057 27965 57069 27999
rect 57103 27965 57115 27999
rect 57238 27996 57244 28008
rect 57199 27968 57244 27996
rect 57057 27959 57115 27965
rect 49090 27900 50292 27928
rect 50632 27900 50936 27928
rect 51629 27931 51687 27937
rect 49090 27897 49102 27900
rect 49044 27891 49102 27897
rect 49234 27860 49240 27872
rect 48792 27832 49240 27860
rect 49234 27820 49240 27832
rect 49292 27820 49298 27872
rect 50264 27860 50292 27900
rect 51629 27897 51641 27931
rect 51675 27897 51687 27931
rect 51629 27891 51687 27897
rect 50709 27863 50767 27869
rect 50709 27860 50721 27863
rect 50264 27832 50721 27860
rect 50709 27829 50721 27832
rect 50755 27829 50767 27863
rect 51644 27860 51672 27891
rect 52178 27888 52184 27940
rect 52236 27928 52242 27940
rect 57072 27928 57100 27959
rect 57238 27956 57244 27968
rect 57296 27956 57302 28008
rect 52236 27900 57100 27928
rect 52236 27888 52242 27900
rect 53466 27860 53472 27872
rect 51644 27832 53472 27860
rect 50709 27823 50767 27829
rect 53466 27820 53472 27832
rect 53524 27820 53530 27872
rect 54018 27860 54024 27872
rect 53979 27832 54024 27860
rect 54018 27820 54024 27832
rect 54076 27820 54082 27872
rect 56502 27860 56508 27872
rect 56463 27832 56508 27860
rect 56502 27820 56508 27832
rect 56560 27820 56566 27872
rect 1104 27770 58880 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 50326 27770
rect 50378 27718 50390 27770
rect 50442 27718 50454 27770
rect 50506 27718 50518 27770
rect 50570 27718 58880 27770
rect 1104 27696 58880 27718
rect 49694 27616 49700 27668
rect 49752 27656 49758 27668
rect 49878 27656 49884 27668
rect 49752 27628 49884 27656
rect 49752 27616 49758 27628
rect 49878 27616 49884 27628
rect 49936 27656 49942 27668
rect 50525 27659 50583 27665
rect 49936 27628 50476 27656
rect 49936 27616 49942 27628
rect 50246 27588 50252 27600
rect 49252 27560 50252 27588
rect 1673 27523 1731 27529
rect 1673 27489 1685 27523
rect 1719 27520 1731 27523
rect 3326 27520 3332 27532
rect 1719 27492 3332 27520
rect 1719 27489 1731 27492
rect 1673 27483 1731 27489
rect 3326 27480 3332 27492
rect 3384 27480 3390 27532
rect 48314 27480 48320 27532
rect 48372 27520 48378 27532
rect 48593 27523 48651 27529
rect 48593 27520 48605 27523
rect 48372 27492 48605 27520
rect 48372 27480 48378 27492
rect 48593 27489 48605 27492
rect 48639 27489 48651 27523
rect 49050 27520 49056 27532
rect 49011 27492 49056 27520
rect 48593 27483 48651 27489
rect 49050 27480 49056 27492
rect 49108 27480 49114 27532
rect 49252 27529 49280 27560
rect 50246 27548 50252 27560
rect 50304 27548 50310 27600
rect 49237 27523 49295 27529
rect 49237 27489 49249 27523
rect 49283 27489 49295 27523
rect 49237 27483 49295 27489
rect 49881 27523 49939 27529
rect 49881 27489 49893 27523
rect 49927 27520 49939 27523
rect 49970 27520 49976 27532
rect 49927 27492 49976 27520
rect 49927 27489 49939 27492
rect 49881 27483 49939 27489
rect 49970 27480 49976 27492
rect 50028 27520 50034 27532
rect 50154 27520 50160 27532
rect 50028 27492 50160 27520
rect 50028 27480 50034 27492
rect 50154 27480 50160 27492
rect 50212 27480 50218 27532
rect 50341 27523 50399 27529
rect 50341 27489 50353 27523
rect 50387 27489 50399 27523
rect 50448 27520 50476 27628
rect 50525 27625 50537 27659
rect 50571 27656 50583 27659
rect 50571 27628 51028 27656
rect 50571 27625 50583 27628
rect 50525 27619 50583 27625
rect 51000 27588 51028 27628
rect 51258 27616 51264 27668
rect 51316 27656 51322 27668
rect 51445 27659 51503 27665
rect 51445 27656 51457 27659
rect 51316 27628 51457 27656
rect 51316 27616 51322 27628
rect 51445 27625 51457 27628
rect 51491 27625 51503 27659
rect 53466 27656 53472 27668
rect 53427 27628 53472 27656
rect 51445 27619 51503 27625
rect 53466 27616 53472 27628
rect 53524 27616 53530 27668
rect 52730 27588 52736 27600
rect 51000 27560 51672 27588
rect 51644 27529 51672 27560
rect 52564 27560 52736 27588
rect 50525 27523 50583 27529
rect 50525 27520 50537 27523
rect 50448 27492 50537 27520
rect 50341 27483 50399 27489
rect 50525 27489 50537 27492
rect 50571 27489 50583 27523
rect 50525 27483 50583 27489
rect 51629 27523 51687 27529
rect 51629 27489 51641 27523
rect 51675 27520 51687 27523
rect 51718 27520 51724 27532
rect 51675 27492 51724 27520
rect 51675 27489 51687 27492
rect 51629 27483 51687 27489
rect 1857 27455 1915 27461
rect 1857 27421 1869 27455
rect 1903 27452 1915 27455
rect 2498 27452 2504 27464
rect 1903 27424 2504 27452
rect 1903 27421 1915 27424
rect 1857 27415 1915 27421
rect 2498 27412 2504 27424
rect 2556 27412 2562 27464
rect 50356 27452 50384 27483
rect 51718 27480 51724 27492
rect 51776 27480 51782 27532
rect 51810 27480 51816 27532
rect 51868 27520 51874 27532
rect 52564 27529 52592 27560
rect 52730 27548 52736 27560
rect 52788 27548 52794 27600
rect 52822 27548 52828 27600
rect 52880 27548 52886 27600
rect 54113 27591 54171 27597
rect 54113 27557 54125 27591
rect 54159 27557 54171 27591
rect 55214 27588 55220 27600
rect 54113 27551 54171 27557
rect 54404 27560 55220 27588
rect 51905 27523 51963 27529
rect 51905 27520 51917 27523
rect 51868 27492 51917 27520
rect 51868 27480 51874 27492
rect 51905 27489 51917 27492
rect 51951 27489 51963 27523
rect 51905 27483 51963 27489
rect 52549 27523 52607 27529
rect 52549 27489 52561 27523
rect 52595 27489 52607 27523
rect 52549 27483 52607 27489
rect 52641 27523 52699 27529
rect 52641 27489 52653 27523
rect 52687 27520 52699 27523
rect 52840 27520 52868 27548
rect 53377 27523 53435 27529
rect 53377 27520 53389 27523
rect 52687 27492 53389 27520
rect 52687 27489 52699 27492
rect 52641 27483 52699 27489
rect 53377 27489 53389 27492
rect 53423 27520 53435 27523
rect 54128 27520 54156 27551
rect 54294 27520 54300 27532
rect 53423 27492 54156 27520
rect 54255 27492 54300 27520
rect 53423 27489 53435 27492
rect 53377 27483 53435 27489
rect 54294 27480 54300 27492
rect 54352 27480 54358 27532
rect 54404 27529 54432 27560
rect 55214 27548 55220 27560
rect 55272 27548 55278 27600
rect 57054 27588 57060 27600
rect 57015 27560 57060 27588
rect 57054 27548 57060 27560
rect 57112 27548 57118 27600
rect 54389 27523 54447 27529
rect 54389 27489 54401 27523
rect 54435 27489 54447 27523
rect 54662 27520 54668 27532
rect 54623 27492 54668 27520
rect 54389 27483 54447 27489
rect 54662 27480 54668 27492
rect 54720 27480 54726 27532
rect 55306 27520 55312 27532
rect 55267 27492 55312 27520
rect 55306 27480 55312 27492
rect 55364 27480 55370 27532
rect 55490 27520 55496 27532
rect 55451 27492 55496 27520
rect 55490 27480 55496 27492
rect 55548 27480 55554 27532
rect 55674 27520 55680 27532
rect 55635 27492 55680 27520
rect 55674 27480 55680 27492
rect 55732 27480 55738 27532
rect 56873 27523 56931 27529
rect 56873 27489 56885 27523
rect 56919 27520 56931 27523
rect 58161 27523 58219 27529
rect 58161 27520 58173 27523
rect 56919 27492 58173 27520
rect 56919 27489 56931 27492
rect 56873 27483 56931 27489
rect 58161 27489 58173 27492
rect 58207 27489 58219 27523
rect 58161 27483 58219 27489
rect 51166 27452 51172 27464
rect 50356 27424 51172 27452
rect 51166 27412 51172 27424
rect 51224 27412 51230 27464
rect 52730 27452 52736 27464
rect 52691 27424 52736 27452
rect 52730 27412 52736 27424
rect 52788 27412 52794 27464
rect 52825 27455 52883 27461
rect 52825 27421 52837 27455
rect 52871 27452 52883 27455
rect 54110 27452 54116 27464
rect 52871 27424 54116 27452
rect 52871 27421 52883 27424
rect 52825 27415 52883 27421
rect 54110 27412 54116 27424
rect 54168 27412 54174 27464
rect 54202 27412 54208 27464
rect 54260 27452 54266 27464
rect 54570 27452 54576 27464
rect 54260 27424 54576 27452
rect 54260 27412 54266 27424
rect 54570 27412 54576 27424
rect 54628 27412 54634 27464
rect 57517 27455 57575 27461
rect 57517 27421 57529 27455
rect 57563 27421 57575 27455
rect 57698 27452 57704 27464
rect 57659 27424 57704 27452
rect 57517 27415 57575 27421
rect 2038 27384 2044 27396
rect 1999 27356 2044 27384
rect 2038 27344 2044 27356
rect 2096 27344 2102 27396
rect 53006 27384 53012 27396
rect 52656 27356 53012 27384
rect 52656 27328 52684 27356
rect 53006 27344 53012 27356
rect 53064 27344 53070 27396
rect 53190 27344 53196 27396
rect 53248 27384 53254 27396
rect 55309 27387 55367 27393
rect 55309 27384 55321 27387
rect 53248 27356 55321 27384
rect 53248 27344 53254 27356
rect 55309 27353 55321 27356
rect 55355 27353 55367 27387
rect 55309 27347 55367 27353
rect 48406 27316 48412 27328
rect 48367 27288 48412 27316
rect 48406 27276 48412 27288
rect 48464 27276 48470 27328
rect 49053 27319 49111 27325
rect 49053 27285 49065 27319
rect 49099 27316 49111 27319
rect 49602 27316 49608 27328
rect 49099 27288 49608 27316
rect 49099 27285 49111 27288
rect 49053 27279 49111 27285
rect 49602 27276 49608 27288
rect 49660 27276 49666 27328
rect 49697 27319 49755 27325
rect 49697 27285 49709 27319
rect 49743 27316 49755 27319
rect 51626 27316 51632 27328
rect 49743 27288 51632 27316
rect 49743 27285 49755 27288
rect 49697 27279 49755 27285
rect 51626 27276 51632 27288
rect 51684 27276 51690 27328
rect 51813 27319 51871 27325
rect 51813 27285 51825 27319
rect 51859 27316 51871 27319
rect 51994 27316 52000 27328
rect 51859 27288 52000 27316
rect 51859 27285 51871 27288
rect 51813 27279 51871 27285
rect 51994 27276 52000 27288
rect 52052 27276 52058 27328
rect 52362 27316 52368 27328
rect 52323 27288 52368 27316
rect 52362 27276 52368 27288
rect 52420 27276 52426 27328
rect 52638 27276 52644 27328
rect 52696 27276 52702 27328
rect 52822 27276 52828 27328
rect 52880 27316 52886 27328
rect 57532 27316 57560 27415
rect 57698 27412 57704 27424
rect 57756 27412 57762 27464
rect 52880 27288 57560 27316
rect 52880 27276 52886 27288
rect 1104 27226 58880 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 58880 27226
rect 1104 27152 58880 27174
rect 2498 27112 2504 27124
rect 2459 27084 2504 27112
rect 2498 27072 2504 27084
rect 2556 27072 2562 27124
rect 3326 27112 3332 27124
rect 3287 27084 3332 27112
rect 3326 27072 3332 27084
rect 3384 27072 3390 27124
rect 49878 27072 49884 27124
rect 49936 27112 49942 27124
rect 49936 27084 51074 27112
rect 49936 27072 49942 27084
rect 51046 26920 51074 27084
rect 51626 27072 51632 27124
rect 51684 27112 51690 27124
rect 54110 27112 54116 27124
rect 51684 27084 52868 27112
rect 54071 27084 54116 27112
rect 51684 27072 51690 27084
rect 52730 27004 52736 27056
rect 52788 27004 52794 27056
rect 52840 27044 52868 27084
rect 54110 27072 54116 27084
rect 54168 27072 54174 27124
rect 55309 27115 55367 27121
rect 55309 27081 55321 27115
rect 55355 27112 55367 27115
rect 55674 27112 55680 27124
rect 55355 27084 55680 27112
rect 55355 27081 55367 27084
rect 55309 27075 55367 27081
rect 55674 27072 55680 27084
rect 55732 27072 55738 27124
rect 57238 27044 57244 27056
rect 52840 27016 57244 27044
rect 57238 27004 57244 27016
rect 57296 27004 57302 27056
rect 51166 26936 51172 26988
rect 51224 26976 51230 26988
rect 52362 26976 52368 26988
rect 51224 26948 52368 26976
rect 51224 26936 51230 26948
rect 2682 26908 2688 26920
rect 2595 26880 2688 26908
rect 2682 26868 2688 26880
rect 2740 26908 2746 26920
rect 2866 26908 2872 26920
rect 2740 26880 2872 26908
rect 2740 26868 2746 26880
rect 2866 26868 2872 26880
rect 2924 26868 2930 26920
rect 49234 26908 49240 26920
rect 49195 26880 49240 26908
rect 49234 26868 49240 26880
rect 49292 26868 49298 26920
rect 50982 26868 50988 26920
rect 51040 26908 51074 26920
rect 51460 26917 51488 26948
rect 52362 26936 52368 26948
rect 52420 26936 52426 26988
rect 52549 26979 52607 26985
rect 52549 26945 52561 26979
rect 52595 26976 52607 26979
rect 52748 26976 52776 27004
rect 53101 26979 53159 26985
rect 53101 26976 53113 26979
rect 52595 26948 53113 26976
rect 52595 26945 52607 26948
rect 52549 26939 52607 26945
rect 53101 26945 53113 26948
rect 53147 26976 53159 26979
rect 54202 26976 54208 26988
rect 53147 26948 54208 26976
rect 53147 26945 53159 26948
rect 53101 26939 53159 26945
rect 54202 26936 54208 26948
rect 54260 26936 54266 26988
rect 55214 26976 55220 26988
rect 54772 26948 55220 26976
rect 51353 26911 51411 26917
rect 51353 26908 51365 26911
rect 51040 26880 51365 26908
rect 51040 26868 51046 26880
rect 51353 26877 51365 26880
rect 51399 26877 51411 26911
rect 51353 26871 51411 26877
rect 51442 26911 51500 26917
rect 51442 26877 51454 26911
rect 51488 26877 51500 26911
rect 51442 26871 51500 26877
rect 51537 26911 51595 26917
rect 51537 26877 51549 26911
rect 51583 26877 51595 26911
rect 51718 26908 51724 26920
rect 51679 26880 51724 26908
rect 51537 26871 51595 26877
rect 1857 26843 1915 26849
rect 1857 26809 1869 26843
rect 1903 26840 1915 26843
rect 2314 26840 2320 26852
rect 1903 26812 2320 26840
rect 1903 26809 1915 26812
rect 1857 26803 1915 26809
rect 2314 26800 2320 26812
rect 2372 26800 2378 26852
rect 49504 26843 49562 26849
rect 49504 26809 49516 26843
rect 49550 26840 49562 26843
rect 51077 26843 51135 26849
rect 51077 26840 51089 26843
rect 49550 26812 51089 26840
rect 49550 26809 49562 26812
rect 49504 26803 49562 26809
rect 51077 26809 51089 26812
rect 51123 26809 51135 26843
rect 51552 26840 51580 26871
rect 51718 26868 51724 26880
rect 51776 26868 51782 26920
rect 52733 26911 52791 26917
rect 52733 26877 52745 26911
rect 52779 26908 52791 26911
rect 53006 26908 53012 26920
rect 52779 26880 53012 26908
rect 52779 26877 52791 26880
rect 52733 26871 52791 26877
rect 53006 26868 53012 26880
rect 53064 26868 53070 26920
rect 53190 26868 53196 26920
rect 53248 26908 53254 26920
rect 54772 26917 54800 26948
rect 55214 26936 55220 26948
rect 55272 26976 55278 26988
rect 55272 26948 56180 26976
rect 55272 26936 55278 26948
rect 54021 26911 54079 26917
rect 54021 26908 54033 26911
rect 53248 26880 54033 26908
rect 53248 26868 53254 26880
rect 54021 26877 54033 26880
rect 54067 26877 54079 26911
rect 54021 26871 54079 26877
rect 54757 26911 54815 26917
rect 54757 26877 54769 26911
rect 54803 26877 54815 26911
rect 54757 26871 54815 26877
rect 55125 26911 55183 26917
rect 55125 26877 55137 26911
rect 55171 26908 55183 26911
rect 55306 26908 55312 26920
rect 55171 26880 55312 26908
rect 55171 26877 55183 26880
rect 55125 26871 55183 26877
rect 55306 26868 55312 26880
rect 55364 26868 55370 26920
rect 56152 26917 56180 26948
rect 56137 26911 56195 26917
rect 56137 26877 56149 26911
rect 56183 26908 56195 26911
rect 56502 26908 56508 26920
rect 56183 26880 56508 26908
rect 56183 26877 56195 26880
rect 56137 26871 56195 26877
rect 56502 26868 56508 26880
rect 56560 26868 56566 26920
rect 57146 26908 57152 26920
rect 57107 26880 57152 26908
rect 57146 26868 57152 26880
rect 57204 26868 57210 26920
rect 57333 26911 57391 26917
rect 57333 26877 57345 26911
rect 57379 26877 57391 26911
rect 57333 26871 57391 26877
rect 52638 26840 52644 26852
rect 51552 26812 52644 26840
rect 51077 26803 51135 26809
rect 52638 26800 52644 26812
rect 52696 26800 52702 26852
rect 53926 26840 53932 26852
rect 52932 26812 53932 26840
rect 1946 26772 1952 26784
rect 1907 26744 1952 26772
rect 1946 26732 1952 26744
rect 2004 26732 2010 26784
rect 50614 26772 50620 26784
rect 50575 26744 50620 26772
rect 50614 26732 50620 26744
rect 50672 26732 50678 26784
rect 52932 26781 52960 26812
rect 53926 26800 53932 26812
rect 53984 26800 53990 26852
rect 54294 26800 54300 26852
rect 54352 26840 54358 26852
rect 54941 26843 54999 26849
rect 54941 26840 54953 26843
rect 54352 26812 54953 26840
rect 54352 26800 54358 26812
rect 54941 26809 54953 26812
rect 54987 26809 54999 26843
rect 54941 26803 54999 26809
rect 55030 26800 55036 26852
rect 55088 26840 55094 26852
rect 55088 26812 55133 26840
rect 55088 26800 55094 26812
rect 55214 26800 55220 26852
rect 55272 26840 55278 26852
rect 57348 26840 57376 26871
rect 55272 26812 57376 26840
rect 55272 26800 55278 26812
rect 52917 26775 52975 26781
rect 52917 26741 52929 26775
rect 52963 26741 52975 26775
rect 52917 26735 52975 26741
rect 53006 26732 53012 26784
rect 53064 26772 53070 26784
rect 54018 26772 54024 26784
rect 53064 26744 54024 26772
rect 53064 26732 53070 26744
rect 54018 26732 54024 26744
rect 54076 26732 54082 26784
rect 54570 26732 54576 26784
rect 54628 26772 54634 26784
rect 56229 26775 56287 26781
rect 56229 26772 56241 26775
rect 54628 26744 56241 26772
rect 54628 26732 54634 26744
rect 56229 26741 56241 26744
rect 56275 26741 56287 26775
rect 56229 26735 56287 26741
rect 57238 26732 57244 26784
rect 57296 26772 57302 26784
rect 57793 26775 57851 26781
rect 57793 26772 57805 26775
rect 57296 26744 57805 26772
rect 57296 26732 57302 26744
rect 57793 26741 57805 26744
rect 57839 26741 57851 26775
rect 57793 26735 57851 26741
rect 1104 26682 58880 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 50326 26682
rect 50378 26630 50390 26682
rect 50442 26630 50454 26682
rect 50506 26630 50518 26682
rect 50570 26630 58880 26682
rect 1104 26608 58880 26630
rect 2314 26568 2320 26580
rect 2275 26540 2320 26568
rect 2314 26528 2320 26540
rect 2372 26528 2378 26580
rect 49697 26571 49755 26577
rect 49697 26537 49709 26571
rect 49743 26537 49755 26571
rect 49697 26531 49755 26537
rect 49712 26500 49740 26531
rect 50982 26528 50988 26580
rect 51040 26568 51046 26580
rect 51445 26571 51503 26577
rect 51445 26568 51457 26571
rect 51040 26540 51457 26568
rect 51040 26528 51046 26540
rect 51445 26537 51457 26540
rect 51491 26537 51503 26571
rect 51445 26531 51503 26537
rect 54294 26528 54300 26580
rect 54352 26568 54358 26580
rect 55030 26568 55036 26580
rect 54352 26540 55036 26568
rect 54352 26528 54358 26540
rect 55030 26528 55036 26540
rect 55088 26568 55094 26580
rect 55490 26568 55496 26580
rect 55088 26540 55496 26568
rect 55088 26528 55094 26540
rect 55490 26528 55496 26540
rect 55548 26528 55554 26580
rect 57330 26568 57336 26580
rect 57291 26540 57336 26568
rect 57330 26528 57336 26540
rect 57388 26528 57394 26580
rect 55214 26500 55220 26512
rect 49712 26472 55220 26500
rect 55214 26460 55220 26472
rect 55272 26460 55278 26512
rect 1673 26435 1731 26441
rect 1673 26401 1685 26435
rect 1719 26432 1731 26435
rect 2961 26435 3019 26441
rect 2961 26432 2973 26435
rect 1719 26404 2973 26432
rect 1719 26401 1731 26404
rect 1673 26395 1731 26401
rect 2961 26401 2973 26404
rect 3007 26401 3019 26435
rect 2961 26395 3019 26401
rect 49881 26435 49939 26441
rect 49881 26401 49893 26435
rect 49927 26432 49939 26435
rect 49970 26432 49976 26444
rect 49927 26404 49976 26432
rect 49927 26401 49939 26404
rect 49881 26395 49939 26401
rect 49970 26392 49976 26404
rect 50028 26392 50034 26444
rect 50341 26435 50399 26441
rect 50341 26401 50353 26435
rect 50387 26432 50399 26435
rect 50614 26432 50620 26444
rect 50387 26404 50620 26432
rect 50387 26401 50399 26404
rect 50341 26395 50399 26401
rect 50614 26392 50620 26404
rect 50672 26432 50678 26444
rect 51629 26435 51687 26441
rect 51629 26432 51641 26435
rect 50672 26404 51641 26432
rect 50672 26392 50678 26404
rect 51629 26401 51641 26404
rect 51675 26401 51687 26435
rect 51629 26395 51687 26401
rect 51718 26392 51724 26444
rect 51776 26432 51782 26444
rect 51776 26404 51821 26432
rect 51776 26392 51782 26404
rect 51902 26392 51908 26444
rect 51960 26432 51966 26444
rect 51997 26435 52055 26441
rect 51997 26432 52009 26435
rect 51960 26404 52009 26432
rect 51960 26392 51966 26404
rect 51997 26401 52009 26404
rect 52043 26401 52055 26435
rect 52914 26432 52920 26444
rect 52875 26404 52920 26432
rect 51997 26395 52055 26401
rect 52914 26392 52920 26404
rect 52972 26392 52978 26444
rect 53184 26435 53242 26441
rect 53184 26401 53196 26435
rect 53230 26432 53242 26435
rect 54110 26432 54116 26444
rect 53230 26404 54116 26432
rect 53230 26401 53242 26404
rect 53184 26395 53242 26401
rect 54110 26392 54116 26404
rect 54168 26392 54174 26444
rect 54386 26392 54392 26444
rect 54444 26432 54450 26444
rect 54941 26435 54999 26441
rect 54941 26432 54953 26435
rect 54444 26404 54953 26432
rect 54444 26392 54450 26404
rect 54941 26401 54953 26404
rect 54987 26401 54999 26435
rect 54941 26395 54999 26401
rect 55033 26435 55091 26441
rect 55033 26401 55045 26435
rect 55079 26401 55091 26435
rect 55033 26395 55091 26401
rect 55309 26435 55367 26441
rect 55309 26401 55321 26435
rect 55355 26432 55367 26435
rect 55508 26432 55536 26528
rect 57238 26500 57244 26512
rect 57199 26472 57244 26500
rect 57238 26460 57244 26472
rect 57296 26460 57302 26512
rect 57974 26432 57980 26444
rect 55355 26404 55536 26432
rect 57935 26404 57980 26432
rect 55355 26401 55367 26404
rect 55309 26395 55367 26401
rect 1854 26364 1860 26376
rect 1815 26336 1860 26364
rect 1854 26324 1860 26336
rect 1912 26324 1918 26376
rect 50154 26324 50160 26376
rect 50212 26364 50218 26376
rect 50433 26367 50491 26373
rect 50433 26364 50445 26367
rect 50212 26336 50445 26364
rect 50212 26324 50218 26336
rect 50433 26333 50445 26336
rect 50479 26364 50491 26367
rect 51920 26364 51948 26392
rect 50479 26336 51948 26364
rect 50479 26333 50491 26336
rect 50433 26327 50491 26333
rect 54202 26324 54208 26376
rect 54260 26364 54266 26376
rect 54757 26367 54815 26373
rect 54757 26364 54769 26367
rect 54260 26336 54769 26364
rect 54260 26324 54266 26336
rect 54757 26333 54769 26336
rect 54803 26333 54815 26367
rect 54757 26327 54815 26333
rect 54846 26324 54852 26376
rect 54904 26364 54910 26376
rect 55048 26364 55076 26395
rect 57974 26392 57980 26404
rect 58032 26392 58038 26444
rect 54904 26336 55076 26364
rect 54904 26324 54910 26336
rect 49237 26299 49295 26305
rect 49237 26265 49249 26299
rect 49283 26296 49295 26299
rect 52822 26296 52828 26308
rect 49283 26268 52828 26296
rect 49283 26265 49295 26268
rect 49237 26259 49295 26265
rect 52822 26256 52828 26268
rect 52880 26256 52886 26308
rect 55490 26296 55496 26308
rect 53852 26268 55496 26296
rect 49418 26188 49424 26240
rect 49476 26228 49482 26240
rect 51810 26228 51816 26240
rect 49476 26200 51816 26228
rect 49476 26188 49482 26200
rect 51810 26188 51816 26200
rect 51868 26188 51874 26240
rect 51905 26231 51963 26237
rect 51905 26197 51917 26231
rect 51951 26228 51963 26231
rect 51994 26228 52000 26240
rect 51951 26200 52000 26228
rect 51951 26197 51963 26200
rect 51905 26191 51963 26197
rect 51994 26188 52000 26200
rect 52052 26188 52058 26240
rect 52454 26188 52460 26240
rect 52512 26228 52518 26240
rect 53852 26228 53880 26268
rect 55490 26256 55496 26268
rect 55548 26256 55554 26308
rect 57882 26256 57888 26308
rect 57940 26296 57946 26308
rect 58161 26299 58219 26305
rect 58161 26296 58173 26299
rect 57940 26268 58173 26296
rect 57940 26256 57946 26268
rect 58161 26265 58173 26268
rect 58207 26265 58219 26299
rect 58161 26259 58219 26265
rect 52512 26200 53880 26228
rect 55217 26231 55275 26237
rect 52512 26188 52518 26200
rect 55217 26197 55229 26231
rect 55263 26228 55275 26231
rect 55306 26228 55312 26240
rect 55263 26200 55312 26228
rect 55263 26197 55275 26200
rect 55217 26191 55275 26197
rect 55306 26188 55312 26200
rect 55364 26228 55370 26240
rect 56318 26228 56324 26240
rect 55364 26200 56324 26228
rect 55364 26188 55370 26200
rect 56318 26188 56324 26200
rect 56376 26188 56382 26240
rect 1104 26138 58880 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 58880 26138
rect 1104 26064 58880 26086
rect 1854 25984 1860 26036
rect 1912 26024 1918 26036
rect 2501 26027 2559 26033
rect 2501 26024 2513 26027
rect 1912 25996 2513 26024
rect 1912 25984 1918 25996
rect 2501 25993 2513 25996
rect 2547 25993 2559 26027
rect 46198 26024 46204 26036
rect 2501 25987 2559 25993
rect 6886 25996 46204 26024
rect 1302 25916 1308 25968
rect 1360 25956 1366 25968
rect 6886 25956 6914 25996
rect 46198 25984 46204 25996
rect 46256 25984 46262 26036
rect 49234 25984 49240 26036
rect 49292 26024 49298 26036
rect 50614 26024 50620 26036
rect 49292 25996 50620 26024
rect 49292 25984 49298 25996
rect 50614 25984 50620 25996
rect 50672 25984 50678 26036
rect 51718 25984 51724 26036
rect 51776 26024 51782 26036
rect 51997 26027 52055 26033
rect 51997 26024 52009 26027
rect 51776 25996 52009 26024
rect 51776 25984 51782 25996
rect 51997 25993 52009 25996
rect 52043 25993 52055 26027
rect 51997 25987 52055 25993
rect 1360 25928 6914 25956
rect 1360 25916 1366 25928
rect 49988 25860 50752 25888
rect 2685 25823 2743 25829
rect 2685 25789 2697 25823
rect 2731 25789 2743 25823
rect 2685 25783 2743 25789
rect 1854 25752 1860 25764
rect 1815 25724 1860 25752
rect 1854 25712 1860 25724
rect 1912 25712 1918 25764
rect 2038 25752 2044 25764
rect 1999 25724 2044 25752
rect 2038 25712 2044 25724
rect 2096 25712 2102 25764
rect 2700 25752 2728 25783
rect 2774 25780 2780 25832
rect 2832 25820 2838 25832
rect 49988 25829 50016 25860
rect 3329 25823 3387 25829
rect 3329 25820 3341 25823
rect 2832 25792 3341 25820
rect 2832 25780 2838 25792
rect 3329 25789 3341 25792
rect 3375 25789 3387 25823
rect 3329 25783 3387 25789
rect 49329 25823 49387 25829
rect 49329 25789 49341 25823
rect 49375 25789 49387 25823
rect 49329 25783 49387 25789
rect 49973 25823 50031 25829
rect 49973 25789 49985 25823
rect 50019 25789 50031 25823
rect 50154 25820 50160 25832
rect 50115 25792 50160 25820
rect 49973 25783 50031 25789
rect 3142 25752 3148 25764
rect 2700 25724 3148 25752
rect 3142 25712 3148 25724
rect 3200 25712 3206 25764
rect 49344 25684 49372 25783
rect 50154 25780 50160 25792
rect 50212 25780 50218 25832
rect 50614 25820 50620 25832
rect 50575 25792 50620 25820
rect 50614 25780 50620 25792
rect 50672 25780 50678 25832
rect 50724 25820 50752 25860
rect 52012 25820 52040 25987
rect 52086 25984 52092 26036
rect 52144 26024 52150 26036
rect 52549 26027 52607 26033
rect 52549 26024 52561 26027
rect 52144 25996 52561 26024
rect 52144 25984 52150 25996
rect 52549 25993 52561 25996
rect 52595 25993 52607 26027
rect 57146 26024 57152 26036
rect 52549 25987 52607 25993
rect 52656 25996 57152 26024
rect 52086 25848 52092 25900
rect 52144 25888 52150 25900
rect 52656 25888 52684 25996
rect 57146 25984 57152 25996
rect 57204 25984 57210 26036
rect 57974 26024 57980 26036
rect 57935 25996 57980 26024
rect 57974 25984 57980 25996
rect 58032 25984 58038 26036
rect 56318 25956 56324 25968
rect 56231 25928 56324 25956
rect 56318 25916 56324 25928
rect 56376 25956 56382 25968
rect 56376 25928 56824 25956
rect 56376 25916 56382 25928
rect 52144 25860 52684 25888
rect 52144 25848 52150 25860
rect 52730 25848 52736 25900
rect 52788 25888 52794 25900
rect 56594 25888 56600 25900
rect 52788 25860 55070 25888
rect 52788 25848 52794 25860
rect 52457 25823 52515 25829
rect 52457 25820 52469 25823
rect 50724 25792 51074 25820
rect 52012 25792 52469 25820
rect 51046 25764 51074 25792
rect 52457 25789 52469 25792
rect 52503 25789 52515 25823
rect 54294 25820 54300 25832
rect 54255 25792 54300 25820
rect 52457 25783 52515 25789
rect 54294 25780 54300 25792
rect 54352 25780 54358 25832
rect 54754 25780 54760 25832
rect 54812 25820 54818 25832
rect 54941 25823 54999 25829
rect 54941 25820 54953 25823
rect 54812 25792 54953 25820
rect 54812 25780 54818 25792
rect 54941 25789 54953 25792
rect 54987 25789 54999 25823
rect 55042 25820 55070 25860
rect 55968 25860 56600 25888
rect 55968 25820 55996 25860
rect 56594 25848 56600 25860
rect 56652 25848 56658 25900
rect 56796 25829 56824 25928
rect 55042 25792 55996 25820
rect 56781 25823 56839 25829
rect 54941 25783 54999 25789
rect 56781 25789 56793 25823
rect 56827 25789 56839 25823
rect 56781 25783 56839 25789
rect 57517 25823 57575 25829
rect 57517 25789 57529 25823
rect 57563 25789 57575 25823
rect 57698 25820 57704 25832
rect 57659 25792 57704 25820
rect 57517 25783 57575 25789
rect 50065 25755 50123 25761
rect 50065 25721 50077 25755
rect 50111 25752 50123 25755
rect 50862 25755 50920 25761
rect 50862 25752 50874 25755
rect 50111 25724 50874 25752
rect 50111 25721 50123 25724
rect 50065 25715 50123 25721
rect 50862 25721 50874 25724
rect 50908 25721 50920 25755
rect 51046 25724 51080 25764
rect 50862 25715 50920 25721
rect 51074 25712 51080 25724
rect 51132 25712 51138 25764
rect 51626 25712 51632 25764
rect 51684 25752 51690 25764
rect 54846 25752 54852 25764
rect 51684 25724 54852 25752
rect 51684 25712 51690 25724
rect 54846 25712 54852 25724
rect 54904 25712 54910 25764
rect 54956 25752 54984 25783
rect 55030 25752 55036 25764
rect 54956 25724 55036 25752
rect 55030 25712 55036 25724
rect 55088 25712 55094 25764
rect 55122 25712 55128 25764
rect 55180 25761 55186 25764
rect 55180 25755 55244 25761
rect 55180 25721 55198 25755
rect 55232 25721 55244 25755
rect 55180 25715 55244 25721
rect 55180 25712 55186 25715
rect 55306 25712 55312 25764
rect 55364 25752 55370 25764
rect 57532 25752 57560 25783
rect 57698 25780 57704 25792
rect 57756 25780 57762 25832
rect 55364 25724 57560 25752
rect 55364 25712 55370 25724
rect 52454 25684 52460 25696
rect 49344 25656 52460 25684
rect 52454 25644 52460 25656
rect 52512 25644 52518 25696
rect 54386 25684 54392 25696
rect 54347 25656 54392 25684
rect 54386 25644 54392 25656
rect 54444 25644 54450 25696
rect 54864 25684 54892 25712
rect 56873 25687 56931 25693
rect 56873 25684 56885 25687
rect 54864 25656 56885 25684
rect 56873 25653 56885 25656
rect 56919 25653 56931 25687
rect 56873 25647 56931 25653
rect 1104 25594 58880 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 50326 25594
rect 50378 25542 50390 25594
rect 50442 25542 50454 25594
rect 50506 25542 50518 25594
rect 50570 25542 58880 25594
rect 1104 25520 58880 25542
rect 1854 25440 1860 25492
rect 1912 25480 1918 25492
rect 2501 25483 2559 25489
rect 2501 25480 2513 25483
rect 1912 25452 2513 25480
rect 1912 25440 1918 25452
rect 2501 25449 2513 25452
rect 2547 25449 2559 25483
rect 2501 25443 2559 25449
rect 51810 25440 51816 25492
rect 51868 25480 51874 25492
rect 54113 25483 54171 25489
rect 54113 25480 54125 25483
rect 51868 25452 54125 25480
rect 51868 25440 51874 25452
rect 54113 25449 54125 25452
rect 54159 25449 54171 25483
rect 55122 25480 55128 25492
rect 55083 25452 55128 25480
rect 54113 25443 54171 25449
rect 55122 25440 55128 25452
rect 55180 25440 55186 25492
rect 46198 25372 46204 25424
rect 46256 25412 46262 25424
rect 52825 25415 52883 25421
rect 52825 25412 52837 25415
rect 46256 25384 52837 25412
rect 46256 25372 46262 25384
rect 52825 25381 52837 25384
rect 52871 25381 52883 25415
rect 52825 25375 52883 25381
rect 54386 25372 54392 25424
rect 54444 25412 54450 25424
rect 58158 25412 58164 25424
rect 54444 25384 55260 25412
rect 58119 25384 58164 25412
rect 54444 25372 54450 25384
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 2774 25344 2780 25356
rect 1903 25316 2780 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 2774 25304 2780 25316
rect 2832 25304 2838 25356
rect 3142 25344 3148 25356
rect 3103 25316 3148 25344
rect 3142 25304 3148 25316
rect 3200 25304 3206 25356
rect 49050 25304 49056 25356
rect 49108 25344 49114 25356
rect 50341 25347 50399 25353
rect 50341 25344 50353 25347
rect 49108 25316 50353 25344
rect 49108 25304 49114 25316
rect 50341 25313 50353 25316
rect 50387 25313 50399 25347
rect 50341 25307 50399 25313
rect 50525 25347 50583 25353
rect 50525 25313 50537 25347
rect 50571 25344 50583 25347
rect 51626 25344 51632 25356
rect 50571 25316 51632 25344
rect 50571 25313 50583 25316
rect 50525 25307 50583 25313
rect 51626 25304 51632 25316
rect 51684 25304 51690 25356
rect 51721 25347 51779 25353
rect 51721 25313 51733 25347
rect 51767 25344 51779 25347
rect 51994 25344 52000 25356
rect 51767 25316 52000 25344
rect 51767 25313 51779 25316
rect 51721 25307 51779 25313
rect 51994 25304 52000 25316
rect 52052 25344 52058 25356
rect 52365 25347 52423 25353
rect 52365 25344 52377 25347
rect 52052 25316 52377 25344
rect 52052 25304 52058 25316
rect 52365 25313 52377 25316
rect 52411 25313 52423 25347
rect 52365 25307 52423 25313
rect 54938 25304 54944 25356
rect 54996 25344 55002 25356
rect 55232 25353 55260 25384
rect 58158 25372 58164 25384
rect 58216 25372 58222 25424
rect 55033 25347 55091 25353
rect 55033 25344 55045 25347
rect 54996 25316 55045 25344
rect 54996 25304 55002 25316
rect 55033 25313 55045 25316
rect 55079 25313 55091 25347
rect 55033 25307 55091 25313
rect 55217 25347 55275 25353
rect 55217 25313 55229 25347
rect 55263 25313 55275 25347
rect 55217 25307 55275 25313
rect 56686 25304 56692 25356
rect 56744 25344 56750 25356
rect 56781 25347 56839 25353
rect 56781 25344 56793 25347
rect 56744 25316 56793 25344
rect 56744 25304 56750 25316
rect 56781 25313 56793 25316
rect 56827 25313 56839 25347
rect 56781 25307 56839 25313
rect 57425 25347 57483 25353
rect 57425 25313 57437 25347
rect 57471 25344 57483 25347
rect 57977 25347 58035 25353
rect 57977 25344 57989 25347
rect 57471 25316 57989 25344
rect 57471 25313 57483 25316
rect 57425 25307 57483 25313
rect 57977 25313 57989 25316
rect 58023 25313 58035 25347
rect 57977 25307 58035 25313
rect 2041 25279 2099 25285
rect 2041 25245 2053 25279
rect 2087 25245 2099 25279
rect 2041 25239 2099 25245
rect 49881 25279 49939 25285
rect 49881 25245 49893 25279
rect 49927 25276 49939 25279
rect 55306 25276 55312 25288
rect 49927 25248 55312 25276
rect 49927 25245 49939 25248
rect 49881 25239 49939 25245
rect 2056 25208 2084 25239
rect 55306 25236 55312 25248
rect 55364 25236 55370 25288
rect 56965 25279 57023 25285
rect 56965 25245 56977 25279
rect 57011 25245 57023 25279
rect 56965 25239 57023 25245
rect 2961 25211 3019 25217
rect 2961 25208 2973 25211
rect 2056 25180 2973 25208
rect 2961 25177 2973 25180
rect 3007 25177 3019 25211
rect 2961 25171 3019 25177
rect 51537 25211 51595 25217
rect 51537 25177 51549 25211
rect 51583 25208 51595 25211
rect 51583 25180 53604 25208
rect 51583 25177 51595 25180
rect 51537 25171 51595 25177
rect 50341 25143 50399 25149
rect 50341 25109 50353 25143
rect 50387 25140 50399 25143
rect 52086 25140 52092 25152
rect 50387 25112 52092 25140
rect 50387 25109 50399 25112
rect 50341 25103 50399 25109
rect 52086 25100 52092 25112
rect 52144 25100 52150 25152
rect 52181 25143 52239 25149
rect 52181 25109 52193 25143
rect 52227 25140 52239 25143
rect 52730 25140 52736 25152
rect 52227 25112 52736 25140
rect 52227 25109 52239 25112
rect 52181 25103 52239 25109
rect 52730 25100 52736 25112
rect 52788 25100 52794 25152
rect 53576 25140 53604 25180
rect 53650 25168 53656 25220
rect 53708 25208 53714 25220
rect 56980 25208 57008 25239
rect 53708 25180 57008 25208
rect 53708 25168 53714 25180
rect 57698 25140 57704 25152
rect 53576 25112 57704 25140
rect 57698 25100 57704 25112
rect 57756 25100 57762 25152
rect 1104 25050 58880 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 58880 25050
rect 1104 24976 58880 24998
rect 50798 24896 50804 24948
rect 50856 24936 50862 24948
rect 53650 24936 53656 24948
rect 50856 24908 53656 24936
rect 50856 24896 50862 24908
rect 53650 24896 53656 24908
rect 53708 24896 53714 24948
rect 55214 24936 55220 24948
rect 53760 24908 55220 24936
rect 2774 24800 2780 24812
rect 2735 24772 2780 24800
rect 2774 24760 2780 24772
rect 2832 24760 2838 24812
rect 49528 24772 51856 24800
rect 3142 24692 3148 24744
rect 3200 24732 3206 24744
rect 49528 24741 49556 24772
rect 3421 24735 3479 24741
rect 3421 24732 3433 24735
rect 3200 24704 3433 24732
rect 3200 24692 3206 24704
rect 3421 24701 3433 24704
rect 3467 24701 3479 24735
rect 3421 24695 3479 24701
rect 49513 24735 49571 24741
rect 49513 24701 49525 24735
rect 49559 24701 49571 24735
rect 50154 24732 50160 24744
rect 50115 24704 50160 24732
rect 49513 24695 49571 24701
rect 50154 24692 50160 24704
rect 50212 24692 50218 24744
rect 50614 24692 50620 24744
rect 50672 24732 50678 24744
rect 51721 24735 51779 24741
rect 51721 24732 51733 24735
rect 50672 24704 51733 24732
rect 50672 24692 50678 24704
rect 51721 24701 51733 24704
rect 51767 24701 51779 24735
rect 51828 24732 51856 24772
rect 53760 24732 53788 24908
rect 55214 24896 55220 24908
rect 55272 24896 55278 24948
rect 53944 24840 54248 24868
rect 53834 24760 53840 24812
rect 53892 24800 53898 24812
rect 53944 24800 53972 24840
rect 54110 24800 54116 24812
rect 53892 24772 53972 24800
rect 54071 24772 54116 24800
rect 53892 24760 53898 24772
rect 54110 24760 54116 24772
rect 54168 24760 54174 24812
rect 51828 24704 53788 24732
rect 51721 24695 51779 24701
rect 53926 24692 53932 24744
rect 53984 24732 53990 24744
rect 54220 24741 54248 24840
rect 54754 24760 54760 24812
rect 54812 24800 54818 24812
rect 54941 24803 54999 24809
rect 54941 24800 54953 24803
rect 54812 24772 54953 24800
rect 54812 24760 54818 24772
rect 54941 24769 54953 24772
rect 54987 24769 54999 24803
rect 54941 24763 54999 24769
rect 54021 24735 54079 24741
rect 54021 24732 54033 24735
rect 53984 24704 54033 24732
rect 53984 24692 53990 24704
rect 54021 24701 54033 24704
rect 54067 24701 54079 24735
rect 54021 24695 54079 24701
rect 54205 24735 54263 24741
rect 54205 24701 54217 24735
rect 54251 24701 54263 24735
rect 54205 24695 54263 24701
rect 57241 24735 57299 24741
rect 57241 24701 57253 24735
rect 57287 24732 57299 24735
rect 57330 24732 57336 24744
rect 57287 24704 57336 24732
rect 57287 24701 57299 24704
rect 57241 24695 57299 24701
rect 57330 24692 57336 24704
rect 57388 24732 57394 24744
rect 58342 24732 58348 24744
rect 57388 24704 58348 24732
rect 57388 24692 57394 24704
rect 58342 24692 58348 24704
rect 58400 24692 58406 24744
rect 1857 24667 1915 24673
rect 1857 24633 1869 24667
rect 1903 24664 1915 24667
rect 2038 24664 2044 24676
rect 1903 24636 2044 24664
rect 1903 24633 1915 24636
rect 1857 24627 1915 24633
rect 2038 24624 2044 24636
rect 2096 24624 2102 24676
rect 2590 24664 2596 24676
rect 2551 24636 2596 24664
rect 2590 24624 2596 24636
rect 2648 24624 2654 24676
rect 50062 24624 50068 24676
rect 50120 24664 50126 24676
rect 50893 24667 50951 24673
rect 50893 24664 50905 24667
rect 50120 24636 50905 24664
rect 50120 24624 50126 24636
rect 50893 24633 50905 24636
rect 50939 24664 50951 24667
rect 50982 24664 50988 24676
rect 50939 24636 50988 24664
rect 50939 24633 50951 24636
rect 50893 24627 50951 24633
rect 50982 24624 50988 24636
rect 51040 24624 51046 24676
rect 51074 24624 51080 24676
rect 51132 24664 51138 24676
rect 51988 24667 52046 24673
rect 51132 24636 51225 24664
rect 51132 24624 51138 24636
rect 51988 24633 52000 24667
rect 52034 24664 52046 24667
rect 52362 24664 52368 24676
rect 52034 24636 52368 24664
rect 52034 24633 52046 24636
rect 51988 24627 52046 24633
rect 52362 24624 52368 24636
rect 52420 24624 52426 24676
rect 54846 24664 54852 24676
rect 52472 24636 54852 24664
rect 1946 24596 1952 24608
rect 1907 24568 1952 24596
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 3234 24596 3240 24608
rect 3195 24568 3240 24596
rect 3234 24556 3240 24568
rect 3292 24556 3298 24608
rect 49970 24556 49976 24608
rect 50028 24596 50034 24608
rect 50341 24599 50399 24605
rect 50341 24596 50353 24599
rect 50028 24568 50353 24596
rect 50028 24556 50034 24568
rect 50341 24565 50353 24568
rect 50387 24565 50399 24599
rect 51092 24596 51120 24624
rect 52472 24596 52500 24636
rect 54846 24624 54852 24636
rect 54904 24624 54910 24676
rect 55030 24624 55036 24676
rect 55088 24664 55094 24676
rect 55186 24667 55244 24673
rect 55186 24664 55198 24667
rect 55088 24636 55198 24664
rect 55088 24624 55094 24636
rect 55186 24633 55198 24636
rect 55232 24633 55244 24667
rect 55186 24627 55244 24633
rect 56226 24624 56232 24676
rect 56284 24664 56290 24676
rect 57974 24664 57980 24676
rect 56284 24636 57468 24664
rect 57935 24636 57980 24664
rect 56284 24624 56290 24636
rect 51092 24568 52500 24596
rect 53101 24599 53159 24605
rect 50341 24559 50399 24565
rect 53101 24565 53113 24599
rect 53147 24596 53159 24599
rect 53742 24596 53748 24608
rect 53147 24568 53748 24596
rect 53147 24565 53159 24568
rect 53101 24559 53159 24565
rect 53742 24556 53748 24568
rect 53800 24556 53806 24608
rect 54202 24556 54208 24608
rect 54260 24596 54266 24608
rect 55950 24596 55956 24608
rect 54260 24568 55956 24596
rect 54260 24556 54266 24568
rect 55950 24556 55956 24568
rect 56008 24596 56014 24608
rect 57440 24605 57468 24636
rect 57974 24624 57980 24636
rect 58032 24624 58038 24676
rect 58158 24664 58164 24676
rect 58119 24636 58164 24664
rect 58158 24624 58164 24636
rect 58216 24624 58222 24676
rect 56321 24599 56379 24605
rect 56321 24596 56333 24599
rect 56008 24568 56333 24596
rect 56008 24556 56014 24568
rect 56321 24565 56333 24568
rect 56367 24565 56379 24599
rect 56321 24559 56379 24565
rect 57425 24599 57483 24605
rect 57425 24565 57437 24599
rect 57471 24565 57483 24599
rect 57425 24559 57483 24565
rect 1104 24506 58880 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 50326 24506
rect 50378 24454 50390 24506
rect 50442 24454 50454 24506
rect 50506 24454 50518 24506
rect 50570 24454 58880 24506
rect 1104 24432 58880 24454
rect 2317 24395 2375 24401
rect 2317 24361 2329 24395
rect 2363 24392 2375 24395
rect 2590 24392 2596 24404
rect 2363 24364 2596 24392
rect 2363 24361 2375 24364
rect 2317 24355 2375 24361
rect 2590 24352 2596 24364
rect 2648 24352 2654 24404
rect 51902 24392 51908 24404
rect 51863 24364 51908 24392
rect 51902 24352 51908 24364
rect 51960 24352 51966 24404
rect 54389 24395 54447 24401
rect 54389 24392 54401 24395
rect 53116 24364 54401 24392
rect 53006 24324 53012 24336
rect 52748 24296 53012 24324
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24256 1731 24259
rect 2961 24259 3019 24265
rect 2961 24256 2973 24259
rect 1719 24228 2973 24256
rect 1719 24225 1731 24228
rect 1673 24219 1731 24225
rect 2961 24225 2973 24228
rect 3007 24225 3019 24259
rect 52086 24256 52092 24268
rect 52047 24228 52092 24256
rect 2961 24219 3019 24225
rect 52086 24216 52092 24228
rect 52144 24216 52150 24268
rect 52748 24265 52776 24296
rect 53006 24284 53012 24296
rect 53064 24284 53070 24336
rect 52733 24259 52791 24265
rect 52733 24225 52745 24259
rect 52779 24225 52791 24259
rect 52733 24219 52791 24225
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24188 1915 24191
rect 3234 24188 3240 24200
rect 1903 24160 3240 24188
rect 1903 24157 1915 24160
rect 1857 24151 1915 24157
rect 3234 24148 3240 24160
rect 3292 24148 3298 24200
rect 52549 24191 52607 24197
rect 52549 24157 52561 24191
rect 52595 24188 52607 24191
rect 52822 24188 52828 24200
rect 52595 24160 52828 24188
rect 52595 24157 52607 24160
rect 52549 24151 52607 24157
rect 52822 24148 52828 24160
rect 52880 24188 52886 24200
rect 53116 24197 53144 24364
rect 54389 24361 54401 24364
rect 54435 24361 54447 24395
rect 54389 24355 54447 24361
rect 54570 24352 54576 24404
rect 54628 24392 54634 24404
rect 54628 24364 55260 24392
rect 54628 24352 54634 24364
rect 53653 24327 53711 24333
rect 53653 24293 53665 24327
rect 53699 24324 53711 24327
rect 54662 24324 54668 24336
rect 53699 24296 54668 24324
rect 53699 24293 53711 24296
rect 53653 24287 53711 24293
rect 54662 24284 54668 24296
rect 54720 24324 54726 24336
rect 54720 24296 54800 24324
rect 54720 24284 54726 24296
rect 53561 24259 53619 24265
rect 53561 24225 53573 24259
rect 53607 24225 53619 24259
rect 53742 24256 53748 24268
rect 53703 24228 53748 24256
rect 53561 24219 53619 24225
rect 53101 24191 53159 24197
rect 53101 24188 53113 24191
rect 52880 24160 53113 24188
rect 52880 24148 52886 24160
rect 53101 24157 53113 24160
rect 53147 24157 53159 24191
rect 53576 24188 53604 24219
rect 53742 24216 53748 24228
rect 53800 24256 53806 24268
rect 54389 24259 54447 24265
rect 54389 24256 54401 24259
rect 53800 24228 54401 24256
rect 53800 24216 53806 24228
rect 54389 24225 54401 24228
rect 54435 24256 54447 24259
rect 54570 24256 54576 24268
rect 54435 24228 54576 24256
rect 54435 24225 54447 24228
rect 54389 24219 54447 24225
rect 54570 24216 54576 24228
rect 54628 24216 54634 24268
rect 54772 24265 54800 24296
rect 55232 24265 55260 24364
rect 57974 24352 57980 24404
rect 58032 24392 58038 24404
rect 58161 24395 58219 24401
rect 58161 24392 58173 24395
rect 58032 24364 58173 24392
rect 58032 24352 58038 24364
rect 58161 24361 58173 24364
rect 58207 24361 58219 24395
rect 58161 24355 58219 24361
rect 54757 24259 54815 24265
rect 54757 24225 54769 24259
rect 54803 24225 54815 24259
rect 54757 24219 54815 24225
rect 55217 24259 55275 24265
rect 55217 24225 55229 24259
rect 55263 24225 55275 24259
rect 56870 24256 56876 24268
rect 56831 24228 56876 24256
rect 55217 24219 55275 24225
rect 56870 24216 56876 24228
rect 56928 24216 56934 24268
rect 54202 24188 54208 24200
rect 53576 24160 54208 24188
rect 53101 24151 53159 24157
rect 54202 24148 54208 24160
rect 54260 24148 54266 24200
rect 57517 24191 57575 24197
rect 57517 24157 57529 24191
rect 57563 24157 57575 24191
rect 57698 24188 57704 24200
rect 57659 24160 57704 24188
rect 57517 24151 57575 24157
rect 50525 24123 50583 24129
rect 50525 24089 50537 24123
rect 50571 24120 50583 24123
rect 57532 24120 57560 24151
rect 57698 24148 57704 24160
rect 57756 24148 57762 24200
rect 50571 24092 54340 24120
rect 50571 24089 50583 24092
rect 50525 24083 50583 24089
rect 52454 24012 52460 24064
rect 52512 24052 52518 24064
rect 52825 24055 52883 24061
rect 52825 24052 52837 24055
rect 52512 24024 52837 24052
rect 52512 24012 52518 24024
rect 52825 24021 52837 24024
rect 52871 24021 52883 24055
rect 54312 24052 54340 24092
rect 54772 24092 57560 24120
rect 54772 24052 54800 24092
rect 54312 24024 54800 24052
rect 52825 24015 52883 24021
rect 55122 24012 55128 24064
rect 55180 24052 55186 24064
rect 55309 24055 55367 24061
rect 55309 24052 55321 24055
rect 55180 24024 55321 24052
rect 55180 24012 55186 24024
rect 55309 24021 55321 24024
rect 55355 24021 55367 24055
rect 56962 24052 56968 24064
rect 56923 24024 56968 24052
rect 55309 24015 55367 24021
rect 56962 24012 56968 24024
rect 57020 24012 57026 24064
rect 1104 23962 58880 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 58880 23962
rect 1104 23888 58880 23910
rect 2038 23848 2044 23860
rect 1999 23820 2044 23848
rect 2038 23808 2044 23820
rect 2096 23808 2102 23860
rect 50525 23851 50583 23857
rect 50525 23817 50537 23851
rect 50571 23848 50583 23851
rect 50798 23848 50804 23860
rect 50571 23820 50804 23848
rect 50571 23817 50583 23820
rect 50525 23811 50583 23817
rect 50798 23808 50804 23820
rect 50856 23808 50862 23860
rect 52362 23808 52368 23860
rect 52420 23848 52426 23860
rect 52457 23851 52515 23857
rect 52457 23848 52469 23851
rect 52420 23820 52469 23848
rect 52420 23808 52426 23820
rect 52457 23817 52469 23820
rect 52503 23817 52515 23851
rect 52457 23811 52515 23817
rect 53006 23808 53012 23860
rect 53064 23848 53070 23860
rect 54021 23851 54079 23857
rect 54021 23848 54033 23851
rect 53064 23820 54033 23848
rect 53064 23808 53070 23820
rect 54021 23817 54033 23820
rect 54067 23817 54079 23851
rect 54021 23811 54079 23817
rect 54941 23851 54999 23857
rect 54941 23817 54953 23851
rect 54987 23848 54999 23851
rect 55030 23848 55036 23860
rect 54987 23820 55036 23848
rect 54987 23817 54999 23820
rect 54941 23811 54999 23817
rect 55030 23808 55036 23820
rect 55088 23808 55094 23860
rect 51813 23783 51871 23789
rect 51813 23749 51825 23783
rect 51859 23780 51871 23783
rect 57698 23780 57704 23792
rect 51859 23752 57704 23780
rect 51859 23749 51871 23752
rect 51813 23743 51871 23749
rect 57698 23740 57704 23752
rect 57756 23740 57762 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 2961 23715 3019 23721
rect 2961 23712 2973 23715
rect 1719 23684 2973 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2961 23681 2973 23684
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 50154 23672 50160 23724
rect 50212 23712 50218 23724
rect 50798 23712 50804 23724
rect 50212 23684 50804 23712
rect 50212 23672 50218 23684
rect 50798 23672 50804 23684
rect 50856 23712 50862 23724
rect 52086 23712 52092 23724
rect 50856 23684 51074 23712
rect 51999 23684 52092 23712
rect 50856 23672 50862 23684
rect 1854 23644 1860 23656
rect 1815 23616 1860 23644
rect 1854 23604 1860 23616
rect 1912 23604 1918 23656
rect 49237 23647 49295 23653
rect 49237 23613 49249 23647
rect 49283 23613 49295 23647
rect 49237 23607 49295 23613
rect 50065 23647 50123 23653
rect 50065 23613 50077 23647
rect 50111 23644 50123 23647
rect 50706 23644 50712 23656
rect 50111 23616 50712 23644
rect 50111 23613 50123 23616
rect 50065 23607 50123 23613
rect 49252 23576 49280 23607
rect 50706 23604 50712 23616
rect 50764 23604 50770 23656
rect 51046 23644 51074 23684
rect 52012 23653 52040 23684
rect 52086 23672 52092 23684
rect 52144 23712 52150 23724
rect 56226 23712 56232 23724
rect 52144 23684 56232 23712
rect 52144 23672 52150 23684
rect 56226 23672 56232 23684
rect 56284 23672 56290 23724
rect 51169 23647 51227 23653
rect 51169 23644 51181 23647
rect 51046 23616 51181 23644
rect 51169 23613 51181 23616
rect 51215 23613 51227 23647
rect 51169 23607 51227 23613
rect 51997 23647 52055 23653
rect 51997 23613 52009 23647
rect 52043 23613 52055 23647
rect 52454 23644 52460 23656
rect 52415 23616 52460 23644
rect 51997 23607 52055 23613
rect 52454 23604 52460 23616
rect 52512 23604 52518 23656
rect 52546 23604 52552 23656
rect 52604 23644 52610 23656
rect 52641 23647 52699 23653
rect 52641 23644 52653 23647
rect 52604 23616 52653 23644
rect 52604 23604 52610 23616
rect 52641 23613 52653 23616
rect 52687 23613 52699 23647
rect 52641 23607 52699 23613
rect 52730 23604 52736 23656
rect 52788 23644 52794 23656
rect 54205 23647 54263 23653
rect 54205 23644 54217 23647
rect 52788 23616 54217 23644
rect 52788 23604 52794 23616
rect 54205 23613 54217 23616
rect 54251 23613 54263 23647
rect 54386 23644 54392 23656
rect 54347 23616 54392 23644
rect 54205 23607 54263 23613
rect 54386 23604 54392 23616
rect 54444 23604 54450 23656
rect 54478 23604 54484 23656
rect 54536 23644 54542 23656
rect 54938 23644 54944 23656
rect 54536 23616 54581 23644
rect 54899 23616 54944 23644
rect 54536 23604 54542 23616
rect 54938 23604 54944 23616
rect 54996 23604 55002 23656
rect 55122 23644 55128 23656
rect 55083 23616 55128 23644
rect 55122 23604 55128 23616
rect 55180 23604 55186 23656
rect 55950 23644 55956 23656
rect 55911 23616 55956 23644
rect 55950 23604 55956 23616
rect 56008 23604 56014 23656
rect 55214 23576 55220 23588
rect 49252 23548 55220 23576
rect 55214 23536 55220 23548
rect 55272 23536 55278 23588
rect 57238 23576 57244 23588
rect 57199 23548 57244 23576
rect 57238 23536 57244 23548
rect 57296 23536 57302 23588
rect 57422 23576 57428 23588
rect 57383 23548 57428 23576
rect 57422 23536 57428 23548
rect 57480 23536 57486 23588
rect 57974 23576 57980 23588
rect 57935 23548 57980 23576
rect 57974 23536 57980 23548
rect 58032 23536 58038 23588
rect 49878 23508 49884 23520
rect 49839 23480 49884 23508
rect 49878 23468 49884 23480
rect 49936 23468 49942 23520
rect 50706 23468 50712 23520
rect 50764 23508 50770 23520
rect 51353 23511 51411 23517
rect 51353 23508 51365 23511
rect 50764 23480 51365 23508
rect 50764 23468 50770 23480
rect 51353 23477 51365 23480
rect 51399 23477 51411 23511
rect 51353 23471 51411 23477
rect 52546 23468 52552 23520
rect 52604 23508 52610 23520
rect 53650 23508 53656 23520
rect 52604 23480 53656 23508
rect 52604 23468 52610 23480
rect 53650 23468 53656 23480
rect 53708 23468 53714 23520
rect 56042 23508 56048 23520
rect 56003 23480 56048 23508
rect 56042 23468 56048 23480
rect 56100 23468 56106 23520
rect 57882 23468 57888 23520
rect 57940 23508 57946 23520
rect 58069 23511 58127 23517
rect 58069 23508 58081 23511
rect 57940 23480 58081 23508
rect 57940 23468 57946 23480
rect 58069 23477 58081 23480
rect 58115 23477 58127 23511
rect 58069 23471 58127 23477
rect 1104 23418 58880 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 50326 23418
rect 50378 23366 50390 23418
rect 50442 23366 50454 23418
rect 50506 23366 50518 23418
rect 50570 23366 58880 23418
rect 1104 23344 58880 23366
rect 1854 23264 1860 23316
rect 1912 23304 1918 23316
rect 2501 23307 2559 23313
rect 2501 23304 2513 23307
rect 1912 23276 2513 23304
rect 1912 23264 1918 23276
rect 2501 23273 2513 23276
rect 2547 23273 2559 23307
rect 2501 23267 2559 23273
rect 49878 23264 49884 23316
rect 49936 23304 49942 23316
rect 49936 23276 57376 23304
rect 49936 23264 49942 23276
rect 50430 23236 50436 23248
rect 50391 23208 50436 23236
rect 50430 23196 50436 23208
rect 50488 23196 50494 23248
rect 56042 23236 56048 23248
rect 51046 23208 56048 23236
rect 1854 23168 1860 23180
rect 1815 23140 1860 23168
rect 1854 23128 1860 23140
rect 1912 23128 1918 23180
rect 2685 23171 2743 23177
rect 2685 23137 2697 23171
rect 2731 23168 2743 23171
rect 3142 23168 3148 23180
rect 2731 23140 3148 23168
rect 2731 23137 2743 23140
rect 2685 23131 2743 23137
rect 3142 23128 3148 23140
rect 3200 23128 3206 23180
rect 49878 23128 49884 23180
rect 49936 23168 49942 23180
rect 50341 23171 50399 23177
rect 50341 23168 50353 23171
rect 49936 23140 50353 23168
rect 49936 23128 49942 23140
rect 50341 23137 50353 23140
rect 50387 23137 50399 23171
rect 50341 23131 50399 23137
rect 50525 23171 50583 23177
rect 50525 23137 50537 23171
rect 50571 23168 50583 23171
rect 51046 23168 51074 23208
rect 50571 23140 51074 23168
rect 51445 23171 51503 23177
rect 50571 23137 50583 23140
rect 50525 23131 50583 23137
rect 51445 23137 51457 23171
rect 51491 23168 51503 23171
rect 51721 23171 51779 23177
rect 51721 23168 51733 23171
rect 51491 23140 51733 23168
rect 51491 23137 51503 23140
rect 51445 23131 51503 23137
rect 51721 23137 51733 23140
rect 51767 23137 51779 23171
rect 51721 23131 51779 23137
rect 52086 23128 52092 23180
rect 52144 23168 52150 23180
rect 52437 23171 52495 23177
rect 52437 23168 52449 23171
rect 52144 23140 52449 23168
rect 52144 23128 52150 23140
rect 52437 23137 52449 23140
rect 52483 23137 52495 23171
rect 52437 23131 52495 23137
rect 54202 23128 54208 23180
rect 54260 23168 54266 23180
rect 54478 23168 54484 23180
rect 54260 23140 54484 23168
rect 54260 23128 54266 23140
rect 54478 23128 54484 23140
rect 54536 23128 54542 23180
rect 54772 23177 54800 23208
rect 56042 23196 56048 23208
rect 56100 23196 56106 23248
rect 54757 23171 54815 23177
rect 54757 23137 54769 23171
rect 54803 23137 54815 23171
rect 54757 23131 54815 23137
rect 54941 23171 54999 23177
rect 54941 23137 54953 23171
rect 54987 23168 54999 23171
rect 55122 23168 55128 23180
rect 54987 23140 55128 23168
rect 54987 23137 54999 23140
rect 54941 23131 54999 23137
rect 55122 23128 55128 23140
rect 55180 23128 55186 23180
rect 55582 23168 55588 23180
rect 55543 23140 55588 23168
rect 55582 23128 55588 23140
rect 55640 23128 55646 23180
rect 57146 23168 57152 23180
rect 57107 23140 57152 23168
rect 57146 23128 57152 23140
rect 57204 23128 57210 23180
rect 57348 23177 57376 23276
rect 57333 23171 57391 23177
rect 57333 23137 57345 23171
rect 57379 23137 57391 23171
rect 57333 23131 57391 23137
rect 49970 23060 49976 23112
rect 50028 23100 50034 23112
rect 52181 23103 52239 23109
rect 52181 23100 52193 23103
rect 50028 23072 52193 23100
rect 50028 23060 50034 23072
rect 52181 23069 52193 23072
rect 52227 23069 52239 23103
rect 54662 23100 54668 23112
rect 54623 23072 54668 23100
rect 52181 23063 52239 23069
rect 54662 23060 54668 23072
rect 54720 23060 54726 23112
rect 1578 22992 1584 23044
rect 1636 23032 1642 23044
rect 3329 23035 3387 23041
rect 3329 23032 3341 23035
rect 1636 23004 3341 23032
rect 1636 22992 1642 23004
rect 3329 23001 3341 23004
rect 3375 23001 3387 23035
rect 3329 22995 3387 23001
rect 53834 22992 53840 23044
rect 53892 23032 53898 23044
rect 54297 23035 54355 23041
rect 54297 23032 54309 23035
rect 53892 23004 54309 23032
rect 53892 22992 53898 23004
rect 54297 23001 54309 23004
rect 54343 23001 54355 23035
rect 54297 22995 54355 23001
rect 54386 22992 54392 23044
rect 54444 23032 54450 23044
rect 54573 23035 54631 23041
rect 54573 23032 54585 23035
rect 54444 23004 54585 23032
rect 54444 22992 54450 23004
rect 54573 23001 54585 23004
rect 54619 23032 54631 23035
rect 55677 23035 55735 23041
rect 55677 23032 55689 23035
rect 54619 23004 55689 23032
rect 54619 23001 54631 23004
rect 54573 22995 54631 23001
rect 55677 23001 55689 23004
rect 55723 23001 55735 23035
rect 55677 22995 55735 23001
rect 56870 22992 56876 23044
rect 56928 23032 56934 23044
rect 57517 23035 57575 23041
rect 57517 23032 57529 23035
rect 56928 23004 57529 23032
rect 56928 22992 56934 23004
rect 57517 23001 57529 23004
rect 57563 23001 57575 23035
rect 57517 22995 57575 23001
rect 1946 22964 1952 22976
rect 1907 22936 1952 22964
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 49786 22924 49792 22976
rect 49844 22964 49850 22976
rect 51445 22967 51503 22973
rect 51445 22964 51457 22967
rect 49844 22936 51457 22964
rect 49844 22924 49850 22936
rect 51445 22933 51457 22936
rect 51491 22933 51503 22967
rect 51445 22927 51503 22933
rect 51537 22967 51595 22973
rect 51537 22933 51549 22967
rect 51583 22964 51595 22967
rect 51994 22964 52000 22976
rect 51583 22936 52000 22964
rect 51583 22933 51595 22936
rect 51537 22927 51595 22933
rect 51994 22924 52000 22936
rect 52052 22924 52058 22976
rect 53561 22967 53619 22973
rect 53561 22933 53573 22967
rect 53607 22964 53619 22967
rect 54110 22964 54116 22976
rect 53607 22936 54116 22964
rect 53607 22933 53619 22936
rect 53561 22927 53619 22933
rect 54110 22924 54116 22936
rect 54168 22924 54174 22976
rect 1104 22874 58880 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 58880 22874
rect 1104 22800 58880 22822
rect 1854 22720 1860 22772
rect 1912 22760 1918 22772
rect 1949 22763 2007 22769
rect 1949 22760 1961 22763
rect 1912 22732 1961 22760
rect 1912 22720 1918 22732
rect 1949 22729 1961 22732
rect 1995 22729 2007 22763
rect 1949 22723 2007 22729
rect 2869 22763 2927 22769
rect 2869 22729 2881 22763
rect 2915 22760 2927 22763
rect 3142 22760 3148 22772
rect 2915 22732 3148 22760
rect 2915 22729 2927 22732
rect 2869 22723 2927 22729
rect 3142 22720 3148 22732
rect 3200 22720 3206 22772
rect 51537 22763 51595 22769
rect 51537 22729 51549 22763
rect 51583 22760 51595 22763
rect 51718 22760 51724 22772
rect 51583 22732 51724 22760
rect 51583 22729 51595 22732
rect 51537 22723 51595 22729
rect 51718 22720 51724 22732
rect 51776 22720 51782 22772
rect 52086 22760 52092 22772
rect 52047 22732 52092 22760
rect 52086 22720 52092 22732
rect 52144 22720 52150 22772
rect 53742 22720 53748 22772
rect 53800 22760 53806 22772
rect 53800 22732 54064 22760
rect 53800 22720 53806 22732
rect 3329 22695 3387 22701
rect 3329 22692 3341 22695
rect 1780 22664 3341 22692
rect 1578 22624 1584 22636
rect 1539 22596 1584 22624
rect 1578 22584 1584 22596
rect 1636 22584 1642 22636
rect 1780 22633 1808 22664
rect 3329 22661 3341 22664
rect 3375 22661 3387 22695
rect 3329 22655 3387 22661
rect 50801 22695 50859 22701
rect 50801 22661 50813 22695
rect 50847 22692 50859 22695
rect 50847 22664 53880 22692
rect 50847 22661 50859 22664
rect 50801 22655 50859 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 50249 22627 50307 22633
rect 50249 22593 50261 22627
rect 50295 22624 50307 22627
rect 53742 22624 53748 22636
rect 50295 22596 53748 22624
rect 50295 22593 50307 22596
rect 50249 22587 50307 22593
rect 53742 22584 53748 22596
rect 53800 22584 53806 22636
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22556 2743 22559
rect 2958 22556 2964 22568
rect 2731 22528 2964 22556
rect 2731 22525 2743 22528
rect 2685 22519 2743 22525
rect 2958 22516 2964 22528
rect 3016 22516 3022 22568
rect 3142 22516 3148 22568
rect 3200 22556 3206 22568
rect 3513 22559 3571 22565
rect 3513 22556 3525 22559
rect 3200 22528 3525 22556
rect 3200 22516 3206 22528
rect 3513 22525 3525 22528
rect 3559 22525 3571 22559
rect 3513 22519 3571 22525
rect 49878 22516 49884 22568
rect 49936 22556 49942 22568
rect 50157 22559 50215 22565
rect 50157 22556 50169 22559
rect 49936 22528 50169 22556
rect 49936 22516 49942 22528
rect 50157 22525 50169 22528
rect 50203 22525 50215 22559
rect 50157 22519 50215 22525
rect 50341 22559 50399 22565
rect 50341 22525 50353 22559
rect 50387 22556 50399 22559
rect 50614 22556 50620 22568
rect 50387 22528 50620 22556
rect 50387 22525 50399 22528
rect 50341 22519 50399 22525
rect 50614 22516 50620 22528
rect 50672 22516 50678 22568
rect 50706 22516 50712 22568
rect 50764 22556 50770 22568
rect 50985 22559 51043 22565
rect 50985 22556 50997 22559
rect 50764 22528 50997 22556
rect 50764 22516 50770 22528
rect 50985 22525 50997 22528
rect 51031 22525 51043 22559
rect 50985 22519 51043 22525
rect 51445 22559 51503 22565
rect 51445 22525 51457 22559
rect 51491 22525 51503 22559
rect 51445 22519 51503 22525
rect 51629 22559 51687 22565
rect 51629 22525 51641 22559
rect 51675 22556 51687 22559
rect 52362 22556 52368 22568
rect 51675 22528 52368 22556
rect 51675 22525 51687 22528
rect 51629 22519 51687 22525
rect 51460 22488 51488 22519
rect 52362 22516 52368 22528
rect 52420 22516 52426 22568
rect 52454 22559 52512 22565
rect 52454 22525 52466 22559
rect 52500 22525 52512 22559
rect 52454 22519 52512 22525
rect 52549 22559 52607 22565
rect 52549 22525 52561 22559
rect 52595 22525 52607 22559
rect 52730 22556 52736 22568
rect 52691 22528 52736 22556
rect 52549 22519 52607 22525
rect 52270 22488 52276 22500
rect 51460 22460 52276 22488
rect 52270 22448 52276 22460
rect 52328 22488 52334 22500
rect 52469 22488 52497 22519
rect 52328 22460 52497 22488
rect 52564 22488 52592 22519
rect 52730 22516 52736 22528
rect 52788 22516 52794 22568
rect 52638 22488 52644 22500
rect 52564 22460 52644 22488
rect 52328 22448 52334 22460
rect 52638 22448 52644 22460
rect 52696 22448 52702 22500
rect 53852 22488 53880 22664
rect 54036 22624 54064 22732
rect 55582 22720 55588 22772
rect 55640 22760 55646 22772
rect 56226 22760 56232 22772
rect 55640 22732 56232 22760
rect 55640 22720 55646 22732
rect 56226 22720 56232 22732
rect 56284 22720 56290 22772
rect 57238 22720 57244 22772
rect 57296 22760 57302 22772
rect 57333 22763 57391 22769
rect 57333 22760 57345 22763
rect 57296 22732 57345 22760
rect 57296 22720 57302 22732
rect 57333 22729 57345 22732
rect 57379 22729 57391 22763
rect 57333 22723 57391 22729
rect 54036 22596 54984 22624
rect 54110 22556 54116 22568
rect 54071 22528 54116 22556
rect 54110 22516 54116 22528
rect 54168 22516 54174 22568
rect 54846 22556 54852 22568
rect 54807 22528 54852 22556
rect 54846 22516 54852 22528
rect 54904 22516 54910 22568
rect 54956 22556 54984 22596
rect 56965 22559 57023 22565
rect 56965 22556 56977 22559
rect 54956 22528 56977 22556
rect 56965 22525 56977 22528
rect 57011 22525 57023 22559
rect 56965 22519 57023 22525
rect 57149 22559 57207 22565
rect 57149 22525 57161 22559
rect 57195 22525 57207 22559
rect 57149 22519 57207 22525
rect 53852 22460 54892 22488
rect 51994 22380 52000 22432
rect 52052 22420 52058 22432
rect 53374 22420 53380 22432
rect 52052 22392 53380 22420
rect 52052 22380 52058 22392
rect 53374 22380 53380 22392
rect 53432 22380 53438 22432
rect 54202 22420 54208 22432
rect 54163 22392 54208 22420
rect 54202 22380 54208 22392
rect 54260 22380 54266 22432
rect 54864 22420 54892 22460
rect 54938 22448 54944 22500
rect 54996 22488 55002 22500
rect 55094 22491 55152 22497
rect 55094 22488 55106 22491
rect 54996 22460 55106 22488
rect 54996 22448 55002 22460
rect 55094 22457 55106 22460
rect 55140 22457 55152 22491
rect 55094 22451 55152 22457
rect 57164 22420 57192 22519
rect 54864 22392 57192 22420
rect 1104 22330 58880 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 50326 22330
rect 50378 22278 50390 22330
rect 50442 22278 50454 22330
rect 50506 22278 50518 22330
rect 50570 22278 58880 22330
rect 1104 22256 58880 22278
rect 50614 22176 50620 22228
rect 50672 22216 50678 22228
rect 54294 22216 54300 22228
rect 50672 22188 54300 22216
rect 50672 22176 50678 22188
rect 54294 22176 54300 22188
rect 54352 22176 54358 22228
rect 54938 22216 54944 22228
rect 54899 22188 54944 22216
rect 54938 22176 54944 22188
rect 54996 22176 55002 22228
rect 2593 22151 2651 22157
rect 2593 22117 2605 22151
rect 2639 22148 2651 22151
rect 2958 22148 2964 22160
rect 2639 22120 2964 22148
rect 2639 22117 2651 22120
rect 2593 22111 2651 22117
rect 2958 22108 2964 22120
rect 3016 22108 3022 22160
rect 51350 22108 51356 22160
rect 51408 22148 51414 22160
rect 51537 22151 51595 22157
rect 51537 22148 51549 22151
rect 51408 22120 51549 22148
rect 51408 22108 51414 22120
rect 51537 22117 51549 22120
rect 51583 22117 51595 22151
rect 51537 22111 51595 22117
rect 52362 22108 52368 22160
rect 52420 22148 52426 22160
rect 52420 22120 52960 22148
rect 52420 22108 52426 22120
rect 1854 22080 1860 22092
rect 1815 22052 1860 22080
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 49237 22083 49295 22089
rect 49237 22049 49249 22083
rect 49283 22080 49295 22083
rect 49326 22080 49332 22092
rect 49283 22052 49332 22080
rect 49283 22049 49295 22052
rect 49237 22043 49295 22049
rect 49326 22040 49332 22052
rect 49384 22040 49390 22092
rect 49697 22083 49755 22089
rect 49697 22049 49709 22083
rect 49743 22049 49755 22083
rect 49697 22043 49755 22049
rect 51721 22083 51779 22089
rect 51721 22049 51733 22083
rect 51767 22080 51779 22083
rect 52546 22080 52552 22092
rect 51767 22052 52552 22080
rect 51767 22049 51779 22052
rect 51721 22043 51779 22049
rect 2866 22012 2872 22024
rect 2827 21984 2872 22012
rect 2866 21972 2872 21984
rect 2924 22012 2930 22024
rect 2924 21984 6914 22012
rect 2924 21972 2930 21984
rect 2038 21944 2044 21956
rect 1999 21916 2044 21944
rect 2038 21904 2044 21916
rect 2096 21904 2102 21956
rect 6886 21876 6914 21984
rect 49712 21944 49740 22043
rect 52546 22040 52552 22052
rect 52604 22040 52610 22092
rect 52656 22089 52684 22120
rect 52641 22083 52699 22089
rect 52641 22049 52653 22083
rect 52687 22080 52699 22083
rect 52822 22080 52828 22092
rect 52687 22052 52721 22080
rect 52783 22052 52828 22080
rect 52687 22049 52699 22052
rect 52641 22043 52699 22049
rect 52822 22040 52828 22052
rect 52880 22040 52886 22092
rect 52932 22080 52960 22120
rect 54202 22108 54208 22160
rect 54260 22148 54266 22160
rect 56873 22151 56931 22157
rect 54260 22120 55076 22148
rect 54260 22108 54266 22120
rect 53837 22083 53895 22089
rect 53837 22080 53849 22083
rect 52932 22052 53849 22080
rect 53837 22049 53849 22052
rect 53883 22049 53895 22083
rect 54018 22080 54024 22092
rect 53979 22052 54024 22080
rect 53837 22043 53895 22049
rect 54018 22040 54024 22052
rect 54076 22040 54082 22092
rect 54404 22089 54432 22120
rect 54113 22083 54171 22089
rect 54113 22049 54125 22083
rect 54159 22080 54171 22083
rect 54389 22083 54447 22089
rect 54159 22052 54340 22080
rect 54159 22049 54171 22052
rect 54113 22043 54171 22049
rect 50525 22015 50583 22021
rect 50525 21981 50537 22015
rect 50571 22012 50583 22015
rect 54312 22012 54340 22052
rect 54389 22049 54401 22083
rect 54435 22049 54447 22083
rect 54389 22043 54447 22049
rect 54754 22040 54760 22092
rect 54812 22080 54818 22092
rect 54849 22083 54907 22089
rect 54849 22080 54861 22083
rect 54812 22052 54861 22080
rect 54812 22040 54818 22052
rect 54849 22049 54861 22052
rect 54895 22080 54907 22083
rect 54938 22080 54944 22092
rect 54895 22052 54944 22080
rect 54895 22049 54907 22052
rect 54849 22043 54907 22049
rect 54938 22040 54944 22052
rect 54996 22040 55002 22092
rect 55048 22089 55076 22120
rect 56873 22117 56885 22151
rect 56919 22148 56931 22151
rect 58066 22148 58072 22160
rect 56919 22120 58072 22148
rect 56919 22117 56931 22120
rect 56873 22111 56931 22117
rect 58066 22108 58072 22120
rect 58124 22108 58130 22160
rect 55033 22083 55091 22089
rect 55033 22049 55045 22083
rect 55079 22049 55091 22083
rect 55033 22043 55091 22049
rect 55122 22040 55128 22092
rect 55180 22080 55186 22092
rect 55493 22083 55551 22089
rect 55493 22080 55505 22083
rect 55180 22052 55505 22080
rect 55180 22040 55186 22052
rect 55493 22049 55505 22052
rect 55539 22049 55551 22083
rect 55674 22080 55680 22092
rect 55635 22052 55680 22080
rect 55493 22043 55551 22049
rect 55674 22040 55680 22052
rect 55732 22040 55738 22092
rect 56226 22012 56232 22024
rect 50571 21984 54156 22012
rect 54312 21984 56232 22012
rect 50571 21981 50583 21984
rect 50525 21975 50583 21981
rect 54128 21956 54156 21984
rect 56226 21972 56232 21984
rect 56284 21972 56290 22024
rect 57517 22015 57575 22021
rect 57517 21981 57529 22015
rect 57563 21981 57575 22015
rect 57698 22012 57704 22024
rect 57659 21984 57704 22012
rect 57517 21975 57575 21981
rect 49712 21916 54064 21944
rect 31294 21876 31300 21888
rect 6886 21848 31300 21876
rect 31294 21836 31300 21848
rect 31352 21836 31358 21888
rect 49050 21876 49056 21888
rect 49011 21848 49056 21876
rect 49050 21836 49056 21848
rect 49108 21836 49114 21888
rect 52638 21836 52644 21888
rect 52696 21876 52702 21888
rect 52733 21879 52791 21885
rect 52733 21876 52745 21879
rect 52696 21848 52745 21876
rect 52696 21836 52702 21848
rect 52733 21845 52745 21848
rect 52779 21845 52791 21879
rect 54036 21876 54064 21916
rect 54110 21904 54116 21956
rect 54168 21904 54174 21956
rect 54294 21944 54300 21956
rect 54255 21916 54300 21944
rect 54294 21904 54300 21916
rect 54352 21904 54358 21956
rect 54386 21904 54392 21956
rect 54444 21944 54450 21956
rect 57532 21944 57560 21975
rect 57698 21972 57704 21984
rect 57756 21972 57762 22024
rect 57974 21944 57980 21956
rect 54444 21916 57560 21944
rect 57935 21916 57980 21944
rect 54444 21904 54450 21916
rect 57974 21904 57980 21916
rect 58032 21904 58038 21956
rect 55214 21876 55220 21888
rect 54036 21848 55220 21876
rect 52733 21839 52791 21845
rect 55214 21836 55220 21848
rect 55272 21836 55278 21888
rect 55490 21876 55496 21888
rect 55451 21848 55496 21876
rect 55490 21836 55496 21848
rect 55548 21836 55554 21888
rect 56502 21836 56508 21888
rect 56560 21876 56566 21888
rect 56965 21879 57023 21885
rect 56965 21876 56977 21879
rect 56560 21848 56977 21876
rect 56560 21836 56566 21848
rect 56965 21845 56977 21848
rect 57011 21845 57023 21879
rect 56965 21839 57023 21845
rect 1104 21786 58880 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 58880 21786
rect 1104 21712 58880 21734
rect 1854 21632 1860 21684
rect 1912 21672 1918 21684
rect 2041 21675 2099 21681
rect 2041 21672 2053 21675
rect 1912 21644 2053 21672
rect 1912 21632 1918 21644
rect 2041 21641 2053 21644
rect 2087 21641 2099 21675
rect 4249 21675 4307 21681
rect 4249 21672 4261 21675
rect 2041 21635 2099 21641
rect 2884 21644 4261 21672
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 2884 21536 2912 21644
rect 4249 21641 4261 21644
rect 4295 21641 4307 21675
rect 4249 21635 4307 21641
rect 51810 21632 51816 21684
rect 51868 21672 51874 21684
rect 52457 21675 52515 21681
rect 52457 21672 52469 21675
rect 51868 21644 52469 21672
rect 51868 21632 51874 21644
rect 52457 21641 52469 21644
rect 52503 21641 52515 21675
rect 53190 21672 53196 21684
rect 52457 21635 52515 21641
rect 52840 21644 53196 21672
rect 3142 21604 3148 21616
rect 1719 21508 2912 21536
rect 2976 21576 3148 21604
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 2976 21477 3004 21576
rect 3142 21564 3148 21576
rect 3200 21564 3206 21616
rect 51718 21564 51724 21616
rect 51776 21604 51782 21616
rect 52730 21604 52736 21616
rect 51776 21576 52736 21604
rect 51776 21564 51782 21576
rect 52730 21564 52736 21576
rect 52788 21564 52794 21616
rect 52840 21613 52868 21644
rect 53190 21632 53196 21644
rect 53248 21632 53254 21684
rect 53374 21632 53380 21684
rect 53432 21672 53438 21684
rect 57698 21672 57704 21684
rect 53432 21644 57704 21672
rect 53432 21632 53438 21644
rect 57698 21632 57704 21644
rect 57756 21632 57762 21684
rect 58066 21672 58072 21684
rect 58027 21644 58072 21672
rect 58066 21632 58072 21644
rect 58124 21632 58130 21684
rect 52825 21607 52883 21613
rect 52825 21573 52837 21607
rect 52871 21573 52883 21607
rect 52825 21567 52883 21573
rect 52914 21564 52920 21616
rect 52972 21604 52978 21616
rect 52972 21576 54800 21604
rect 52972 21564 52978 21576
rect 54297 21539 54355 21545
rect 51920 21508 54248 21536
rect 1857 21471 1915 21477
rect 1857 21437 1869 21471
rect 1903 21437 1915 21471
rect 1857 21431 1915 21437
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21437 3019 21471
rect 2961 21431 3019 21437
rect 1872 21400 1900 21431
rect 3050 21428 3056 21480
rect 3108 21468 3114 21480
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 3108 21440 3617 21468
rect 3108 21428 3114 21440
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 49878 21468 49884 21480
rect 49839 21440 49884 21468
rect 3605 21431 3663 21437
rect 49878 21428 49884 21440
rect 49936 21428 49942 21480
rect 50065 21471 50123 21477
rect 50065 21437 50077 21471
rect 50111 21437 50123 21471
rect 50065 21431 50123 21437
rect 3234 21400 3240 21412
rect 1872 21372 3240 21400
rect 3234 21360 3240 21372
rect 3292 21360 3298 21412
rect 2777 21335 2835 21341
rect 2777 21301 2789 21335
rect 2823 21332 2835 21335
rect 2866 21332 2872 21344
rect 2823 21304 2872 21332
rect 2823 21301 2835 21304
rect 2777 21295 2835 21301
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 49970 21332 49976 21344
rect 49931 21304 49976 21332
rect 49970 21292 49976 21304
rect 50028 21292 50034 21344
rect 50080 21332 50108 21431
rect 50154 21428 50160 21480
rect 50212 21468 50218 21480
rect 50525 21471 50583 21477
rect 50525 21468 50537 21471
rect 50212 21440 50537 21468
rect 50212 21428 50218 21440
rect 50525 21437 50537 21440
rect 50571 21437 50583 21471
rect 50525 21431 50583 21437
rect 50614 21360 50620 21412
rect 50672 21400 50678 21412
rect 50770 21403 50828 21409
rect 50770 21400 50782 21403
rect 50672 21372 50782 21400
rect 50672 21360 50678 21372
rect 50770 21369 50782 21372
rect 50816 21369 50828 21403
rect 50770 21363 50828 21369
rect 51626 21332 51632 21344
rect 50080 21304 51632 21332
rect 51626 21292 51632 21304
rect 51684 21292 51690 21344
rect 51920 21341 51948 21508
rect 52641 21471 52699 21477
rect 52641 21437 52653 21471
rect 52687 21437 52699 21471
rect 52641 21431 52699 21437
rect 51905 21335 51963 21341
rect 51905 21301 51917 21335
rect 51951 21301 51963 21335
rect 52656 21332 52684 21431
rect 52730 21428 52736 21480
rect 52788 21468 52794 21480
rect 52917 21471 52975 21477
rect 52788 21440 52833 21468
rect 52788 21428 52794 21440
rect 52917 21437 52929 21471
rect 52963 21468 52975 21471
rect 54110 21468 54116 21480
rect 52963 21440 54116 21468
rect 52963 21437 52975 21440
rect 52917 21431 52975 21437
rect 54110 21428 54116 21440
rect 54168 21428 54174 21480
rect 54220 21477 54248 21508
rect 54297 21505 54309 21539
rect 54343 21505 54355 21539
rect 54478 21536 54484 21548
rect 54439 21508 54484 21536
rect 54297 21499 54355 21505
rect 54205 21471 54263 21477
rect 54205 21437 54217 21471
rect 54251 21437 54263 21471
rect 54312 21468 54340 21499
rect 54478 21496 54484 21508
rect 54536 21496 54542 21548
rect 54772 21536 54800 21576
rect 57701 21539 57759 21545
rect 57701 21536 57713 21539
rect 54772 21508 55260 21536
rect 54312 21440 54984 21468
rect 54205 21431 54263 21437
rect 54220 21400 54248 21431
rect 54570 21400 54576 21412
rect 54220 21372 54576 21400
rect 54570 21360 54576 21372
rect 54628 21360 54634 21412
rect 53282 21332 53288 21344
rect 52656 21304 53288 21332
rect 51905 21295 51963 21301
rect 53282 21292 53288 21304
rect 53340 21292 53346 21344
rect 54018 21292 54024 21344
rect 54076 21332 54082 21344
rect 54481 21335 54539 21341
rect 54481 21332 54493 21335
rect 54076 21304 54493 21332
rect 54076 21292 54082 21304
rect 54481 21301 54493 21304
rect 54527 21301 54539 21335
rect 54956 21332 54984 21440
rect 55030 21428 55036 21480
rect 55088 21468 55094 21480
rect 55125 21471 55183 21477
rect 55125 21468 55137 21471
rect 55088 21440 55137 21468
rect 55088 21428 55094 21440
rect 55125 21437 55137 21440
rect 55171 21437 55183 21471
rect 55232 21468 55260 21508
rect 56152 21508 57713 21536
rect 56152 21468 56180 21508
rect 57701 21505 57713 21508
rect 57747 21505 57759 21539
rect 57701 21499 57759 21505
rect 55232 21440 56180 21468
rect 55125 21431 55183 21437
rect 56594 21428 56600 21480
rect 56652 21468 56658 21480
rect 57517 21471 57575 21477
rect 57517 21468 57529 21471
rect 56652 21440 57529 21468
rect 56652 21428 56658 21440
rect 57517 21437 57529 21440
rect 57563 21437 57575 21471
rect 57517 21431 57575 21437
rect 55392 21403 55450 21409
rect 55392 21369 55404 21403
rect 55438 21400 55450 21403
rect 55490 21400 55496 21412
rect 55438 21372 55496 21400
rect 55438 21369 55450 21372
rect 55392 21363 55450 21369
rect 55490 21360 55496 21372
rect 55548 21360 55554 21412
rect 56042 21332 56048 21344
rect 54956 21304 56048 21332
rect 54481 21295 54539 21301
rect 56042 21292 56048 21304
rect 56100 21332 56106 21344
rect 56505 21335 56563 21341
rect 56505 21332 56517 21335
rect 56100 21304 56517 21332
rect 56100 21292 56106 21304
rect 56505 21301 56517 21304
rect 56551 21301 56563 21335
rect 56505 21295 56563 21301
rect 1104 21242 58880 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 50326 21242
rect 50378 21190 50390 21242
rect 50442 21190 50454 21242
rect 50506 21190 50518 21242
rect 50570 21190 58880 21242
rect 1104 21168 58880 21190
rect 49053 21131 49111 21137
rect 49053 21128 49065 21131
rect 48608 21100 49065 21128
rect 1854 20992 1860 21004
rect 1815 20964 1860 20992
rect 1854 20952 1860 20964
rect 1912 20952 1918 21004
rect 2590 20992 2596 21004
rect 2551 20964 2596 20992
rect 2590 20952 2596 20964
rect 2648 20952 2654 21004
rect 2774 20992 2780 21004
rect 2735 20964 2780 20992
rect 2774 20952 2780 20964
rect 2832 20952 2838 21004
rect 47854 20952 47860 21004
rect 47912 20992 47918 21004
rect 48608 21001 48636 21100
rect 49053 21097 49065 21100
rect 49099 21097 49111 21131
rect 49053 21091 49111 21097
rect 49970 21088 49976 21140
rect 50028 21128 50034 21140
rect 50028 21100 54064 21128
rect 50028 21088 50034 21100
rect 50433 21063 50491 21069
rect 50433 21029 50445 21063
rect 50479 21060 50491 21063
rect 50614 21060 50620 21072
rect 50479 21032 50620 21060
rect 50479 21029 50491 21032
rect 50433 21023 50491 21029
rect 50614 21020 50620 21032
rect 50672 21020 50678 21072
rect 52546 21060 52552 21072
rect 51736 21032 52552 21060
rect 48593 20995 48651 21001
rect 48593 20992 48605 20995
rect 47912 20964 48605 20992
rect 47912 20952 47918 20964
rect 48593 20961 48605 20964
rect 48639 20961 48651 20995
rect 48593 20955 48651 20961
rect 49050 20952 49056 21004
rect 49108 20992 49114 21004
rect 49237 20995 49295 21001
rect 49237 20992 49249 20995
rect 49108 20964 49249 20992
rect 49108 20952 49114 20964
rect 49237 20961 49249 20964
rect 49283 20961 49295 20995
rect 49237 20955 49295 20961
rect 49786 20952 49792 21004
rect 49844 20992 49850 21004
rect 49881 20995 49939 21001
rect 49881 20992 49893 20995
rect 49844 20964 49893 20992
rect 49844 20952 49850 20964
rect 49881 20961 49893 20964
rect 49927 20961 49939 20995
rect 49881 20955 49939 20961
rect 50341 20995 50399 21001
rect 50341 20961 50353 20995
rect 50387 20961 50399 20995
rect 50341 20955 50399 20961
rect 50525 20995 50583 21001
rect 50525 20961 50537 20995
rect 50571 20992 50583 20995
rect 51736 20992 51764 21032
rect 52546 21020 52552 21032
rect 52604 21020 52610 21072
rect 53282 21020 53288 21072
rect 53340 21060 53346 21072
rect 54036 21060 54064 21100
rect 54110 21088 54116 21140
rect 54168 21128 54174 21140
rect 54481 21131 54539 21137
rect 54481 21128 54493 21131
rect 54168 21100 54493 21128
rect 54168 21088 54174 21100
rect 54481 21097 54493 21100
rect 54527 21097 54539 21131
rect 54481 21091 54539 21097
rect 53340 21032 53972 21060
rect 54036 21032 57100 21060
rect 53340 21020 53346 21032
rect 50571 20964 51764 20992
rect 51905 20995 51963 21001
rect 50571 20961 50583 20964
rect 50525 20955 50583 20961
rect 51905 20961 51917 20995
rect 51951 20961 51963 20995
rect 52638 20992 52644 21004
rect 52599 20964 52644 20992
rect 51905 20955 51963 20961
rect 50356 20924 50384 20955
rect 51258 20924 51264 20936
rect 50356 20896 51264 20924
rect 51258 20884 51264 20896
rect 51316 20884 51322 20936
rect 49697 20859 49755 20865
rect 49697 20825 49709 20859
rect 49743 20856 49755 20859
rect 51718 20856 51724 20868
rect 49743 20828 51724 20856
rect 49743 20825 49755 20828
rect 49697 20819 49755 20825
rect 51718 20816 51724 20828
rect 51776 20816 51782 20868
rect 51920 20856 51948 20955
rect 52638 20952 52644 20964
rect 52696 20952 52702 21004
rect 52825 20995 52883 21001
rect 52825 20961 52837 20995
rect 52871 20961 52883 20995
rect 52825 20955 52883 20961
rect 52546 20884 52552 20936
rect 52604 20924 52610 20936
rect 52730 20924 52736 20936
rect 52604 20896 52736 20924
rect 52604 20884 52610 20896
rect 52730 20884 52736 20896
rect 52788 20884 52794 20936
rect 52840 20924 52868 20955
rect 52914 20952 52920 21004
rect 52972 20992 52978 21004
rect 53742 20992 53748 21004
rect 52972 20964 53017 20992
rect 53703 20964 53748 20992
rect 52972 20952 52978 20964
rect 53742 20952 53748 20964
rect 53800 20952 53806 21004
rect 53944 21001 53972 21032
rect 53929 20995 53987 21001
rect 53929 20961 53941 20995
rect 53975 20961 53987 20995
rect 54294 20992 54300 21004
rect 54255 20964 54300 20992
rect 53929 20955 53987 20961
rect 54294 20952 54300 20964
rect 54352 20952 54358 21004
rect 54570 20952 54576 21004
rect 54628 20992 54634 21004
rect 55217 20995 55275 21001
rect 55217 20992 55229 20995
rect 54628 20964 55229 20992
rect 54628 20952 54634 20964
rect 55217 20961 55229 20964
rect 55263 20961 55275 20995
rect 55217 20955 55275 20961
rect 55309 20995 55367 21001
rect 55309 20961 55321 20995
rect 55355 20961 55367 20995
rect 55309 20955 55367 20961
rect 55585 20995 55643 21001
rect 55585 20961 55597 20995
rect 55631 20992 55643 20995
rect 55674 20992 55680 21004
rect 55631 20964 55680 20992
rect 55631 20961 55643 20964
rect 55585 20955 55643 20961
rect 53098 20924 53104 20936
rect 52840 20896 53104 20924
rect 53098 20884 53104 20896
rect 53156 20924 53162 20936
rect 53650 20924 53656 20936
rect 53156 20896 53656 20924
rect 53156 20884 53162 20896
rect 53650 20884 53656 20896
rect 53708 20884 53714 20936
rect 54021 20927 54079 20933
rect 54021 20893 54033 20927
rect 54067 20893 54079 20927
rect 54021 20887 54079 20893
rect 53834 20856 53840 20868
rect 51920 20828 53840 20856
rect 53834 20816 53840 20828
rect 53892 20816 53898 20868
rect 54036 20856 54064 20887
rect 54110 20884 54116 20936
rect 54168 20924 54174 20936
rect 55324 20924 55352 20955
rect 55674 20952 55680 20964
rect 55732 20952 55738 21004
rect 57072 21001 57100 21032
rect 57057 20995 57115 21001
rect 57057 20961 57069 20995
rect 57103 20961 57115 20995
rect 57057 20955 57115 20961
rect 56042 20924 56048 20936
rect 54168 20896 54213 20924
rect 55324 20896 56048 20924
rect 54168 20884 54174 20896
rect 56042 20884 56048 20896
rect 56100 20884 56106 20936
rect 57238 20924 57244 20936
rect 57199 20896 57244 20924
rect 57238 20884 57244 20896
rect 57296 20884 57302 20936
rect 53944 20828 54064 20856
rect 1946 20788 1952 20800
rect 1907 20760 1952 20788
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 48406 20788 48412 20800
rect 48367 20760 48412 20788
rect 48406 20748 48412 20760
rect 48464 20748 48470 20800
rect 51994 20788 52000 20800
rect 51955 20760 52000 20788
rect 51994 20748 52000 20760
rect 52052 20748 52058 20800
rect 52914 20748 52920 20800
rect 52972 20788 52978 20800
rect 53944 20788 53972 20828
rect 54294 20816 54300 20868
rect 54352 20856 54358 20868
rect 56594 20856 56600 20868
rect 54352 20828 56600 20856
rect 54352 20816 54358 20828
rect 56594 20816 56600 20828
rect 56652 20816 56658 20868
rect 52972 20760 53972 20788
rect 52972 20748 52978 20760
rect 54018 20748 54024 20800
rect 54076 20788 54082 20800
rect 55033 20791 55091 20797
rect 55033 20788 55045 20791
rect 54076 20760 55045 20788
rect 54076 20748 54082 20760
rect 55033 20757 55045 20760
rect 55079 20757 55091 20791
rect 55490 20788 55496 20800
rect 55451 20760 55496 20788
rect 55033 20751 55091 20757
rect 55490 20748 55496 20760
rect 55548 20748 55554 20800
rect 57422 20788 57428 20800
rect 57383 20760 57428 20788
rect 57422 20748 57428 20760
rect 57480 20748 57486 20800
rect 1104 20698 58880 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 58880 20698
rect 1104 20624 58880 20646
rect 2409 20587 2467 20593
rect 2409 20553 2421 20587
rect 2455 20584 2467 20587
rect 2590 20584 2596 20596
rect 2455 20556 2596 20584
rect 2455 20553 2467 20556
rect 2409 20547 2467 20553
rect 2590 20544 2596 20556
rect 2648 20544 2654 20596
rect 3234 20584 3240 20596
rect 3195 20556 3240 20584
rect 3234 20544 3240 20556
rect 3292 20544 3298 20596
rect 49881 20587 49939 20593
rect 49881 20553 49893 20587
rect 49927 20584 49939 20587
rect 51258 20584 51264 20596
rect 49927 20556 51074 20584
rect 51219 20556 51264 20584
rect 49927 20553 49939 20556
rect 49881 20547 49939 20553
rect 50341 20519 50399 20525
rect 50341 20485 50353 20519
rect 50387 20485 50399 20519
rect 51046 20516 51074 20556
rect 51258 20544 51264 20556
rect 51316 20544 51322 20596
rect 54294 20584 54300 20596
rect 52472 20556 54300 20584
rect 52472 20516 52500 20556
rect 54294 20544 54300 20556
rect 54352 20544 54358 20596
rect 54478 20544 54484 20596
rect 54536 20584 54542 20596
rect 54849 20587 54907 20593
rect 54849 20584 54861 20587
rect 54536 20556 54861 20584
rect 54536 20544 54542 20556
rect 54849 20553 54861 20556
rect 54895 20553 54907 20587
rect 54849 20547 54907 20553
rect 55401 20587 55459 20593
rect 55401 20553 55413 20587
rect 55447 20584 55459 20587
rect 55674 20584 55680 20596
rect 55447 20556 55680 20584
rect 55447 20553 55459 20556
rect 55401 20547 55459 20553
rect 55674 20544 55680 20556
rect 55732 20544 55738 20596
rect 57238 20516 57244 20528
rect 51046 20488 52500 20516
rect 52564 20488 57244 20516
rect 50341 20479 50399 20485
rect 1949 20451 2007 20457
rect 1949 20417 1961 20451
rect 1995 20448 2007 20451
rect 2866 20448 2872 20460
rect 1995 20420 2872 20448
rect 1995 20417 2007 20420
rect 1949 20411 2007 20417
rect 2866 20408 2872 20420
rect 2924 20408 2930 20460
rect 50356 20448 50384 20479
rect 52564 20448 52592 20488
rect 57238 20476 57244 20488
rect 57296 20476 57302 20528
rect 57425 20519 57483 20525
rect 57425 20485 57437 20519
rect 57471 20516 57483 20519
rect 57514 20516 57520 20528
rect 57471 20488 57520 20516
rect 57471 20485 57483 20488
rect 57425 20479 57483 20485
rect 57514 20476 57520 20488
rect 57572 20476 57578 20528
rect 52822 20448 52828 20460
rect 50356 20420 52592 20448
rect 52783 20420 52828 20448
rect 52822 20408 52828 20420
rect 52880 20408 52886 20460
rect 53009 20451 53067 20457
rect 53009 20417 53021 20451
rect 53055 20448 53067 20451
rect 53282 20448 53288 20460
rect 53055 20420 53288 20448
rect 53055 20417 53067 20420
rect 53009 20411 53067 20417
rect 53282 20408 53288 20420
rect 53340 20408 53346 20460
rect 54588 20420 55352 20448
rect 54588 20392 54616 20420
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 3050 20380 3056 20392
rect 1811 20352 3056 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 3050 20340 3056 20352
rect 3108 20340 3114 20392
rect 3234 20340 3240 20392
rect 3292 20380 3298 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3292 20352 3433 20380
rect 3292 20340 3298 20352
rect 3421 20349 3433 20352
rect 3467 20380 3479 20383
rect 4065 20383 4123 20389
rect 4065 20380 4077 20383
rect 3467 20352 4077 20380
rect 3467 20349 3479 20352
rect 3421 20343 3479 20349
rect 4065 20349 4077 20352
rect 4111 20349 4123 20383
rect 4065 20343 4123 20349
rect 49053 20383 49111 20389
rect 49053 20349 49065 20383
rect 49099 20380 49111 20383
rect 50062 20380 50068 20392
rect 49099 20352 50068 20380
rect 49099 20349 49111 20352
rect 49053 20343 49111 20349
rect 50062 20340 50068 20352
rect 50120 20340 50126 20392
rect 50525 20383 50583 20389
rect 50525 20349 50537 20383
rect 50571 20380 50583 20383
rect 50706 20380 50712 20392
rect 50571 20352 50712 20380
rect 50571 20349 50583 20352
rect 50525 20343 50583 20349
rect 50706 20340 50712 20352
rect 50764 20340 50770 20392
rect 50985 20383 51043 20389
rect 50985 20349 50997 20383
rect 51031 20349 51043 20383
rect 50985 20343 51043 20349
rect 51169 20383 51227 20389
rect 51169 20349 51181 20383
rect 51215 20380 51227 20383
rect 51442 20380 51448 20392
rect 51215 20352 51448 20380
rect 51215 20349 51227 20352
rect 51169 20343 51227 20349
rect 51000 20312 51028 20343
rect 51442 20340 51448 20352
rect 51500 20340 51506 20392
rect 51537 20383 51595 20389
rect 51537 20349 51549 20383
rect 51583 20349 51595 20383
rect 51537 20343 51595 20349
rect 52733 20383 52791 20389
rect 52733 20349 52745 20383
rect 52779 20349 52791 20383
rect 52733 20343 52791 20349
rect 52908 20383 52966 20389
rect 52908 20349 52920 20383
rect 52954 20380 52966 20383
rect 53098 20380 53104 20392
rect 52954 20352 53104 20380
rect 52954 20349 52966 20352
rect 52908 20343 52966 20349
rect 51552 20312 51580 20343
rect 52748 20312 52776 20343
rect 53098 20340 53104 20352
rect 53156 20340 53162 20392
rect 54294 20380 54300 20392
rect 54255 20352 54300 20380
rect 54294 20340 54300 20352
rect 54352 20340 54358 20392
rect 54570 20380 54576 20392
rect 54531 20352 54576 20380
rect 54570 20340 54576 20352
rect 54628 20340 54634 20392
rect 55324 20389 55352 20420
rect 55490 20408 55496 20460
rect 55548 20448 55554 20460
rect 56137 20451 56195 20457
rect 56137 20448 56149 20451
rect 55548 20420 56149 20448
rect 55548 20408 55554 20420
rect 56137 20417 56149 20420
rect 56183 20417 56195 20451
rect 56137 20411 56195 20417
rect 54665 20383 54723 20389
rect 54665 20349 54677 20383
rect 54711 20349 54723 20383
rect 54665 20343 54723 20349
rect 55309 20383 55367 20389
rect 55309 20349 55321 20383
rect 55355 20349 55367 20383
rect 56042 20380 56048 20392
rect 56003 20352 56048 20380
rect 55309 20343 55367 20349
rect 52822 20312 52828 20324
rect 51000 20284 52684 20312
rect 52748 20284 52828 20312
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 50614 20204 50620 20256
rect 50672 20244 50678 20256
rect 50982 20244 50988 20256
rect 50672 20216 50988 20244
rect 50672 20204 50678 20216
rect 50982 20204 50988 20216
rect 51040 20204 51046 20256
rect 51442 20244 51448 20256
rect 51403 20216 51448 20244
rect 51442 20204 51448 20216
rect 51500 20204 51506 20256
rect 52270 20204 52276 20256
rect 52328 20244 52334 20256
rect 52549 20247 52607 20253
rect 52549 20244 52561 20247
rect 52328 20216 52561 20244
rect 52328 20204 52334 20216
rect 52549 20213 52561 20216
rect 52595 20213 52607 20247
rect 52656 20244 52684 20284
rect 52822 20272 52828 20284
rect 52880 20272 52886 20324
rect 53110 20244 53138 20340
rect 54478 20312 54484 20324
rect 54439 20284 54484 20312
rect 54478 20272 54484 20284
rect 54536 20272 54542 20324
rect 54680 20312 54708 20343
rect 56042 20340 56048 20352
rect 56100 20340 56106 20392
rect 57241 20383 57299 20389
rect 57241 20349 57253 20383
rect 57287 20380 57299 20383
rect 57422 20380 57428 20392
rect 57287 20352 57428 20380
rect 57287 20349 57299 20352
rect 57241 20343 57299 20349
rect 57422 20340 57428 20352
rect 57480 20340 57486 20392
rect 56060 20312 56088 20340
rect 57974 20312 57980 20324
rect 54680 20284 56088 20312
rect 57935 20284 57980 20312
rect 57974 20272 57980 20284
rect 58032 20272 58038 20324
rect 58158 20312 58164 20324
rect 58119 20284 58164 20312
rect 58158 20272 58164 20284
rect 58216 20272 58222 20324
rect 52656 20216 53138 20244
rect 52549 20207 52607 20213
rect 54294 20204 54300 20256
rect 54352 20244 54358 20256
rect 55122 20244 55128 20256
rect 54352 20216 55128 20244
rect 54352 20204 54358 20216
rect 55122 20204 55128 20216
rect 55180 20204 55186 20256
rect 1104 20154 58880 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 50326 20154
rect 50378 20102 50390 20154
rect 50442 20102 50454 20154
rect 50506 20102 50518 20154
rect 50570 20102 58880 20154
rect 1104 20080 58880 20102
rect 1854 20000 1860 20052
rect 1912 20040 1918 20052
rect 2409 20043 2467 20049
rect 2409 20040 2421 20043
rect 1912 20012 2421 20040
rect 1912 20000 1918 20012
rect 2409 20009 2421 20012
rect 2455 20009 2467 20043
rect 2409 20003 2467 20009
rect 51442 20000 51448 20052
rect 51500 20040 51506 20052
rect 52181 20043 52239 20049
rect 52181 20040 52193 20043
rect 51500 20012 52193 20040
rect 51500 20000 51506 20012
rect 52181 20009 52193 20012
rect 52227 20009 52239 20043
rect 52181 20003 52239 20009
rect 52270 20000 52276 20052
rect 52328 20040 52334 20052
rect 55306 20040 55312 20052
rect 52328 20012 55312 20040
rect 52328 20000 52334 20012
rect 55306 20000 55312 20012
rect 55364 20000 55370 20052
rect 57974 20000 57980 20052
rect 58032 20040 58038 20052
rect 58161 20043 58219 20049
rect 58161 20040 58173 20043
rect 58032 20012 58173 20040
rect 58032 20000 58038 20012
rect 58161 20009 58173 20012
rect 58207 20009 58219 20043
rect 58161 20003 58219 20009
rect 3878 19972 3884 19984
rect 1964 19944 3884 19972
rect 1964 19913 1992 19944
rect 3878 19932 3884 19944
rect 3936 19932 3942 19984
rect 49896 19944 57560 19972
rect 1949 19907 2007 19913
rect 1949 19873 1961 19907
rect 1995 19873 2007 19907
rect 1949 19867 2007 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 2958 19904 2964 19916
rect 2915 19876 2964 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 49050 19864 49056 19916
rect 49108 19904 49114 19916
rect 49896 19913 49924 19944
rect 49237 19907 49295 19913
rect 49237 19904 49249 19907
rect 49108 19876 49249 19904
rect 49108 19864 49114 19876
rect 49237 19873 49249 19876
rect 49283 19873 49295 19907
rect 49237 19867 49295 19873
rect 49881 19907 49939 19913
rect 49881 19873 49893 19907
rect 49927 19873 49939 19907
rect 49881 19867 49939 19873
rect 50525 19907 50583 19913
rect 50525 19873 50537 19907
rect 50571 19904 50583 19907
rect 50706 19904 50712 19916
rect 50571 19876 50712 19904
rect 50571 19873 50583 19876
rect 50525 19867 50583 19873
rect 50706 19864 50712 19876
rect 50764 19864 50770 19916
rect 50890 19864 50896 19916
rect 50948 19904 50954 19916
rect 51537 19907 51595 19913
rect 51537 19904 51549 19907
rect 50948 19876 51549 19904
rect 50948 19864 50954 19876
rect 51537 19873 51549 19876
rect 51583 19873 51595 19907
rect 52362 19904 52368 19916
rect 52323 19876 52368 19904
rect 51537 19867 51595 19873
rect 52362 19864 52368 19876
rect 52420 19864 52426 19916
rect 52549 19907 52607 19913
rect 52549 19873 52561 19907
rect 52595 19904 52607 19907
rect 53006 19904 53012 19916
rect 52595 19876 53012 19904
rect 52595 19873 52607 19876
rect 52549 19867 52607 19873
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 1780 19768 1808 19799
rect 50062 19796 50068 19848
rect 50120 19836 50126 19848
rect 52270 19836 52276 19848
rect 50120 19808 52276 19836
rect 50120 19796 50126 19808
rect 52270 19796 52276 19808
rect 52328 19796 52334 19848
rect 4433 19771 4491 19777
rect 4433 19768 4445 19771
rect 1780 19740 4445 19768
rect 4433 19737 4445 19740
rect 4479 19737 4491 19771
rect 50614 19768 50620 19780
rect 4433 19731 4491 19737
rect 50080 19740 50620 19768
rect 50080 19712 50108 19740
rect 50614 19728 50620 19740
rect 50672 19768 50678 19780
rect 50890 19768 50896 19780
rect 50672 19740 50896 19768
rect 50672 19728 50678 19740
rect 50890 19728 50896 19740
rect 50948 19728 50954 19780
rect 51442 19728 51448 19780
rect 51500 19768 51506 19780
rect 52564 19768 52592 19867
rect 53006 19864 53012 19876
rect 53064 19864 53070 19916
rect 53098 19864 53104 19916
rect 53156 19904 53162 19916
rect 53374 19913 53380 19916
rect 53156 19876 53201 19904
rect 53156 19864 53162 19876
rect 53368 19867 53380 19913
rect 53432 19904 53438 19916
rect 53432 19876 53468 19904
rect 53374 19864 53380 19867
rect 53432 19864 53438 19876
rect 54754 19864 54760 19916
rect 54812 19904 54818 19916
rect 54941 19907 54999 19913
rect 54941 19904 54953 19907
rect 54812 19876 54953 19904
rect 54812 19864 54818 19876
rect 54941 19873 54953 19876
rect 54987 19873 54999 19907
rect 55122 19904 55128 19916
rect 55083 19876 55128 19904
rect 54941 19867 54999 19873
rect 55122 19864 55128 19876
rect 55180 19864 55186 19916
rect 55214 19864 55220 19916
rect 55272 19904 55278 19916
rect 55585 19907 55643 19913
rect 55585 19904 55597 19907
rect 55272 19876 55597 19904
rect 55272 19864 55278 19876
rect 55585 19873 55597 19876
rect 55631 19873 55643 19907
rect 56870 19904 56876 19916
rect 56831 19876 56876 19904
rect 55585 19867 55643 19873
rect 56870 19864 56876 19876
rect 56928 19864 56934 19916
rect 57532 19913 57560 19944
rect 57517 19907 57575 19913
rect 57517 19873 57529 19907
rect 57563 19873 57575 19907
rect 57517 19867 57575 19873
rect 52641 19839 52699 19845
rect 52641 19805 52653 19839
rect 52687 19805 52699 19839
rect 52641 19799 52699 19805
rect 51500 19740 52592 19768
rect 51500 19728 51506 19740
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 3234 19700 3240 19712
rect 3099 19672 3240 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 3234 19660 3240 19672
rect 3292 19660 3298 19712
rect 49050 19700 49056 19712
rect 49011 19672 49056 19700
rect 49050 19660 49056 19672
rect 49108 19660 49114 19712
rect 50062 19660 50068 19712
rect 50120 19660 50126 19712
rect 50341 19703 50399 19709
rect 50341 19669 50353 19703
rect 50387 19700 50399 19703
rect 50706 19700 50712 19712
rect 50387 19672 50712 19700
rect 50387 19669 50399 19672
rect 50341 19663 50399 19669
rect 50706 19660 50712 19672
rect 50764 19660 50770 19712
rect 51534 19660 51540 19712
rect 51592 19700 51598 19712
rect 51629 19703 51687 19709
rect 51629 19700 51641 19703
rect 51592 19672 51641 19700
rect 51592 19660 51598 19672
rect 51629 19669 51641 19672
rect 51675 19669 51687 19703
rect 52656 19700 52684 19799
rect 54386 19796 54392 19848
rect 54444 19836 54450 19848
rect 57701 19839 57759 19845
rect 57701 19836 57713 19839
rect 54444 19808 57713 19836
rect 54444 19796 54450 19808
rect 57701 19805 57713 19808
rect 57747 19805 57759 19839
rect 57701 19799 57759 19805
rect 55122 19768 55128 19780
rect 54312 19740 55128 19768
rect 54202 19700 54208 19712
rect 52656 19672 54208 19700
rect 51629 19663 51687 19669
rect 54202 19660 54208 19672
rect 54260 19700 54266 19712
rect 54312 19700 54340 19740
rect 55122 19728 55128 19740
rect 55180 19728 55186 19780
rect 57054 19768 57060 19780
rect 57015 19740 57060 19768
rect 57054 19728 57060 19740
rect 57112 19728 57118 19780
rect 54478 19700 54484 19712
rect 54260 19672 54340 19700
rect 54439 19672 54484 19700
rect 54260 19660 54266 19672
rect 54478 19660 54484 19672
rect 54536 19660 54542 19712
rect 54941 19703 54999 19709
rect 54941 19669 54953 19703
rect 54987 19700 54999 19703
rect 55214 19700 55220 19712
rect 54987 19672 55220 19700
rect 54987 19669 54999 19672
rect 54941 19663 54999 19669
rect 55214 19660 55220 19672
rect 55272 19660 55278 19712
rect 55306 19660 55312 19712
rect 55364 19700 55370 19712
rect 55677 19703 55735 19709
rect 55677 19700 55689 19703
rect 55364 19672 55689 19700
rect 55364 19660 55370 19672
rect 55677 19669 55689 19672
rect 55723 19669 55735 19703
rect 55677 19663 55735 19669
rect 1104 19610 58880 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 58880 19610
rect 1104 19536 58880 19558
rect 49605 19499 49663 19505
rect 49605 19465 49617 19499
rect 49651 19496 49663 19499
rect 49651 19468 52316 19496
rect 49651 19465 49663 19468
rect 49605 19459 49663 19465
rect 52288 19428 52316 19468
rect 52362 19456 52368 19508
rect 52420 19496 52426 19508
rect 53098 19496 53104 19508
rect 52420 19468 53104 19496
rect 52420 19456 52426 19468
rect 53098 19456 53104 19468
rect 53156 19456 53162 19508
rect 54294 19456 54300 19508
rect 54352 19496 54358 19508
rect 56321 19499 56379 19505
rect 56321 19496 56333 19499
rect 54352 19468 56333 19496
rect 54352 19456 54358 19468
rect 56321 19465 56333 19468
rect 56367 19465 56379 19499
rect 56321 19459 56379 19465
rect 56870 19456 56876 19508
rect 56928 19496 56934 19508
rect 57333 19499 57391 19505
rect 57333 19496 57345 19499
rect 56928 19468 57345 19496
rect 56928 19456 56934 19468
rect 57333 19465 57345 19468
rect 57379 19465 57391 19499
rect 57333 19459 57391 19465
rect 54386 19428 54392 19440
rect 52288 19400 54392 19428
rect 54386 19388 54392 19400
rect 54444 19388 54450 19440
rect 53282 19360 53288 19372
rect 49896 19332 50384 19360
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 2924 19264 3433 19292
rect 2924 19252 2930 19264
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 47854 19292 47860 19304
rect 47815 19264 47860 19292
rect 3421 19255 3479 19261
rect 47854 19252 47860 19264
rect 47912 19252 47918 19304
rect 49050 19252 49056 19304
rect 49108 19292 49114 19304
rect 49145 19295 49203 19301
rect 49145 19292 49157 19295
rect 49108 19264 49157 19292
rect 49108 19252 49114 19264
rect 49145 19261 49157 19264
rect 49191 19261 49203 19295
rect 49786 19292 49792 19304
rect 49747 19264 49792 19292
rect 49145 19255 49203 19261
rect 49786 19252 49792 19264
rect 49844 19252 49850 19304
rect 1854 19224 1860 19236
rect 1815 19196 1860 19224
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 2590 19224 2596 19236
rect 2551 19196 2596 19224
rect 2590 19184 2596 19196
rect 2648 19184 2654 19236
rect 2774 19224 2780 19236
rect 2735 19196 2780 19224
rect 2774 19184 2780 19196
rect 2832 19184 2838 19236
rect 49896 19224 49924 19332
rect 49970 19252 49976 19304
rect 50028 19292 50034 19304
rect 50249 19295 50307 19301
rect 50249 19292 50261 19295
rect 50028 19264 50261 19292
rect 50028 19252 50034 19264
rect 50249 19261 50261 19264
rect 50295 19261 50307 19295
rect 50356 19292 50384 19332
rect 52840 19332 53288 19360
rect 52086 19292 52092 19304
rect 50356 19264 52092 19292
rect 50249 19255 50307 19261
rect 47688 19196 49924 19224
rect 50264 19224 50292 19255
rect 52086 19252 52092 19264
rect 52144 19252 52150 19304
rect 52840 19301 52868 19332
rect 53282 19320 53288 19332
rect 53340 19320 53346 19372
rect 54570 19320 54576 19372
rect 54628 19320 54634 19372
rect 52733 19295 52791 19301
rect 52733 19261 52745 19295
rect 52779 19261 52791 19295
rect 52733 19255 52791 19261
rect 52822 19295 52880 19301
rect 52822 19261 52834 19295
rect 52868 19261 52880 19295
rect 52822 19255 52880 19261
rect 52917 19295 52975 19301
rect 52917 19261 52929 19295
rect 52963 19261 52975 19295
rect 52917 19255 52975 19261
rect 50516 19227 50574 19233
rect 50264 19196 50384 19224
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 47688 19165 47716 19196
rect 47673 19159 47731 19165
rect 47673 19125 47685 19159
rect 47719 19125 47731 19159
rect 47673 19119 47731 19125
rect 48961 19159 49019 19165
rect 48961 19125 48973 19159
rect 49007 19156 49019 19159
rect 49694 19156 49700 19168
rect 49007 19128 49700 19156
rect 49007 19125 49019 19128
rect 48961 19119 49019 19125
rect 49694 19116 49700 19128
rect 49752 19156 49758 19168
rect 50154 19156 50160 19168
rect 49752 19128 50160 19156
rect 49752 19116 49758 19128
rect 50154 19116 50160 19128
rect 50212 19116 50218 19168
rect 50356 19156 50384 19196
rect 50516 19193 50528 19227
rect 50562 19224 50574 19227
rect 51902 19224 51908 19236
rect 50562 19196 51908 19224
rect 50562 19193 50574 19196
rect 50516 19187 50574 19193
rect 51902 19184 51908 19196
rect 51960 19184 51966 19236
rect 52457 19227 52515 19233
rect 52457 19193 52469 19227
rect 52503 19224 52515 19227
rect 52546 19224 52552 19236
rect 52503 19196 52552 19224
rect 52503 19193 52515 19196
rect 52457 19187 52515 19193
rect 52546 19184 52552 19196
rect 52604 19184 52610 19236
rect 52748 19168 52776 19255
rect 52932 19224 52960 19255
rect 53098 19252 53104 19304
rect 53156 19292 53162 19304
rect 53156 19264 53201 19292
rect 53156 19252 53162 19264
rect 54110 19252 54116 19304
rect 54168 19292 54174 19304
rect 54297 19295 54355 19301
rect 54297 19292 54309 19295
rect 54168 19264 54309 19292
rect 54168 19252 54174 19264
rect 54297 19261 54309 19264
rect 54343 19292 54355 19295
rect 54478 19292 54484 19304
rect 54343 19264 54484 19292
rect 54343 19261 54355 19264
rect 54297 19255 54355 19261
rect 54478 19252 54484 19264
rect 54536 19252 54542 19304
rect 54588 19236 54616 19320
rect 54662 19252 54668 19304
rect 54720 19292 54726 19304
rect 54941 19295 54999 19301
rect 54941 19292 54953 19295
rect 54720 19264 54953 19292
rect 54720 19252 54726 19264
rect 54941 19261 54953 19264
rect 54987 19292 54999 19295
rect 55030 19292 55036 19304
rect 54987 19264 55036 19292
rect 54987 19261 54999 19264
rect 54941 19255 54999 19261
rect 55030 19252 55036 19264
rect 55088 19252 55094 19304
rect 55214 19301 55220 19304
rect 55208 19292 55220 19301
rect 55175 19264 55220 19292
rect 55208 19255 55220 19264
rect 55214 19252 55220 19255
rect 55272 19252 55278 19304
rect 56962 19292 56968 19304
rect 56923 19264 56968 19292
rect 56962 19252 56968 19264
rect 57020 19252 57026 19304
rect 57146 19292 57152 19304
rect 57107 19264 57152 19292
rect 57146 19252 57152 19264
rect 57204 19252 57210 19304
rect 53834 19224 53840 19236
rect 52932 19196 53840 19224
rect 53834 19184 53840 19196
rect 53892 19184 53898 19236
rect 54202 19184 54208 19236
rect 54260 19224 54266 19236
rect 54386 19224 54392 19236
rect 54260 19196 54392 19224
rect 54260 19184 54266 19196
rect 54386 19184 54392 19196
rect 54444 19184 54450 19236
rect 54570 19184 54576 19236
rect 54628 19224 54634 19236
rect 55306 19224 55312 19236
rect 54628 19196 55312 19224
rect 54628 19184 54634 19196
rect 55306 19184 55312 19196
rect 55364 19184 55370 19236
rect 50890 19156 50896 19168
rect 50356 19128 50896 19156
rect 50890 19116 50896 19128
rect 50948 19116 50954 19168
rect 51626 19156 51632 19168
rect 51587 19128 51632 19156
rect 51626 19116 51632 19128
rect 51684 19116 51690 19168
rect 52730 19156 52736 19168
rect 52643 19128 52736 19156
rect 52730 19116 52736 19128
rect 52788 19156 52794 19168
rect 53926 19156 53932 19168
rect 52788 19128 53932 19156
rect 52788 19116 52794 19128
rect 53926 19116 53932 19128
rect 53984 19116 53990 19168
rect 1104 19066 58880 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 50326 19066
rect 50378 19014 50390 19066
rect 50442 19014 50454 19066
rect 50506 19014 50518 19066
rect 50570 19014 58880 19066
rect 1104 18992 58880 19014
rect 2590 18952 2596 18964
rect 2551 18924 2596 18952
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 49053 18955 49111 18961
rect 49053 18921 49065 18955
rect 49099 18952 49111 18955
rect 49970 18952 49976 18964
rect 49099 18924 49976 18952
rect 49099 18921 49111 18924
rect 49053 18915 49111 18921
rect 49970 18912 49976 18924
rect 50028 18912 50034 18964
rect 50706 18912 50712 18964
rect 50764 18952 50770 18964
rect 57146 18952 57152 18964
rect 50764 18924 57152 18952
rect 50764 18912 50770 18924
rect 57146 18912 57152 18924
rect 57204 18912 57210 18964
rect 55214 18884 55220 18896
rect 49712 18856 55220 18884
rect 1949 18819 2007 18825
rect 1949 18785 1961 18819
rect 1995 18816 2007 18819
rect 2866 18816 2872 18828
rect 1995 18788 2872 18816
rect 1995 18785 2007 18788
rect 1949 18779 2007 18785
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 3234 18816 3240 18828
rect 3195 18788 3240 18816
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 49050 18776 49056 18828
rect 49108 18816 49114 18828
rect 49712 18825 49740 18856
rect 55214 18844 55220 18856
rect 55272 18844 55278 18896
rect 56686 18884 56692 18896
rect 55508 18856 56692 18884
rect 49237 18819 49295 18825
rect 49237 18816 49249 18819
rect 49108 18788 49249 18816
rect 49108 18776 49114 18788
rect 49237 18785 49249 18788
rect 49283 18785 49295 18819
rect 49237 18779 49295 18785
rect 49697 18819 49755 18825
rect 49697 18785 49709 18819
rect 49743 18785 49755 18819
rect 49697 18779 49755 18785
rect 49878 18776 49884 18828
rect 49936 18816 49942 18828
rect 50341 18819 50399 18825
rect 50341 18816 50353 18819
rect 49936 18788 50353 18816
rect 49936 18776 49942 18788
rect 50341 18785 50353 18788
rect 50387 18785 50399 18819
rect 50341 18779 50399 18785
rect 50525 18819 50583 18825
rect 50525 18785 50537 18819
rect 50571 18816 50583 18819
rect 51442 18816 51448 18828
rect 50571 18788 51448 18816
rect 50571 18785 50583 18788
rect 50525 18779 50583 18785
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18748 2191 18751
rect 50356 18748 50384 18779
rect 51442 18776 51448 18788
rect 51500 18776 51506 18828
rect 51626 18816 51632 18828
rect 51587 18788 51632 18816
rect 51626 18776 51632 18788
rect 51684 18776 51690 18828
rect 52549 18819 52607 18825
rect 52549 18785 52561 18819
rect 52595 18816 52607 18819
rect 52638 18816 52644 18828
rect 52595 18788 52644 18816
rect 52595 18785 52607 18788
rect 52549 18779 52607 18785
rect 52638 18776 52644 18788
rect 52696 18776 52702 18828
rect 52914 18776 52920 18828
rect 52972 18816 52978 18828
rect 53374 18816 53380 18828
rect 52972 18788 53380 18816
rect 52972 18776 52978 18788
rect 53374 18776 53380 18788
rect 53432 18776 53438 18828
rect 54110 18816 54116 18828
rect 54071 18788 54116 18816
rect 54110 18776 54116 18788
rect 54168 18776 54174 18828
rect 54205 18819 54263 18825
rect 54205 18785 54217 18819
rect 54251 18816 54263 18819
rect 54294 18816 54300 18828
rect 54251 18788 54300 18816
rect 54251 18785 54263 18788
rect 54205 18779 54263 18785
rect 54294 18776 54300 18788
rect 54352 18776 54358 18828
rect 54386 18776 54392 18828
rect 54444 18816 54450 18828
rect 54481 18819 54539 18825
rect 54481 18816 54493 18819
rect 54444 18788 54493 18816
rect 54444 18776 54450 18788
rect 54481 18785 54493 18788
rect 54527 18785 54539 18819
rect 54481 18779 54539 18785
rect 54941 18819 54999 18825
rect 54941 18785 54953 18819
rect 54987 18816 54999 18819
rect 55508 18816 55536 18856
rect 56686 18844 56692 18856
rect 56744 18884 56750 18896
rect 57330 18884 57336 18896
rect 56744 18856 57336 18884
rect 56744 18844 56750 18856
rect 57330 18844 57336 18856
rect 57388 18844 57394 18896
rect 54987 18788 55536 18816
rect 55585 18819 55643 18825
rect 54987 18785 54999 18788
rect 54941 18779 54999 18785
rect 55585 18785 55597 18819
rect 55631 18816 55643 18819
rect 56134 18816 56140 18828
rect 55631 18788 56140 18816
rect 55631 18785 55643 18788
rect 55585 18779 55643 18785
rect 56134 18776 56140 18788
rect 56192 18776 56198 18828
rect 56778 18816 56784 18828
rect 56739 18788 56784 18816
rect 56778 18776 56784 18788
rect 56836 18776 56842 18828
rect 57974 18816 57980 18828
rect 57935 18788 57980 18816
rect 57974 18776 57980 18788
rect 58032 18776 58038 18828
rect 50614 18748 50620 18760
rect 2179 18720 3096 18748
rect 50356 18720 50620 18748
rect 2179 18717 2191 18720
rect 2133 18711 2191 18717
rect 3068 18689 3096 18720
rect 50614 18708 50620 18720
rect 50672 18708 50678 18760
rect 52270 18708 52276 18760
rect 52328 18748 52334 18760
rect 52365 18751 52423 18757
rect 52365 18748 52377 18751
rect 52328 18720 52377 18748
rect 52328 18708 52334 18720
rect 52365 18717 52377 18720
rect 52411 18717 52423 18751
rect 52365 18711 52423 18717
rect 52472 18720 55168 18748
rect 3053 18683 3111 18689
rect 3053 18649 3065 18683
rect 3099 18649 3111 18683
rect 3053 18643 3111 18649
rect 50341 18683 50399 18689
rect 50341 18649 50353 18683
rect 50387 18680 50399 18683
rect 51074 18680 51080 18692
rect 50387 18652 51080 18680
rect 50387 18649 50399 18652
rect 50341 18643 50399 18649
rect 51074 18640 51080 18652
rect 51132 18640 51138 18692
rect 51258 18640 51264 18692
rect 51316 18680 51322 18692
rect 52472 18680 52500 18720
rect 55140 18689 55168 18720
rect 55125 18683 55183 18689
rect 51316 18652 52500 18680
rect 52656 18652 54524 18680
rect 51316 18640 51322 18652
rect 51442 18572 51448 18624
rect 51500 18612 51506 18624
rect 51721 18615 51779 18621
rect 51721 18612 51733 18615
rect 51500 18584 51733 18612
rect 51500 18572 51506 18584
rect 51721 18581 51733 18584
rect 51767 18581 51779 18615
rect 51721 18575 51779 18581
rect 51810 18572 51816 18624
rect 51868 18612 51874 18624
rect 52656 18612 52684 18652
rect 52822 18612 52828 18624
rect 51868 18584 52684 18612
rect 52735 18584 52828 18612
rect 51868 18572 51874 18584
rect 52822 18572 52828 18584
rect 52880 18612 52886 18624
rect 53282 18612 53288 18624
rect 52880 18584 53288 18612
rect 52880 18572 52886 18584
rect 53282 18572 53288 18584
rect 53340 18572 53346 18624
rect 53926 18612 53932 18624
rect 53839 18584 53932 18612
rect 53926 18572 53932 18584
rect 53984 18612 53990 18624
rect 54202 18612 54208 18624
rect 53984 18584 54208 18612
rect 53984 18572 53990 18584
rect 54202 18572 54208 18584
rect 54260 18572 54266 18624
rect 54386 18612 54392 18624
rect 54347 18584 54392 18612
rect 54386 18572 54392 18584
rect 54444 18572 54450 18624
rect 54496 18612 54524 18652
rect 55125 18649 55137 18683
rect 55171 18649 55183 18683
rect 56965 18683 57023 18689
rect 56965 18680 56977 18683
rect 55125 18643 55183 18649
rect 55232 18652 56977 18680
rect 55232 18612 55260 18652
rect 56965 18649 56977 18652
rect 57011 18649 57023 18683
rect 58158 18680 58164 18692
rect 58119 18652 58164 18680
rect 56965 18643 57023 18649
rect 58158 18640 58164 18652
rect 58216 18640 58222 18692
rect 54496 18584 55260 18612
rect 55582 18572 55588 18624
rect 55640 18612 55646 18624
rect 55677 18615 55735 18621
rect 55677 18612 55689 18615
rect 55640 18584 55689 18612
rect 55640 18572 55646 18584
rect 55677 18581 55689 18584
rect 55723 18581 55735 18615
rect 55677 18575 55735 18581
rect 1104 18522 58880 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 58880 18522
rect 1104 18448 58880 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 1949 18411 2007 18417
rect 1949 18408 1961 18411
rect 1912 18380 1961 18408
rect 1912 18368 1918 18380
rect 1949 18377 1961 18380
rect 1995 18377 2007 18411
rect 1949 18371 2007 18377
rect 50617 18411 50675 18417
rect 50617 18377 50629 18411
rect 50663 18408 50675 18411
rect 56134 18408 56140 18420
rect 50663 18380 55720 18408
rect 56095 18380 56140 18408
rect 50663 18377 50675 18380
rect 50617 18371 50675 18377
rect 51442 18340 51448 18352
rect 49988 18312 51448 18340
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 2869 18275 2927 18281
rect 2869 18272 2881 18275
rect 1627 18244 2881 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2869 18241 2881 18244
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 49988 18213 50016 18312
rect 51442 18300 51448 18312
rect 51500 18300 51506 18352
rect 51902 18340 51908 18352
rect 51863 18312 51908 18340
rect 51902 18300 51908 18312
rect 51960 18300 51966 18352
rect 53098 18300 53104 18352
rect 53156 18340 53162 18352
rect 54113 18343 54171 18349
rect 54113 18340 54125 18343
rect 53156 18312 54125 18340
rect 53156 18300 53162 18312
rect 54113 18309 54125 18312
rect 54159 18309 54171 18343
rect 55692 18340 55720 18380
rect 56134 18368 56140 18380
rect 56192 18368 56198 18420
rect 57974 18408 57980 18420
rect 57935 18380 57980 18408
rect 57974 18368 57980 18380
rect 58032 18368 58038 18420
rect 55692 18312 57744 18340
rect 54113 18303 54171 18309
rect 51353 18275 51411 18281
rect 51353 18241 51365 18275
rect 51399 18272 51411 18275
rect 51994 18272 52000 18284
rect 51399 18244 52000 18272
rect 51399 18241 51411 18244
rect 51353 18235 51411 18241
rect 51994 18232 52000 18244
rect 52052 18272 52058 18284
rect 52052 18244 52868 18272
rect 52052 18232 52058 18244
rect 49973 18207 50031 18213
rect 49973 18173 49985 18207
rect 50019 18173 50031 18207
rect 50154 18204 50160 18216
rect 50115 18176 50160 18204
rect 49973 18167 50031 18173
rect 50154 18164 50160 18176
rect 50212 18164 50218 18216
rect 50706 18164 50712 18216
rect 50764 18204 50770 18216
rect 50801 18207 50859 18213
rect 50801 18204 50813 18207
rect 50764 18176 50813 18204
rect 50764 18164 50770 18176
rect 50801 18173 50813 18176
rect 50847 18173 50859 18207
rect 50801 18167 50859 18173
rect 51166 18164 51172 18216
rect 51224 18204 51230 18216
rect 51261 18207 51319 18213
rect 51261 18204 51273 18207
rect 51224 18176 51273 18204
rect 51224 18164 51230 18176
rect 51261 18173 51273 18176
rect 51307 18173 51319 18207
rect 51261 18167 51319 18173
rect 51534 18164 51540 18216
rect 51592 18204 51598 18216
rect 52104 18213 52132 18244
rect 51905 18207 51963 18213
rect 51905 18204 51917 18207
rect 51592 18176 51917 18204
rect 51592 18164 51598 18176
rect 51905 18173 51917 18176
rect 51951 18173 51963 18207
rect 51905 18167 51963 18173
rect 52089 18207 52147 18213
rect 52089 18173 52101 18207
rect 52135 18173 52147 18207
rect 52089 18167 52147 18173
rect 52454 18164 52460 18216
rect 52512 18204 52518 18216
rect 52840 18213 52868 18244
rect 54662 18232 54668 18284
rect 54720 18272 54726 18284
rect 57716 18281 57744 18312
rect 54757 18275 54815 18281
rect 54757 18272 54769 18275
rect 54720 18244 54769 18272
rect 54720 18232 54726 18244
rect 54757 18241 54769 18244
rect 54803 18241 54815 18275
rect 54757 18235 54815 18241
rect 57701 18275 57759 18281
rect 57701 18241 57713 18275
rect 57747 18241 57759 18275
rect 57701 18235 57759 18241
rect 52549 18207 52607 18213
rect 52549 18204 52561 18207
rect 52512 18176 52561 18204
rect 52512 18164 52518 18176
rect 52549 18173 52561 18176
rect 52595 18173 52607 18207
rect 52549 18167 52607 18173
rect 52733 18207 52791 18213
rect 52733 18173 52745 18207
rect 52779 18173 52791 18207
rect 52733 18167 52791 18173
rect 52825 18207 52883 18213
rect 52825 18173 52837 18207
rect 52871 18173 52883 18207
rect 53006 18204 53012 18216
rect 52967 18176 53012 18204
rect 52825 18167 52883 18173
rect 50065 18139 50123 18145
rect 50065 18105 50077 18139
rect 50111 18136 50123 18139
rect 52362 18136 52368 18148
rect 50111 18108 52368 18136
rect 50111 18105 50123 18108
rect 50065 18099 50123 18105
rect 52362 18096 52368 18108
rect 52420 18096 52426 18148
rect 49786 18028 49792 18080
rect 49844 18068 49850 18080
rect 50706 18068 50712 18080
rect 49844 18040 50712 18068
rect 49844 18028 49850 18040
rect 50706 18028 50712 18040
rect 50764 18028 50770 18080
rect 51442 18028 51448 18080
rect 51500 18068 51506 18080
rect 52748 18068 52776 18167
rect 52840 18136 52868 18167
rect 53006 18164 53012 18176
rect 53064 18164 53070 18216
rect 53101 18207 53159 18213
rect 53101 18173 53113 18207
rect 53147 18204 53159 18207
rect 53147 18176 53236 18204
rect 53147 18173 53159 18176
rect 53101 18167 53159 18173
rect 53208 18148 53236 18176
rect 53282 18164 53288 18216
rect 53340 18204 53346 18216
rect 54021 18207 54079 18213
rect 54021 18204 54033 18207
rect 53340 18176 54033 18204
rect 53340 18164 53346 18176
rect 54021 18173 54033 18176
rect 54067 18173 54079 18207
rect 54202 18204 54208 18216
rect 54163 18176 54208 18204
rect 54021 18167 54079 18173
rect 54202 18164 54208 18176
rect 54260 18164 54266 18216
rect 55582 18204 55588 18216
rect 54772 18176 55588 18204
rect 52914 18136 52920 18148
rect 52840 18108 52920 18136
rect 52914 18096 52920 18108
rect 52972 18096 52978 18148
rect 53190 18096 53196 18148
rect 53248 18136 53254 18148
rect 54772 18136 54800 18176
rect 55582 18164 55588 18176
rect 55640 18164 55646 18216
rect 57514 18204 57520 18216
rect 57475 18176 57520 18204
rect 57514 18164 57520 18176
rect 57572 18164 57578 18216
rect 53248 18108 54800 18136
rect 53248 18096 53254 18108
rect 54846 18096 54852 18148
rect 54904 18136 54910 18148
rect 55002 18139 55060 18145
rect 55002 18136 55014 18139
rect 54904 18108 55014 18136
rect 54904 18096 54910 18108
rect 55002 18105 55014 18108
rect 55048 18105 55060 18139
rect 56870 18136 56876 18148
rect 56831 18108 56876 18136
rect 55002 18099 55060 18105
rect 56870 18096 56876 18108
rect 56928 18096 56934 18148
rect 57054 18136 57060 18148
rect 57015 18108 57060 18136
rect 57054 18096 57060 18108
rect 57112 18096 57118 18148
rect 52822 18068 52828 18080
rect 51500 18040 52828 18068
rect 51500 18028 51506 18040
rect 52822 18028 52828 18040
rect 52880 18028 52886 18080
rect 1104 17978 58880 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 50326 17978
rect 50378 17926 50390 17978
rect 50442 17926 50454 17978
rect 50506 17926 50518 17978
rect 50570 17926 58880 17978
rect 1104 17904 58880 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 1820 17836 2513 17864
rect 1820 17824 1826 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 2501 17827 2559 17833
rect 49697 17867 49755 17873
rect 49697 17833 49709 17867
rect 49743 17833 49755 17867
rect 54846 17864 54852 17876
rect 54807 17836 54852 17864
rect 49697 17827 49755 17833
rect 1854 17728 1860 17740
rect 1815 17700 1860 17728
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17728 2743 17731
rect 3234 17728 3240 17740
rect 2731 17700 3240 17728
rect 2731 17697 2743 17700
rect 2685 17691 2743 17697
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 49712 17660 49740 17827
rect 54846 17824 54852 17836
rect 54904 17824 54910 17876
rect 52730 17796 52736 17808
rect 50356 17768 52736 17796
rect 49786 17688 49792 17740
rect 49844 17728 49850 17740
rect 50356 17737 50384 17768
rect 52730 17756 52736 17768
rect 52788 17796 52794 17808
rect 52788 17768 54061 17796
rect 52788 17756 52794 17768
rect 49881 17731 49939 17737
rect 49881 17728 49893 17731
rect 49844 17700 49893 17728
rect 49844 17688 49850 17700
rect 49881 17697 49893 17700
rect 49927 17697 49939 17731
rect 49881 17691 49939 17697
rect 50341 17731 50399 17737
rect 50341 17697 50353 17731
rect 50387 17697 50399 17731
rect 50522 17728 50528 17740
rect 50483 17700 50528 17728
rect 50341 17691 50399 17697
rect 50522 17688 50528 17700
rect 50580 17688 50586 17740
rect 51166 17688 51172 17740
rect 51224 17728 51230 17740
rect 51629 17731 51687 17737
rect 51629 17728 51641 17731
rect 51224 17700 51641 17728
rect 51224 17688 51230 17700
rect 51629 17697 51641 17700
rect 51675 17697 51687 17731
rect 51629 17691 51687 17697
rect 51718 17688 51724 17740
rect 51776 17728 51782 17740
rect 51994 17728 52000 17740
rect 51776 17700 51821 17728
rect 51955 17700 52000 17728
rect 51776 17688 51782 17700
rect 51994 17688 52000 17700
rect 52052 17688 52058 17740
rect 52454 17728 52460 17740
rect 52415 17700 52460 17728
rect 52454 17688 52460 17700
rect 52512 17688 52518 17740
rect 52546 17688 52552 17740
rect 52604 17728 52610 17740
rect 52641 17731 52699 17737
rect 52641 17728 52653 17731
rect 52604 17700 52653 17728
rect 52604 17688 52610 17700
rect 52641 17697 52653 17700
rect 52687 17697 52699 17731
rect 52822 17728 52828 17740
rect 52783 17700 52828 17728
rect 52641 17691 52699 17697
rect 52822 17688 52828 17700
rect 52880 17688 52886 17740
rect 52914 17688 52920 17740
rect 52972 17728 52978 17740
rect 53009 17731 53067 17737
rect 53009 17728 53021 17731
rect 52972 17700 53021 17728
rect 52972 17688 52978 17700
rect 53009 17697 53021 17700
rect 53055 17697 53067 17731
rect 53009 17691 53067 17697
rect 53193 17731 53251 17737
rect 53193 17697 53205 17731
rect 53239 17728 53251 17731
rect 53374 17728 53380 17740
rect 53239 17700 53380 17728
rect 53239 17697 53251 17700
rect 53193 17691 53251 17697
rect 53374 17688 53380 17700
rect 53432 17688 53438 17740
rect 53926 17728 53932 17740
rect 53887 17700 53932 17728
rect 53926 17688 53932 17700
rect 53984 17688 53990 17740
rect 54033 17737 54061 17768
rect 54018 17731 54076 17737
rect 54018 17697 54030 17731
rect 54064 17697 54076 17731
rect 54018 17691 54076 17697
rect 54113 17731 54171 17737
rect 54113 17697 54125 17731
rect 54159 17697 54171 17731
rect 54113 17691 54171 17697
rect 54297 17731 54355 17737
rect 54297 17697 54309 17731
rect 54343 17697 54355 17731
rect 54754 17728 54760 17740
rect 54715 17700 54760 17728
rect 54297 17691 54355 17697
rect 51350 17660 51356 17672
rect 49712 17632 51356 17660
rect 51350 17620 51356 17632
rect 51408 17620 51414 17672
rect 51442 17620 51448 17672
rect 51500 17660 51506 17672
rect 51905 17663 51963 17669
rect 51905 17660 51917 17663
rect 51500 17632 51917 17660
rect 51500 17620 51506 17632
rect 51905 17629 51917 17632
rect 51951 17629 51963 17663
rect 51905 17623 51963 17629
rect 52733 17663 52791 17669
rect 52733 17629 52745 17663
rect 52779 17660 52791 17663
rect 53466 17660 53472 17672
rect 52779 17632 53472 17660
rect 52779 17629 52791 17632
rect 52733 17623 52791 17629
rect 53466 17620 53472 17632
rect 53524 17620 53530 17672
rect 53834 17620 53840 17672
rect 53892 17660 53898 17672
rect 54128 17660 54156 17691
rect 53892 17632 54156 17660
rect 53892 17620 53898 17632
rect 49237 17595 49295 17601
rect 49237 17561 49249 17595
rect 49283 17592 49295 17595
rect 50433 17595 50491 17601
rect 49283 17564 50200 17592
rect 49283 17561 49295 17564
rect 49237 17555 49295 17561
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 50172 17524 50200 17564
rect 50433 17561 50445 17595
rect 50479 17592 50491 17595
rect 52822 17592 52828 17604
rect 50479 17564 52828 17592
rect 50479 17561 50491 17564
rect 50433 17555 50491 17561
rect 52822 17552 52828 17564
rect 52880 17592 52886 17604
rect 54312 17592 54340 17691
rect 54754 17688 54760 17700
rect 54812 17688 54818 17740
rect 54938 17728 54944 17740
rect 54899 17700 54944 17728
rect 54938 17688 54944 17700
rect 54996 17688 55002 17740
rect 55490 17728 55496 17740
rect 55451 17700 55496 17728
rect 55490 17688 55496 17700
rect 55548 17688 55554 17740
rect 54956 17660 54984 17688
rect 55585 17663 55643 17669
rect 55585 17660 55597 17663
rect 54956 17632 55597 17660
rect 55585 17629 55597 17632
rect 55631 17660 55643 17663
rect 56502 17660 56508 17672
rect 55631 17632 56508 17660
rect 55631 17629 55643 17632
rect 55585 17623 55643 17629
rect 56502 17620 56508 17632
rect 56560 17620 56566 17672
rect 56962 17660 56968 17672
rect 56923 17632 56968 17660
rect 56962 17620 56968 17632
rect 57020 17620 57026 17672
rect 57146 17660 57152 17672
rect 57107 17632 57152 17660
rect 57146 17620 57152 17632
rect 57204 17620 57210 17672
rect 52880 17564 54340 17592
rect 52880 17552 52886 17564
rect 56870 17552 56876 17604
rect 56928 17592 56934 17604
rect 57333 17595 57391 17601
rect 57333 17592 57345 17595
rect 56928 17564 57345 17592
rect 56928 17552 56934 17564
rect 57333 17561 57345 17564
rect 57379 17561 57391 17595
rect 57333 17555 57391 17561
rect 51350 17524 51356 17536
rect 50172 17496 51356 17524
rect 51350 17484 51356 17496
rect 51408 17484 51414 17536
rect 51445 17527 51503 17533
rect 51445 17493 51457 17527
rect 51491 17524 51503 17527
rect 51626 17524 51632 17536
rect 51491 17496 51632 17524
rect 51491 17493 51503 17496
rect 51445 17487 51503 17493
rect 51626 17484 51632 17496
rect 51684 17484 51690 17536
rect 53653 17527 53711 17533
rect 53653 17493 53665 17527
rect 53699 17524 53711 17527
rect 54202 17524 54208 17536
rect 53699 17496 54208 17524
rect 53699 17493 53711 17496
rect 53653 17487 53711 17493
rect 54202 17484 54208 17496
rect 54260 17484 54266 17536
rect 54294 17484 54300 17536
rect 54352 17524 54358 17536
rect 57514 17524 57520 17536
rect 54352 17496 57520 17524
rect 54352 17484 54358 17496
rect 57514 17484 57520 17496
rect 57572 17484 57578 17536
rect 1104 17434 58880 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 58880 17434
rect 1104 17360 58880 17382
rect 1854 17280 1860 17332
rect 1912 17320 1918 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1912 17292 1961 17320
rect 1912 17280 1918 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 55214 17320 55220 17332
rect 1949 17283 2007 17289
rect 49160 17292 55220 17320
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17184 1639 17187
rect 2869 17187 2927 17193
rect 2869 17184 2881 17187
rect 1627 17156 2881 17184
rect 1627 17153 1639 17156
rect 1581 17147 1639 17153
rect 2869 17153 2881 17156
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 2498 17116 2504 17128
rect 1811 17088 2504 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 2498 17076 2504 17088
rect 2556 17076 2562 17128
rect 49160 17125 49188 17292
rect 55214 17280 55220 17292
rect 55272 17280 55278 17332
rect 55490 17320 55496 17332
rect 55451 17292 55496 17320
rect 55490 17280 55496 17292
rect 55548 17280 55554 17332
rect 55674 17280 55680 17332
rect 55732 17320 55738 17332
rect 55953 17323 56011 17329
rect 55953 17320 55965 17323
rect 55732 17292 55965 17320
rect 55732 17280 55738 17292
rect 55953 17289 55965 17292
rect 55999 17289 56011 17323
rect 55953 17283 56011 17289
rect 51166 17252 51172 17264
rect 51127 17224 51172 17252
rect 51166 17212 51172 17224
rect 51224 17212 51230 17264
rect 51350 17212 51356 17264
rect 51408 17252 51414 17264
rect 51408 17224 52316 17252
rect 51408 17212 51414 17224
rect 49694 17144 49700 17196
rect 49752 17184 49758 17196
rect 49789 17187 49847 17193
rect 49789 17184 49801 17187
rect 49752 17156 49801 17184
rect 49752 17144 49758 17156
rect 49789 17153 49801 17156
rect 49835 17153 49847 17187
rect 51626 17184 51632 17196
rect 51587 17156 51632 17184
rect 49789 17147 49847 17153
rect 51626 17144 51632 17156
rect 51684 17184 51690 17196
rect 52181 17187 52239 17193
rect 52181 17184 52193 17187
rect 51684 17156 52193 17184
rect 51684 17144 51690 17156
rect 52181 17153 52193 17156
rect 52227 17153 52239 17187
rect 52288 17184 52316 17224
rect 54110 17212 54116 17264
rect 54168 17212 54174 17264
rect 53098 17184 53104 17196
rect 52288 17156 52960 17184
rect 53059 17156 53104 17184
rect 52181 17147 52239 17153
rect 49145 17119 49203 17125
rect 49145 17085 49157 17119
rect 49191 17085 49203 17119
rect 49145 17079 49203 17085
rect 51813 17119 51871 17125
rect 51813 17085 51825 17119
rect 51859 17116 51871 17119
rect 52822 17116 52828 17128
rect 51859 17088 52132 17116
rect 52783 17088 52828 17116
rect 51859 17085 51871 17088
rect 51813 17079 51871 17085
rect 50056 17051 50114 17057
rect 50056 17017 50068 17051
rect 50102 17048 50114 17051
rect 50154 17048 50160 17060
rect 50102 17020 50160 17048
rect 50102 17017 50114 17020
rect 50056 17011 50114 17017
rect 50154 17008 50160 17020
rect 50212 17008 50218 17060
rect 52104 17057 52132 17088
rect 52822 17076 52828 17088
rect 52880 17076 52886 17128
rect 52089 17051 52147 17057
rect 52089 17017 52101 17051
rect 52135 17048 52147 17051
rect 52641 17051 52699 17057
rect 52641 17048 52653 17051
rect 52135 17020 52653 17048
rect 52135 17017 52147 17020
rect 52089 17011 52147 17017
rect 52641 17017 52653 17020
rect 52687 17017 52699 17051
rect 52932 17048 52960 17156
rect 53098 17144 53104 17156
rect 53156 17144 53162 17196
rect 54128 17184 54156 17212
rect 53208 17156 54156 17184
rect 53006 17076 53012 17128
rect 53064 17116 53070 17128
rect 53064 17088 53109 17116
rect 53064 17076 53070 17088
rect 53208 17048 53236 17156
rect 53926 17076 53932 17128
rect 53984 17116 53990 17128
rect 54113 17119 54171 17125
rect 54113 17116 54125 17119
rect 53984 17088 54125 17116
rect 53984 17076 53990 17088
rect 54113 17085 54125 17088
rect 54159 17085 54171 17119
rect 54113 17079 54171 17085
rect 54202 17076 54208 17128
rect 54260 17116 54266 17128
rect 54369 17119 54427 17125
rect 54369 17116 54381 17119
rect 54260 17088 54381 17116
rect 54260 17076 54266 17088
rect 54369 17085 54381 17088
rect 54415 17085 54427 17119
rect 55508 17116 55536 17280
rect 55582 17212 55588 17264
rect 55640 17252 55646 17264
rect 56413 17255 56471 17261
rect 56413 17252 56425 17255
rect 55640 17224 56425 17252
rect 55640 17212 55646 17224
rect 56413 17221 56425 17224
rect 56459 17221 56471 17255
rect 56413 17215 56471 17221
rect 56137 17119 56195 17125
rect 56137 17116 56149 17119
rect 55508 17088 56149 17116
rect 54369 17079 54427 17085
rect 56137 17085 56149 17088
rect 56183 17085 56195 17119
rect 56137 17079 56195 17085
rect 56226 17076 56232 17128
rect 56284 17116 56290 17128
rect 56502 17116 56508 17128
rect 56284 17088 56329 17116
rect 56463 17088 56508 17116
rect 56284 17076 56290 17088
rect 56502 17076 56508 17088
rect 56560 17076 56566 17128
rect 52932 17020 53236 17048
rect 52641 17011 52699 17017
rect 53466 17008 53472 17060
rect 53524 17048 53530 17060
rect 54570 17048 54576 17060
rect 53524 17020 54576 17048
rect 53524 17008 53530 17020
rect 54570 17008 54576 17020
rect 54628 17048 54634 17060
rect 55214 17048 55220 17060
rect 54628 17020 55220 17048
rect 54628 17008 54634 17020
rect 55214 17008 55220 17020
rect 55272 17008 55278 17060
rect 57238 17048 57244 17060
rect 57199 17020 57244 17048
rect 57238 17008 57244 17020
rect 57296 17008 57302 17060
rect 57422 17048 57428 17060
rect 57383 17020 57428 17048
rect 57422 17008 57428 17020
rect 57480 17008 57486 17060
rect 57974 17048 57980 17060
rect 57935 17020 57980 17048
rect 57974 17008 57980 17020
rect 58032 17008 58038 17060
rect 58158 17048 58164 17060
rect 58119 17020 58164 17048
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 50706 16940 50712 16992
rect 50764 16980 50770 16992
rect 51997 16983 52055 16989
rect 51997 16980 52009 16983
rect 50764 16952 52009 16980
rect 50764 16940 50770 16952
rect 51997 16949 52009 16952
rect 52043 16949 52055 16983
rect 51997 16943 52055 16949
rect 52362 16940 52368 16992
rect 52420 16980 52426 16992
rect 56962 16980 56968 16992
rect 52420 16952 56968 16980
rect 52420 16940 52426 16952
rect 56962 16940 56968 16952
rect 57020 16940 57026 16992
rect 1104 16890 58880 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 50326 16890
rect 50378 16838 50390 16890
rect 50442 16838 50454 16890
rect 50506 16838 50518 16890
rect 50570 16838 58880 16890
rect 1104 16816 58880 16838
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 49697 16779 49755 16785
rect 49697 16745 49709 16779
rect 49743 16776 49755 16779
rect 49878 16776 49884 16788
rect 49743 16748 49884 16776
rect 49743 16745 49755 16748
rect 49697 16739 49755 16745
rect 49878 16736 49884 16748
rect 49936 16736 49942 16788
rect 50154 16736 50160 16788
rect 50212 16776 50218 16788
rect 50433 16779 50491 16785
rect 50433 16776 50445 16779
rect 50212 16748 50445 16776
rect 50212 16736 50218 16748
rect 50433 16745 50445 16748
rect 50479 16745 50491 16779
rect 50433 16739 50491 16745
rect 51629 16779 51687 16785
rect 51629 16745 51641 16779
rect 51675 16776 51687 16779
rect 52546 16776 52552 16788
rect 51675 16748 52552 16776
rect 51675 16745 51687 16748
rect 51629 16739 51687 16745
rect 52546 16736 52552 16748
rect 52604 16736 52610 16788
rect 52730 16736 52736 16788
rect 52788 16776 52794 16788
rect 52917 16779 52975 16785
rect 52917 16776 52929 16779
rect 52788 16748 52929 16776
rect 52788 16736 52794 16748
rect 52917 16745 52929 16748
rect 52963 16745 52975 16779
rect 54665 16779 54723 16785
rect 54665 16776 54677 16779
rect 52917 16739 52975 16745
rect 53116 16748 54677 16776
rect 50706 16708 50712 16720
rect 50356 16680 50712 16708
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 3050 16640 3056 16652
rect 2731 16612 3056 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 3050 16600 3056 16612
rect 3108 16640 3114 16652
rect 3329 16643 3387 16649
rect 3329 16640 3341 16643
rect 3108 16612 3341 16640
rect 3108 16600 3114 16612
rect 3329 16609 3341 16612
rect 3375 16609 3387 16643
rect 3329 16603 3387 16609
rect 49881 16643 49939 16649
rect 49881 16609 49893 16643
rect 49927 16640 49939 16643
rect 49970 16640 49976 16652
rect 49927 16612 49976 16640
rect 49927 16609 49939 16612
rect 49881 16603 49939 16609
rect 49970 16600 49976 16612
rect 50028 16600 50034 16652
rect 50356 16649 50384 16680
rect 50706 16668 50712 16680
rect 50764 16668 50770 16720
rect 52089 16711 52147 16717
rect 52089 16677 52101 16711
rect 52135 16708 52147 16711
rect 53006 16708 53012 16720
rect 52135 16680 53012 16708
rect 52135 16677 52147 16680
rect 52089 16671 52147 16677
rect 53006 16668 53012 16680
rect 53064 16668 53070 16720
rect 53116 16652 53144 16748
rect 54665 16745 54677 16748
rect 54711 16745 54723 16779
rect 54665 16739 54723 16745
rect 54754 16736 54760 16788
rect 54812 16776 54818 16788
rect 54812 16748 57744 16776
rect 54812 16736 54818 16748
rect 55309 16711 55367 16717
rect 55309 16708 55321 16711
rect 53852 16680 55321 16708
rect 50341 16643 50399 16649
rect 50341 16609 50353 16643
rect 50387 16609 50399 16643
rect 50341 16603 50399 16609
rect 50525 16643 50583 16649
rect 50525 16609 50537 16643
rect 50571 16640 50583 16643
rect 51350 16640 51356 16652
rect 50571 16612 51356 16640
rect 50571 16609 50583 16612
rect 50525 16603 50583 16609
rect 51350 16600 51356 16612
rect 51408 16600 51414 16652
rect 51442 16600 51448 16652
rect 51500 16640 51506 16652
rect 51626 16640 51632 16652
rect 51500 16612 51545 16640
rect 51587 16612 51632 16640
rect 51500 16600 51506 16612
rect 51626 16600 51632 16612
rect 51684 16600 51690 16652
rect 52270 16640 52276 16652
rect 52183 16612 52276 16640
rect 52270 16600 52276 16612
rect 52328 16640 52334 16652
rect 52822 16640 52828 16652
rect 52328 16612 52828 16640
rect 52328 16600 52334 16612
rect 52822 16600 52828 16612
rect 52880 16600 52886 16652
rect 53098 16640 53104 16652
rect 53011 16612 53104 16640
rect 53098 16600 53104 16612
rect 53156 16600 53162 16652
rect 53377 16643 53435 16649
rect 53377 16609 53389 16643
rect 53423 16640 53435 16643
rect 53423 16612 53696 16640
rect 53423 16609 53435 16612
rect 53377 16603 53435 16609
rect 51166 16532 51172 16584
rect 51224 16572 51230 16584
rect 52914 16572 52920 16584
rect 51224 16544 52920 16572
rect 51224 16532 51230 16544
rect 52914 16532 52920 16544
rect 52972 16532 52978 16584
rect 53190 16572 53196 16584
rect 53151 16544 53196 16572
rect 53190 16532 53196 16544
rect 53248 16532 53254 16584
rect 53282 16532 53288 16584
rect 53340 16572 53346 16584
rect 53668 16572 53696 16612
rect 53852 16572 53880 16680
rect 55309 16677 55321 16680
rect 55355 16677 55367 16711
rect 55309 16671 55367 16677
rect 53929 16643 53987 16649
rect 53929 16609 53941 16643
rect 53975 16640 53987 16643
rect 54202 16640 54208 16652
rect 53975 16612 54208 16640
rect 53975 16609 53987 16612
rect 53929 16603 53987 16609
rect 54202 16600 54208 16612
rect 54260 16600 54266 16652
rect 54478 16600 54484 16652
rect 54536 16640 54542 16652
rect 54573 16643 54631 16649
rect 54573 16640 54585 16643
rect 54536 16612 54585 16640
rect 54536 16600 54542 16612
rect 54573 16609 54585 16612
rect 54619 16609 54631 16643
rect 55214 16640 55220 16652
rect 55175 16612 55220 16640
rect 54573 16603 54631 16609
rect 55214 16600 55220 16612
rect 55272 16600 55278 16652
rect 56594 16600 56600 16652
rect 56652 16640 56658 16652
rect 57716 16649 57744 16748
rect 57974 16736 57980 16788
rect 58032 16776 58038 16788
rect 58161 16779 58219 16785
rect 58161 16776 58173 16779
rect 58032 16748 58173 16776
rect 58032 16736 58038 16748
rect 58161 16745 58173 16748
rect 58207 16745 58219 16779
rect 58161 16739 58219 16745
rect 56689 16643 56747 16649
rect 56689 16640 56701 16643
rect 56652 16612 56701 16640
rect 56652 16600 56658 16612
rect 56689 16609 56701 16612
rect 56735 16609 56747 16643
rect 56689 16603 56747 16609
rect 57701 16643 57759 16649
rect 57701 16609 57713 16643
rect 57747 16609 57759 16643
rect 57701 16603 57759 16609
rect 53340 16544 53385 16572
rect 53668 16544 53880 16572
rect 57517 16575 57575 16581
rect 53340 16532 53346 16544
rect 57517 16541 57529 16575
rect 57563 16541 57575 16575
rect 57517 16535 57575 16541
rect 49237 16507 49295 16513
rect 49237 16473 49249 16507
rect 49283 16504 49295 16507
rect 57532 16504 57560 16535
rect 49283 16476 57560 16504
rect 49283 16473 49295 16476
rect 49237 16467 49295 16473
rect 1946 16436 1952 16448
rect 1907 16408 1952 16436
rect 1946 16396 1952 16408
rect 2004 16396 2010 16448
rect 3142 16436 3148 16448
rect 3103 16408 3148 16436
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 52454 16436 52460 16448
rect 52415 16408 52460 16436
rect 52454 16396 52460 16408
rect 52512 16396 52518 16448
rect 53006 16396 53012 16448
rect 53064 16436 53070 16448
rect 54021 16439 54079 16445
rect 54021 16436 54033 16439
rect 53064 16408 54033 16436
rect 53064 16396 53070 16408
rect 54021 16405 54033 16408
rect 54067 16405 54079 16439
rect 54021 16399 54079 16405
rect 56686 16396 56692 16448
rect 56744 16436 56750 16448
rect 56873 16439 56931 16445
rect 56873 16436 56885 16439
rect 56744 16408 56885 16436
rect 56744 16396 56750 16408
rect 56873 16405 56885 16408
rect 56919 16405 56931 16439
rect 56873 16399 56931 16405
rect 1104 16346 58880 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 58880 16346
rect 1104 16272 58880 16294
rect 1854 16192 1860 16244
rect 1912 16232 1918 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 1912 16204 2237 16232
rect 1912 16192 1918 16204
rect 2225 16201 2237 16204
rect 2271 16201 2283 16235
rect 2225 16195 2283 16201
rect 49605 16235 49663 16241
rect 49605 16201 49617 16235
rect 49651 16232 49663 16235
rect 49651 16204 55076 16232
rect 49651 16201 49663 16204
rect 49605 16195 49663 16201
rect 4709 16167 4767 16173
rect 4709 16164 4721 16167
rect 1872 16136 4721 16164
rect 1872 16105 1900 16136
rect 4709 16133 4721 16136
rect 4755 16133 4767 16167
rect 4709 16127 4767 16133
rect 1857 16099 1915 16105
rect 1857 16065 1869 16099
rect 1903 16065 1915 16099
rect 1857 16059 1915 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 3142 16096 3148 16108
rect 2087 16068 3148 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 52546 16096 52552 16108
rect 52507 16068 52552 16096
rect 52546 16056 52552 16068
rect 52604 16056 52610 16108
rect 52641 16099 52699 16105
rect 52641 16065 52653 16099
rect 52687 16096 52699 16099
rect 53006 16096 53012 16108
rect 52687 16068 53012 16096
rect 52687 16065 52699 16068
rect 52641 16059 52699 16065
rect 53006 16056 53012 16068
rect 53064 16056 53070 16108
rect 53926 16056 53932 16108
rect 53984 16096 53990 16108
rect 54021 16099 54079 16105
rect 54021 16096 54033 16099
rect 53984 16068 54033 16096
rect 53984 16056 53990 16068
rect 54021 16065 54033 16068
rect 54067 16065 54079 16099
rect 55048 16096 55076 16204
rect 57238 16192 57244 16244
rect 57296 16232 57302 16244
rect 57425 16235 57483 16241
rect 57425 16232 57437 16235
rect 57296 16204 57437 16232
rect 57296 16192 57302 16204
rect 57425 16201 57437 16204
rect 57471 16201 57483 16235
rect 57425 16195 57483 16201
rect 57241 16099 57299 16105
rect 57241 16096 57253 16099
rect 55048 16068 57253 16096
rect 54021 16059 54079 16065
rect 57241 16065 57253 16068
rect 57287 16065 57299 16099
rect 57241 16059 57299 16065
rect 3050 15988 3056 16040
rect 3108 16028 3114 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3108 16000 3433 16028
rect 3108 15988 3114 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 4062 16028 4068 16040
rect 4023 16000 4068 16028
rect 3421 15991 3479 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 49789 16031 49847 16037
rect 49789 15997 49801 16031
rect 49835 16028 49847 16031
rect 50249 16031 50307 16037
rect 49835 16000 50016 16028
rect 49835 15997 49847 16000
rect 49789 15991 49847 15997
rect 49988 15904 50016 16000
rect 50249 15997 50261 16031
rect 50295 16028 50307 16031
rect 50798 16028 50804 16040
rect 50295 16000 50804 16028
rect 50295 15997 50307 16000
rect 50249 15991 50307 15997
rect 50798 15988 50804 16000
rect 50856 15988 50862 16040
rect 50985 16031 51043 16037
rect 50985 15997 50997 16031
rect 51031 16028 51043 16031
rect 51258 16028 51264 16040
rect 51031 16000 51264 16028
rect 51031 15997 51043 16000
rect 50985 15991 51043 15997
rect 51258 15988 51264 16000
rect 51316 16028 51322 16040
rect 51626 16028 51632 16040
rect 51316 16000 51632 16028
rect 51316 15988 51322 16000
rect 51626 15988 51632 16000
rect 51684 15988 51690 16040
rect 51994 15988 52000 16040
rect 52052 16028 52058 16040
rect 52089 16031 52147 16037
rect 52089 16028 52101 16031
rect 52052 16000 52101 16028
rect 52052 15988 52058 16000
rect 52089 15997 52101 16000
rect 52135 16028 52147 16031
rect 53282 16028 53288 16040
rect 52135 16000 53288 16028
rect 52135 15997 52147 16000
rect 52089 15991 52147 15997
rect 53282 15988 53288 16000
rect 53340 15988 53346 16040
rect 54036 16028 54064 16059
rect 54846 16028 54852 16040
rect 54036 16000 54852 16028
rect 54846 15988 54852 16000
rect 54904 15988 54910 16040
rect 55674 15988 55680 16040
rect 55732 16028 55738 16040
rect 55953 16031 56011 16037
rect 55953 16028 55965 16031
rect 55732 16000 55965 16028
rect 55732 15988 55738 16000
rect 55953 15997 55965 16000
rect 55999 15997 56011 16031
rect 57057 16031 57115 16037
rect 57057 16028 57069 16031
rect 55953 15991 56011 15997
rect 56060 16000 57069 16028
rect 51169 15963 51227 15969
rect 51169 15929 51181 15963
rect 51215 15960 51227 15963
rect 51350 15960 51356 15972
rect 51215 15932 51356 15960
rect 51215 15929 51227 15932
rect 51169 15923 51227 15929
rect 51350 15920 51356 15932
rect 51408 15920 51414 15972
rect 53006 15920 53012 15972
rect 53064 15960 53070 15972
rect 54266 15963 54324 15969
rect 54266 15960 54278 15963
rect 53064 15932 54278 15960
rect 53064 15920 53070 15932
rect 54266 15929 54278 15932
rect 54312 15929 54324 15963
rect 56060 15960 56088 16000
rect 57057 15997 57069 16000
rect 57103 15997 57115 16031
rect 57057 15991 57115 15997
rect 54266 15923 54324 15929
rect 54404 15932 56088 15960
rect 56321 15963 56379 15969
rect 3234 15892 3240 15904
rect 3195 15864 3240 15892
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 49970 15852 49976 15904
rect 50028 15892 50034 15904
rect 50433 15895 50491 15901
rect 50433 15892 50445 15895
rect 50028 15864 50445 15892
rect 50028 15852 50034 15864
rect 50433 15861 50445 15864
rect 50479 15861 50491 15895
rect 50433 15855 50491 15861
rect 52273 15895 52331 15901
rect 52273 15861 52285 15895
rect 52319 15892 52331 15895
rect 52546 15892 52552 15904
rect 52319 15864 52552 15892
rect 52319 15861 52331 15864
rect 52273 15855 52331 15861
rect 52546 15852 52552 15864
rect 52604 15852 52610 15904
rect 52638 15852 52644 15904
rect 52696 15892 52702 15904
rect 54404 15892 54432 15932
rect 56321 15929 56333 15963
rect 56367 15929 56379 15963
rect 56321 15923 56379 15929
rect 52696 15864 54432 15892
rect 52696 15852 52702 15864
rect 54478 15852 54484 15904
rect 54536 15892 54542 15904
rect 55401 15895 55459 15901
rect 55401 15892 55413 15895
rect 54536 15864 55413 15892
rect 54536 15852 54542 15864
rect 55401 15861 55413 15864
rect 55447 15861 55459 15895
rect 55401 15855 55459 15861
rect 55490 15852 55496 15904
rect 55548 15892 55554 15904
rect 56336 15892 56364 15923
rect 55548 15864 56364 15892
rect 55548 15852 55554 15864
rect 1104 15802 58880 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 50326 15802
rect 50378 15750 50390 15802
rect 50442 15750 50454 15802
rect 50506 15750 50518 15802
rect 50570 15750 58880 15802
rect 1104 15728 58880 15750
rect 51166 15688 51172 15700
rect 50356 15660 51172 15688
rect 1854 15552 1860 15564
rect 1815 15524 1860 15552
rect 1854 15512 1860 15524
rect 1912 15512 1918 15564
rect 2590 15552 2596 15564
rect 2551 15524 2596 15552
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 49694 15552 49700 15564
rect 49655 15524 49700 15552
rect 49694 15512 49700 15524
rect 49752 15512 49758 15564
rect 50356 15561 50384 15660
rect 51166 15648 51172 15660
rect 51224 15648 51230 15700
rect 52638 15688 52644 15700
rect 51552 15660 52644 15688
rect 50433 15623 50491 15629
rect 50433 15589 50445 15623
rect 50479 15620 50491 15623
rect 51552 15620 51580 15660
rect 52638 15648 52644 15660
rect 52696 15648 52702 15700
rect 52825 15691 52883 15697
rect 52825 15657 52837 15691
rect 52871 15688 52883 15691
rect 53006 15688 53012 15700
rect 52871 15660 53012 15688
rect 52871 15657 52883 15660
rect 52825 15651 52883 15657
rect 53006 15648 53012 15660
rect 53064 15648 53070 15700
rect 53282 15648 53288 15700
rect 53340 15688 53346 15700
rect 55122 15688 55128 15700
rect 53340 15660 55128 15688
rect 53340 15648 53346 15660
rect 55122 15648 55128 15660
rect 55180 15648 55186 15700
rect 55950 15648 55956 15700
rect 56008 15688 56014 15700
rect 56318 15688 56324 15700
rect 56008 15660 56324 15688
rect 56008 15648 56014 15660
rect 56318 15648 56324 15660
rect 56376 15688 56382 15700
rect 56873 15691 56931 15697
rect 56873 15688 56885 15691
rect 56376 15660 56885 15688
rect 56376 15648 56382 15660
rect 56873 15657 56885 15660
rect 56919 15657 56931 15691
rect 56873 15651 56931 15657
rect 51902 15620 51908 15632
rect 50479 15592 51580 15620
rect 51644 15592 51908 15620
rect 50479 15589 50491 15592
rect 50433 15583 50491 15589
rect 50341 15555 50399 15561
rect 50341 15521 50353 15555
rect 50387 15521 50399 15555
rect 50341 15515 50399 15521
rect 50525 15555 50583 15561
rect 50525 15521 50537 15555
rect 50571 15552 50583 15555
rect 50706 15552 50712 15564
rect 50571 15524 50712 15552
rect 50571 15521 50583 15524
rect 50525 15515 50583 15521
rect 50706 15512 50712 15524
rect 50764 15512 50770 15564
rect 51644 15561 51672 15592
rect 51902 15580 51908 15592
rect 51960 15580 51966 15632
rect 53834 15620 53840 15632
rect 53300 15592 53840 15620
rect 53300 15564 53328 15592
rect 53834 15580 53840 15592
rect 53892 15580 53898 15632
rect 51629 15555 51687 15561
rect 51629 15521 51641 15555
rect 51675 15521 51687 15555
rect 51994 15552 52000 15564
rect 51955 15524 52000 15552
rect 51629 15515 51687 15521
rect 51994 15512 52000 15524
rect 52052 15512 52058 15564
rect 53006 15512 53012 15564
rect 53064 15561 53070 15564
rect 53064 15555 53113 15561
rect 53064 15521 53067 15555
rect 53101 15521 53113 15555
rect 53064 15515 53113 15521
rect 53190 15555 53248 15561
rect 53190 15521 53202 15555
rect 53236 15521 53248 15555
rect 53190 15515 53248 15521
rect 53064 15512 53070 15515
rect 51445 15487 51503 15493
rect 51445 15453 51457 15487
rect 51491 15484 51503 15487
rect 52012 15484 52040 15512
rect 51491 15456 52040 15484
rect 51491 15453 51503 15456
rect 51445 15447 51503 15453
rect 2774 15416 2780 15428
rect 2735 15388 2780 15416
rect 2774 15376 2780 15388
rect 2832 15376 2838 15428
rect 53208 15360 53236 15515
rect 53282 15512 53288 15564
rect 53340 15552 53346 15564
rect 53340 15524 53385 15552
rect 53340 15512 53346 15524
rect 53466 15512 53472 15564
rect 53524 15552 53530 15564
rect 53929 15555 53987 15561
rect 53524 15524 53569 15552
rect 53524 15512 53530 15524
rect 53929 15521 53941 15555
rect 53975 15552 53987 15555
rect 54478 15552 54484 15564
rect 53975 15524 54484 15552
rect 53975 15521 53987 15524
rect 53929 15515 53987 15521
rect 54478 15512 54484 15524
rect 54536 15512 54542 15564
rect 55033 15555 55091 15561
rect 55033 15521 55045 15555
rect 55079 15552 55091 15555
rect 55214 15552 55220 15564
rect 55079 15524 55220 15552
rect 55079 15521 55091 15524
rect 55033 15515 55091 15521
rect 55214 15512 55220 15524
rect 55272 15512 55278 15564
rect 55674 15512 55680 15564
rect 55732 15552 55738 15564
rect 56594 15552 56600 15564
rect 55732 15524 56600 15552
rect 55732 15512 55738 15524
rect 56594 15512 56600 15524
rect 56652 15552 56658 15564
rect 56689 15555 56747 15561
rect 56689 15552 56701 15555
rect 56652 15524 56701 15552
rect 56652 15512 56658 15524
rect 56689 15521 56701 15524
rect 56735 15521 56747 15555
rect 57974 15552 57980 15564
rect 57935 15524 57980 15552
rect 56689 15515 56747 15521
rect 57974 15512 57980 15524
rect 58032 15512 58038 15564
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 51258 15308 51264 15360
rect 51316 15348 51322 15360
rect 51721 15351 51779 15357
rect 51721 15348 51733 15351
rect 51316 15320 51733 15348
rect 51316 15308 51322 15320
rect 51721 15317 51733 15320
rect 51767 15317 51779 15351
rect 51721 15311 51779 15317
rect 53190 15308 53196 15360
rect 53248 15308 53254 15360
rect 54018 15348 54024 15360
rect 53979 15320 54024 15348
rect 54018 15308 54024 15320
rect 54076 15348 54082 15360
rect 54662 15348 54668 15360
rect 54076 15320 54668 15348
rect 54076 15308 54082 15320
rect 54662 15308 54668 15320
rect 54720 15308 54726 15360
rect 55125 15351 55183 15357
rect 55125 15317 55137 15351
rect 55171 15348 55183 15351
rect 55766 15348 55772 15360
rect 55171 15320 55772 15348
rect 55171 15317 55183 15320
rect 55125 15311 55183 15317
rect 55766 15308 55772 15320
rect 55824 15308 55830 15360
rect 57882 15308 57888 15360
rect 57940 15348 57946 15360
rect 58069 15351 58127 15357
rect 58069 15348 58081 15351
rect 57940 15320 58081 15348
rect 57940 15308 57946 15320
rect 58069 15317 58081 15320
rect 58115 15317 58127 15351
rect 58069 15311 58127 15317
rect 1104 15258 58880 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 58880 15258
rect 1104 15184 58880 15206
rect 2409 15147 2467 15153
rect 2409 15113 2421 15147
rect 2455 15144 2467 15147
rect 2590 15144 2596 15156
rect 2455 15116 2596 15144
rect 2455 15113 2467 15116
rect 2409 15107 2467 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 49973 15147 50031 15153
rect 49973 15113 49985 15147
rect 50019 15144 50031 15147
rect 50019 15116 51856 15144
rect 50019 15113 50031 15116
rect 49973 15107 50031 15113
rect 4062 15076 4068 15088
rect 1780 15048 4068 15076
rect 1780 15017 1808 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 14977 1823 15011
rect 1765 14971 1823 14977
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 3234 15008 3240 15020
rect 1995 14980 3240 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 49786 14968 49792 15020
rect 49844 15008 49850 15020
rect 50433 15011 50491 15017
rect 50433 15008 50445 15011
rect 49844 14980 50445 15008
rect 49844 14968 49850 14980
rect 50433 14977 50445 14980
rect 50479 14977 50491 15011
rect 51828 15008 51856 15116
rect 51902 15104 51908 15156
rect 51960 15144 51966 15156
rect 52273 15147 52331 15153
rect 52273 15144 52285 15147
rect 51960 15116 52285 15144
rect 51960 15104 51966 15116
rect 52273 15113 52285 15116
rect 52319 15113 52331 15147
rect 52273 15107 52331 15113
rect 52454 15104 52460 15156
rect 52512 15144 52518 15156
rect 53466 15144 53472 15156
rect 52512 15116 53472 15144
rect 52512 15104 52518 15116
rect 53466 15104 53472 15116
rect 53524 15104 53530 15156
rect 54570 15144 54576 15156
rect 54531 15116 54576 15144
rect 54570 15104 54576 15116
rect 54628 15104 54634 15156
rect 57974 15144 57980 15156
rect 54772 15116 57744 15144
rect 57935 15116 57980 15144
rect 51994 15036 52000 15088
rect 52052 15076 52058 15088
rect 54772 15076 54800 15116
rect 52052 15048 54800 15076
rect 52052 15036 52058 15048
rect 57716 15017 57744 15116
rect 57974 15104 57980 15116
rect 58032 15104 58038 15156
rect 57701 15011 57759 15017
rect 51828 14980 55260 15008
rect 50433 14971 50491 14977
rect 2869 14943 2927 14949
rect 2869 14909 2881 14943
rect 2915 14940 2927 14943
rect 2958 14940 2964 14952
rect 2915 14912 2964 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 52454 14940 52460 14952
rect 52415 14912 52460 14940
rect 52454 14900 52460 14912
rect 52512 14900 52518 14952
rect 52546 14900 52552 14952
rect 52604 14940 52610 14952
rect 52641 14943 52699 14949
rect 52641 14940 52653 14943
rect 52604 14912 52653 14940
rect 52604 14900 52610 14912
rect 52641 14909 52653 14912
rect 52687 14909 52699 14943
rect 52641 14903 52699 14909
rect 52730 14900 52736 14952
rect 52788 14940 52794 14952
rect 54018 14940 54024 14952
rect 52788 14912 54024 14940
rect 52788 14900 52794 14912
rect 54018 14900 54024 14912
rect 54076 14900 54082 14952
rect 54294 14940 54300 14952
rect 54255 14912 54300 14940
rect 54294 14900 54300 14912
rect 54352 14900 54358 14952
rect 54481 14943 54539 14949
rect 54481 14940 54493 14943
rect 54404 14912 54493 14940
rect 50700 14875 50758 14881
rect 50700 14841 50712 14875
rect 50746 14872 50758 14875
rect 51442 14872 51448 14884
rect 50746 14844 51448 14872
rect 50746 14841 50758 14844
rect 50700 14835 50758 14841
rect 51442 14832 51448 14844
rect 51500 14832 51506 14884
rect 51813 14807 51871 14813
rect 51813 14773 51825 14807
rect 51859 14804 51871 14807
rect 54110 14804 54116 14816
rect 51859 14776 54116 14804
rect 51859 14773 51871 14776
rect 51813 14767 51871 14773
rect 54110 14764 54116 14776
rect 54168 14804 54174 14816
rect 54404 14804 54432 14912
rect 54481 14909 54493 14912
rect 54527 14909 54539 14943
rect 54481 14903 54539 14909
rect 54938 14900 54944 14952
rect 54996 14940 55002 14952
rect 55125 14943 55183 14949
rect 55125 14940 55137 14943
rect 54996 14912 55137 14940
rect 54996 14900 55002 14912
rect 55125 14909 55137 14912
rect 55171 14909 55183 14943
rect 55232 14940 55260 14980
rect 57701 14977 57713 15011
rect 57747 14977 57759 15011
rect 57701 14971 57759 14977
rect 57517 14943 57575 14949
rect 57517 14940 57529 14943
rect 55232 14912 57529 14940
rect 55125 14903 55183 14909
rect 57517 14909 57529 14912
rect 57563 14909 57575 14943
rect 57517 14903 57575 14909
rect 54665 14875 54723 14881
rect 54665 14841 54677 14875
rect 54711 14872 54723 14875
rect 54754 14872 54760 14884
rect 54711 14844 54760 14872
rect 54711 14841 54723 14844
rect 54665 14835 54723 14841
rect 54754 14832 54760 14844
rect 54812 14832 54818 14884
rect 55306 14832 55312 14884
rect 55364 14881 55370 14884
rect 55364 14875 55428 14881
rect 55364 14841 55382 14875
rect 55416 14841 55428 14875
rect 55364 14835 55428 14841
rect 55364 14832 55370 14835
rect 55214 14804 55220 14816
rect 54168 14776 55220 14804
rect 54168 14764 54174 14776
rect 55214 14764 55220 14776
rect 55272 14764 55278 14816
rect 55582 14764 55588 14816
rect 55640 14804 55646 14816
rect 56505 14807 56563 14813
rect 56505 14804 56517 14807
rect 55640 14776 56517 14804
rect 55640 14764 55646 14776
rect 56505 14773 56517 14776
rect 56551 14773 56563 14807
rect 56505 14767 56563 14773
rect 1104 14714 58880 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 50326 14714
rect 50378 14662 50390 14714
rect 50442 14662 50454 14714
rect 50506 14662 50518 14714
rect 50570 14662 58880 14714
rect 1104 14640 58880 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 2501 14603 2559 14609
rect 2501 14600 2513 14603
rect 1912 14572 2513 14600
rect 1912 14560 1918 14572
rect 2501 14569 2513 14572
rect 2547 14569 2559 14603
rect 54018 14600 54024 14612
rect 2501 14563 2559 14569
rect 49712 14572 54024 14600
rect 49712 14473 49740 14572
rect 54018 14560 54024 14572
rect 54076 14560 54082 14612
rect 54202 14600 54208 14612
rect 54163 14572 54208 14600
rect 54202 14560 54208 14572
rect 54260 14560 54266 14612
rect 54294 14560 54300 14612
rect 54352 14600 54358 14612
rect 54570 14600 54576 14612
rect 54352 14572 54576 14600
rect 54352 14560 54358 14572
rect 54570 14560 54576 14572
rect 54628 14600 54634 14612
rect 55582 14600 55588 14612
rect 54628 14572 55588 14600
rect 54628 14560 54634 14572
rect 55582 14560 55588 14572
rect 55640 14560 55646 14612
rect 49789 14535 49847 14541
rect 49789 14501 49801 14535
rect 49835 14532 49847 14535
rect 49835 14504 57284 14532
rect 49835 14501 49847 14504
rect 49789 14495 49847 14501
rect 49697 14467 49755 14473
rect 49697 14433 49709 14467
rect 49743 14433 49755 14467
rect 49697 14427 49755 14433
rect 49881 14467 49939 14473
rect 49881 14433 49893 14467
rect 49927 14433 49939 14467
rect 49881 14427 49939 14433
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14365 1915 14399
rect 1857 14359 1915 14365
rect 2041 14399 2099 14405
rect 2041 14365 2053 14399
rect 2087 14396 2099 14399
rect 2498 14396 2504 14408
rect 2087 14368 2504 14396
rect 2087 14365 2099 14368
rect 2041 14359 2099 14365
rect 1872 14328 1900 14359
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 49896 14396 49924 14427
rect 49970 14424 49976 14476
rect 50028 14464 50034 14476
rect 50525 14467 50583 14473
rect 50525 14464 50537 14467
rect 50028 14436 50537 14464
rect 50028 14424 50034 14436
rect 50525 14433 50537 14436
rect 50571 14433 50583 14467
rect 50525 14427 50583 14433
rect 51258 14424 51264 14476
rect 51316 14464 51322 14476
rect 51445 14467 51503 14473
rect 51445 14464 51457 14467
rect 51316 14436 51457 14464
rect 51316 14424 51322 14436
rect 51445 14433 51457 14436
rect 51491 14433 51503 14467
rect 51445 14427 51503 14433
rect 51629 14467 51687 14473
rect 51629 14433 51641 14467
rect 51675 14433 51687 14467
rect 52362 14464 52368 14476
rect 52323 14436 52368 14464
rect 51629 14427 51687 14433
rect 50246 14396 50252 14408
rect 49896 14368 50252 14396
rect 50246 14356 50252 14368
rect 50304 14356 50310 14408
rect 51350 14356 51356 14408
rect 51408 14396 51414 14408
rect 51644 14396 51672 14427
rect 52362 14424 52368 14436
rect 52420 14424 52426 14476
rect 52638 14473 52644 14476
rect 52632 14427 52644 14473
rect 52696 14464 52702 14476
rect 54386 14464 54392 14476
rect 52696 14436 52732 14464
rect 54347 14436 54392 14464
rect 52638 14424 52644 14427
rect 52696 14424 52702 14436
rect 54386 14424 54392 14436
rect 54444 14424 54450 14476
rect 54478 14424 54484 14476
rect 54536 14464 54542 14476
rect 54536 14436 54581 14464
rect 54536 14424 54542 14436
rect 54662 14424 54668 14476
rect 54720 14464 54726 14476
rect 54757 14467 54815 14473
rect 54757 14464 54769 14467
rect 54720 14436 54769 14464
rect 54720 14424 54726 14436
rect 54757 14433 54769 14436
rect 54803 14433 54815 14467
rect 54757 14427 54815 14433
rect 55214 14424 55220 14476
rect 55272 14464 55278 14476
rect 55401 14467 55459 14473
rect 55401 14464 55413 14467
rect 55272 14436 55413 14464
rect 55272 14424 55278 14436
rect 55401 14433 55413 14436
rect 55447 14433 55459 14467
rect 55401 14427 55459 14433
rect 55493 14467 55551 14473
rect 55493 14433 55505 14467
rect 55539 14464 55551 14467
rect 55582 14464 55588 14476
rect 55539 14436 55588 14464
rect 55539 14433 55551 14436
rect 55493 14427 55551 14433
rect 55582 14424 55588 14436
rect 55640 14424 55646 14476
rect 55766 14464 55772 14476
rect 55727 14436 55772 14464
rect 55766 14424 55772 14436
rect 55824 14464 55830 14476
rect 55950 14464 55956 14476
rect 55824 14436 55956 14464
rect 55824 14424 55830 14436
rect 55950 14424 55956 14436
rect 56008 14424 56014 14476
rect 57256 14473 57284 14504
rect 57241 14467 57299 14473
rect 57241 14433 57253 14467
rect 57287 14433 57299 14467
rect 57241 14427 57299 14433
rect 57425 14399 57483 14405
rect 57425 14396 57437 14399
rect 51408 14368 51672 14396
rect 53668 14368 57437 14396
rect 51408 14356 51414 14368
rect 3970 14328 3976 14340
rect 1872 14300 3976 14328
rect 3970 14288 3976 14300
rect 4028 14288 4034 14340
rect 51442 14328 51448 14340
rect 51403 14300 51448 14328
rect 51442 14288 51448 14300
rect 51500 14288 51506 14340
rect 50341 14263 50399 14269
rect 50341 14229 50353 14263
rect 50387 14260 50399 14263
rect 53668 14260 53696 14368
rect 57425 14365 57437 14368
rect 57471 14365 57483 14399
rect 57425 14359 57483 14365
rect 53745 14331 53803 14337
rect 53745 14297 53757 14331
rect 53791 14328 53803 14331
rect 54478 14328 54484 14340
rect 53791 14300 54484 14328
rect 53791 14297 53803 14300
rect 53745 14291 53803 14297
rect 54478 14288 54484 14300
rect 54536 14288 54542 14340
rect 55677 14331 55735 14337
rect 55677 14328 55689 14331
rect 54588 14300 55689 14328
rect 50387 14232 53696 14260
rect 50387 14229 50399 14232
rect 50341 14223 50399 14229
rect 54018 14220 54024 14272
rect 54076 14260 54082 14272
rect 54588 14260 54616 14300
rect 55677 14297 55689 14300
rect 55723 14297 55735 14331
rect 55677 14291 55735 14297
rect 54076 14232 54616 14260
rect 54076 14220 54082 14232
rect 54662 14220 54668 14272
rect 54720 14260 54726 14272
rect 54720 14232 54765 14260
rect 54720 14220 54726 14232
rect 55122 14220 55128 14272
rect 55180 14260 55186 14272
rect 55217 14263 55275 14269
rect 55217 14260 55229 14263
rect 55180 14232 55229 14260
rect 55180 14220 55186 14232
rect 55217 14229 55229 14232
rect 55263 14229 55275 14263
rect 55217 14223 55275 14229
rect 55766 14220 55772 14272
rect 55824 14260 55830 14272
rect 57609 14263 57667 14269
rect 57609 14260 57621 14263
rect 55824 14232 57621 14260
rect 55824 14220 55830 14232
rect 57609 14229 57621 14232
rect 57655 14229 57667 14263
rect 57609 14223 57667 14229
rect 1104 14170 58880 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 58880 14170
rect 1104 14096 58880 14118
rect 2498 14056 2504 14068
rect 2459 14028 2504 14056
rect 2498 14016 2504 14028
rect 2556 14016 2562 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 49694 14016 49700 14068
rect 49752 14056 49758 14068
rect 50982 14056 50988 14068
rect 49752 14028 50988 14056
rect 49752 14016 49758 14028
rect 50982 14016 50988 14028
rect 51040 14016 51046 14068
rect 51905 14059 51963 14065
rect 51905 14025 51917 14059
rect 51951 14056 51963 14059
rect 51994 14056 52000 14068
rect 51951 14028 52000 14056
rect 51951 14025 51963 14028
rect 51905 14019 51963 14025
rect 51994 14016 52000 14028
rect 52052 14016 52058 14068
rect 52549 14059 52607 14065
rect 52549 14025 52561 14059
rect 52595 14056 52607 14059
rect 52638 14056 52644 14068
rect 52595 14028 52644 14056
rect 52595 14025 52607 14028
rect 52549 14019 52607 14025
rect 52638 14016 52644 14028
rect 52696 14016 52702 14068
rect 53926 14016 53932 14068
rect 53984 14056 53990 14068
rect 54662 14056 54668 14068
rect 53984 14028 54668 14056
rect 53984 14016 53990 14028
rect 54662 14016 54668 14028
rect 54720 14016 54726 14068
rect 54754 13948 54760 14000
rect 54812 13988 54818 14000
rect 55490 13988 55496 14000
rect 54812 13960 54857 13988
rect 55451 13960 55496 13988
rect 54812 13948 54818 13960
rect 55490 13948 55496 13960
rect 55548 13948 55554 14000
rect 57885 13991 57943 13997
rect 57885 13957 57897 13991
rect 57931 13957 57943 13991
rect 57885 13951 57943 13957
rect 49804 13892 51120 13920
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 3050 13852 3056 13864
rect 2731 13824 3056 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 3050 13812 3056 13824
rect 3108 13852 3114 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 3108 13824 3341 13852
rect 3108 13812 3114 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 49142 13852 49148 13864
rect 49103 13824 49148 13852
rect 3329 13815 3387 13821
rect 49142 13812 49148 13824
rect 49200 13812 49206 13864
rect 49804 13861 49832 13892
rect 49789 13855 49847 13861
rect 49789 13821 49801 13855
rect 49835 13821 49847 13855
rect 50430 13852 50436 13864
rect 50391 13824 50436 13852
rect 49789 13815 49847 13821
rect 50430 13812 50436 13824
rect 50488 13812 50494 13864
rect 50617 13855 50675 13861
rect 50617 13821 50629 13855
rect 50663 13852 50675 13855
rect 50706 13852 50712 13864
rect 50663 13824 50712 13852
rect 50663 13821 50675 13824
rect 50617 13815 50675 13821
rect 1857 13787 1915 13793
rect 1857 13753 1869 13787
rect 1903 13784 1915 13787
rect 2038 13784 2044 13796
rect 1903 13756 2044 13784
rect 1903 13753 1915 13756
rect 1857 13747 1915 13753
rect 2038 13744 2044 13756
rect 2096 13744 2102 13796
rect 49418 13744 49424 13796
rect 49476 13784 49482 13796
rect 50246 13784 50252 13796
rect 49476 13756 50252 13784
rect 49476 13744 49482 13756
rect 50246 13744 50252 13756
rect 50304 13784 50310 13796
rect 50632 13784 50660 13815
rect 50706 13812 50712 13824
rect 50764 13812 50770 13864
rect 51092 13852 51120 13892
rect 52914 13880 52920 13932
rect 52972 13920 52978 13932
rect 55674 13920 55680 13932
rect 52972 13892 55680 13920
rect 52972 13880 52978 13892
rect 55674 13880 55680 13892
rect 55732 13880 55738 13932
rect 57900 13920 57928 13951
rect 56888 13892 57928 13920
rect 51258 13852 51264 13864
rect 51092 13824 51264 13852
rect 51258 13812 51264 13824
rect 51316 13812 51322 13864
rect 51353 13855 51411 13861
rect 51353 13821 51365 13855
rect 51399 13852 51411 13855
rect 51534 13852 51540 13864
rect 51399 13824 51540 13852
rect 51399 13821 51411 13824
rect 51353 13815 51411 13821
rect 51534 13812 51540 13824
rect 51592 13852 51598 13864
rect 52086 13852 52092 13864
rect 51592 13824 51948 13852
rect 52047 13824 52092 13852
rect 51592 13812 51598 13824
rect 50304 13756 50660 13784
rect 51169 13787 51227 13793
rect 50304 13744 50310 13756
rect 51169 13753 51181 13787
rect 51215 13784 51227 13787
rect 51626 13784 51632 13796
rect 51215 13756 51632 13784
rect 51215 13753 51227 13756
rect 51169 13747 51227 13753
rect 51626 13744 51632 13756
rect 51684 13744 51690 13796
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 3142 13716 3148 13728
rect 3103 13688 3148 13716
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 50525 13719 50583 13725
rect 50525 13685 50537 13719
rect 50571 13716 50583 13719
rect 51074 13716 51080 13728
rect 50571 13688 51080 13716
rect 50571 13685 50583 13688
rect 50525 13679 50583 13685
rect 51074 13676 51080 13688
rect 51132 13676 51138 13728
rect 51920 13716 51948 13824
rect 52086 13812 52092 13824
rect 52144 13812 52150 13864
rect 52546 13812 52552 13864
rect 52604 13852 52610 13864
rect 52730 13852 52736 13864
rect 52604 13824 52649 13852
rect 52691 13824 52736 13852
rect 52604 13812 52610 13824
rect 52730 13812 52736 13824
rect 52788 13812 52794 13864
rect 54205 13855 54263 13861
rect 54205 13821 54217 13855
rect 54251 13852 54263 13855
rect 54294 13852 54300 13864
rect 54251 13824 54300 13852
rect 54251 13821 54263 13824
rect 54205 13815 54263 13821
rect 54294 13812 54300 13824
rect 54352 13812 54358 13864
rect 54386 13812 54392 13864
rect 54444 13852 54450 13864
rect 54573 13855 54631 13861
rect 54444 13824 54489 13852
rect 54444 13812 54450 13824
rect 54573 13821 54585 13855
rect 54619 13821 54631 13855
rect 54573 13815 54631 13821
rect 55309 13855 55367 13861
rect 55309 13821 55321 13855
rect 55355 13852 55367 13855
rect 55766 13852 55772 13864
rect 55355 13824 55772 13852
rect 55355 13821 55367 13824
rect 55309 13815 55367 13821
rect 54110 13744 54116 13796
rect 54168 13784 54174 13796
rect 54481 13787 54539 13793
rect 54481 13784 54493 13787
rect 54168 13756 54493 13784
rect 54168 13744 54174 13756
rect 54481 13753 54493 13756
rect 54527 13753 54539 13787
rect 54481 13747 54539 13753
rect 54588 13728 54616 13815
rect 55766 13812 55772 13824
rect 55824 13812 55830 13864
rect 56042 13852 56048 13864
rect 56003 13824 56048 13852
rect 56042 13812 56048 13824
rect 56100 13812 56106 13864
rect 56888 13861 56916 13892
rect 56873 13855 56931 13861
rect 56873 13821 56885 13855
rect 56919 13821 56931 13855
rect 57054 13852 57060 13864
rect 57015 13824 57060 13852
rect 56873 13815 56931 13821
rect 57054 13812 57060 13824
rect 57112 13812 57118 13864
rect 57514 13852 57520 13864
rect 57475 13824 57520 13852
rect 57514 13812 57520 13824
rect 57572 13812 57578 13864
rect 57698 13852 57704 13864
rect 57659 13824 57704 13852
rect 57698 13812 57704 13824
rect 57756 13812 57762 13864
rect 52546 13716 52552 13728
rect 51920 13688 52552 13716
rect 52546 13676 52552 13688
rect 52604 13676 52610 13728
rect 54570 13676 54576 13728
rect 54628 13676 54634 13728
rect 56134 13716 56140 13728
rect 56095 13688 56140 13716
rect 56134 13676 56140 13688
rect 56192 13676 56198 13728
rect 1104 13626 58880 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 50326 13626
rect 50378 13574 50390 13626
rect 50442 13574 50454 13626
rect 50506 13574 50518 13626
rect 50570 13574 58880 13626
rect 1104 13552 58880 13574
rect 49697 13515 49755 13521
rect 49697 13481 49709 13515
rect 49743 13512 49755 13515
rect 55306 13512 55312 13524
rect 49743 13484 55214 13512
rect 55267 13484 55312 13512
rect 49743 13481 49755 13484
rect 49697 13475 49755 13481
rect 51074 13404 51080 13456
rect 51132 13444 51138 13456
rect 51905 13447 51963 13453
rect 51905 13444 51917 13447
rect 51132 13416 51580 13444
rect 51132 13404 51138 13416
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 2961 13379 3019 13385
rect 2961 13376 2973 13379
rect 1719 13348 2973 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 2961 13345 2973 13348
rect 3007 13345 3019 13379
rect 5074 13376 5080 13388
rect 5035 13348 5080 13376
rect 2961 13339 3019 13345
rect 5074 13336 5080 13348
rect 5132 13336 5138 13388
rect 47486 13376 47492 13388
rect 26206 13348 47492 13376
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 3142 13308 3148 13320
rect 1903 13280 3148 13308
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 2038 13240 2044 13252
rect 1999 13212 2044 13240
rect 2038 13200 2044 13212
rect 2096 13200 2102 13252
rect 5074 13172 5080 13184
rect 5035 13144 5080 13172
rect 5074 13132 5080 13144
rect 5132 13172 5138 13184
rect 26206 13172 26234 13348
rect 47486 13336 47492 13348
rect 47544 13376 47550 13388
rect 47857 13379 47915 13385
rect 47857 13376 47869 13379
rect 47544 13348 47869 13376
rect 47544 13336 47550 13348
rect 47857 13345 47869 13348
rect 47903 13345 47915 13379
rect 49878 13376 49884 13388
rect 49839 13348 49884 13376
rect 47857 13339 47915 13345
rect 49878 13336 49884 13348
rect 49936 13336 49942 13388
rect 50341 13379 50399 13385
rect 50341 13345 50353 13379
rect 50387 13345 50399 13379
rect 50341 13339 50399 13345
rect 50525 13379 50583 13385
rect 50525 13345 50537 13379
rect 50571 13376 50583 13379
rect 51350 13376 51356 13388
rect 50571 13348 51356 13376
rect 50571 13345 50583 13348
rect 50525 13339 50583 13345
rect 50356 13240 50384 13339
rect 51350 13336 51356 13348
rect 51408 13336 51414 13388
rect 50430 13268 50436 13320
rect 50488 13308 50494 13320
rect 51442 13308 51448 13320
rect 50488 13280 50533 13308
rect 51403 13280 51448 13308
rect 50488 13268 50494 13280
rect 51442 13268 51448 13280
rect 51500 13268 51506 13320
rect 51552 13308 51580 13416
rect 51644 13416 51917 13444
rect 51644 13385 51672 13416
rect 51905 13413 51917 13416
rect 51951 13444 51963 13447
rect 52641 13447 52699 13453
rect 52641 13444 52653 13447
rect 51951 13416 52653 13444
rect 51951 13413 51963 13416
rect 51905 13407 51963 13413
rect 52641 13413 52653 13416
rect 52687 13413 52699 13447
rect 53926 13444 53932 13456
rect 53887 13416 53932 13444
rect 52641 13407 52699 13413
rect 53926 13404 53932 13416
rect 53984 13404 53990 13456
rect 54018 13404 54024 13456
rect 54076 13444 54082 13456
rect 54665 13447 54723 13453
rect 54665 13444 54677 13447
rect 54076 13416 54677 13444
rect 54076 13404 54082 13416
rect 54665 13413 54677 13416
rect 54711 13413 54723 13447
rect 55186 13444 55214 13484
rect 55306 13472 55312 13484
rect 55364 13472 55370 13524
rect 55186 13416 57284 13444
rect 54665 13407 54723 13413
rect 51629 13379 51687 13385
rect 51629 13345 51641 13379
rect 51675 13345 51687 13379
rect 51629 13339 51687 13345
rect 52825 13379 52883 13385
rect 52825 13345 52837 13379
rect 52871 13376 52883 13379
rect 53190 13376 53196 13388
rect 52871 13348 53196 13376
rect 52871 13345 52883 13348
rect 52825 13339 52883 13345
rect 53190 13336 53196 13348
rect 53248 13336 53254 13388
rect 53837 13379 53895 13385
rect 53837 13345 53849 13379
rect 53883 13376 53895 13379
rect 54386 13376 54392 13388
rect 53883 13348 54392 13376
rect 53883 13345 53895 13348
rect 53837 13339 53895 13345
rect 54386 13336 54392 13348
rect 54444 13336 54450 13388
rect 54570 13376 54576 13388
rect 54531 13348 54576 13376
rect 54570 13336 54576 13348
rect 54628 13336 54634 13388
rect 55214 13376 55220 13388
rect 55127 13348 55220 13376
rect 55214 13336 55220 13348
rect 55272 13336 55278 13388
rect 55401 13379 55459 13385
rect 55401 13345 55413 13379
rect 55447 13376 55459 13379
rect 55950 13376 55956 13388
rect 55447 13348 55956 13376
rect 55447 13345 55459 13348
rect 55401 13339 55459 13345
rect 55950 13336 55956 13348
rect 56008 13336 56014 13388
rect 57256 13385 57284 13416
rect 57241 13379 57299 13385
rect 57241 13345 57253 13379
rect 57287 13345 57299 13379
rect 57241 13339 57299 13345
rect 51552 13280 51948 13308
rect 51721 13243 51779 13249
rect 51721 13240 51733 13243
rect 50356 13212 51733 13240
rect 51721 13209 51733 13212
rect 51767 13209 51779 13243
rect 51920 13240 51948 13280
rect 51994 13268 52000 13320
rect 52052 13308 52058 13320
rect 53101 13311 53159 13317
rect 52052 13280 52097 13308
rect 52052 13268 52058 13280
rect 53101 13277 53113 13311
rect 53147 13308 53159 13311
rect 54294 13308 54300 13320
rect 53147 13280 54300 13308
rect 53147 13277 53159 13280
rect 53101 13271 53159 13277
rect 54294 13268 54300 13280
rect 54352 13268 54358 13320
rect 55232 13308 55260 13336
rect 55766 13308 55772 13320
rect 55232 13280 55772 13308
rect 55766 13268 55772 13280
rect 55824 13268 55830 13320
rect 57057 13311 57115 13317
rect 57057 13277 57069 13311
rect 57103 13277 57115 13311
rect 57057 13271 57115 13277
rect 57072 13240 57100 13271
rect 51920 13212 57100 13240
rect 51721 13203 51779 13209
rect 5132 13144 26234 13172
rect 5132 13132 5138 13144
rect 47578 13132 47584 13184
rect 47636 13172 47642 13184
rect 48133 13175 48191 13181
rect 48133 13172 48145 13175
rect 47636 13144 48145 13172
rect 47636 13132 47642 13144
rect 48133 13141 48145 13144
rect 48179 13172 48191 13175
rect 52914 13172 52920 13184
rect 48179 13144 52920 13172
rect 48179 13141 48191 13144
rect 48133 13135 48191 13141
rect 52914 13132 52920 13144
rect 52972 13132 52978 13184
rect 53009 13175 53067 13181
rect 53009 13141 53021 13175
rect 53055 13172 53067 13175
rect 53098 13172 53104 13184
rect 53055 13144 53104 13172
rect 53055 13141 53067 13144
rect 53009 13135 53067 13141
rect 53098 13132 53104 13144
rect 53156 13132 53162 13184
rect 57238 13132 57244 13184
rect 57296 13172 57302 13184
rect 57425 13175 57483 13181
rect 57425 13172 57437 13175
rect 57296 13144 57437 13172
rect 57296 13132 57302 13144
rect 57425 13141 57437 13144
rect 57471 13141 57483 13175
rect 57425 13135 57483 13141
rect 1104 13082 58880 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 58880 13082
rect 1104 13008 58880 13030
rect 2958 12968 2964 12980
rect 2919 12940 2964 12968
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 50982 12968 50988 12980
rect 49804 12940 50988 12968
rect 49804 12841 49832 12940
rect 50982 12928 50988 12940
rect 51040 12928 51046 12980
rect 51442 12928 51448 12980
rect 51500 12968 51506 12980
rect 51994 12968 52000 12980
rect 51500 12940 52000 12968
rect 51500 12928 51506 12940
rect 51994 12928 52000 12940
rect 52052 12968 52058 12980
rect 54202 12968 54208 12980
rect 52052 12940 54208 12968
rect 52052 12928 52058 12940
rect 54202 12928 54208 12940
rect 54260 12928 54266 12980
rect 55214 12968 55220 12980
rect 54496 12940 55220 12968
rect 54496 12900 54524 12940
rect 55214 12928 55220 12940
rect 55272 12928 55278 12980
rect 57330 12968 57336 12980
rect 57291 12940 57336 12968
rect 57330 12928 57336 12940
rect 57388 12928 57394 12980
rect 52840 12872 54524 12900
rect 49789 12835 49847 12841
rect 49789 12801 49801 12835
rect 49835 12801 49847 12835
rect 49789 12795 49847 12801
rect 51258 12792 51264 12844
rect 51316 12832 51322 12844
rect 52840 12832 52868 12872
rect 54294 12832 54300 12844
rect 51316 12804 52868 12832
rect 53024 12804 54300 12832
rect 51316 12792 51322 12804
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 5074 12764 5080 12776
rect 2915 12736 5080 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 49329 12767 49387 12773
rect 49329 12733 49341 12767
rect 49375 12733 49387 12767
rect 49329 12727 49387 12733
rect 50056 12767 50114 12773
rect 50056 12733 50068 12767
rect 50102 12764 50114 12767
rect 50430 12764 50436 12776
rect 50102 12736 50436 12764
rect 50102 12733 50114 12736
rect 50056 12727 50114 12733
rect 1854 12696 1860 12708
rect 1815 12668 1860 12696
rect 1854 12656 1860 12668
rect 1912 12656 1918 12708
rect 49344 12696 49372 12727
rect 50430 12724 50436 12736
rect 50488 12724 50494 12776
rect 51629 12767 51687 12773
rect 51629 12733 51641 12767
rect 51675 12764 51687 12767
rect 51718 12764 51724 12776
rect 51675 12736 51724 12764
rect 51675 12733 51687 12736
rect 51629 12727 51687 12733
rect 51718 12724 51724 12736
rect 51776 12724 51782 12776
rect 51810 12724 51816 12776
rect 51868 12764 51874 12776
rect 52733 12767 52791 12773
rect 52733 12764 52745 12767
rect 51868 12736 52745 12764
rect 51868 12724 51874 12736
rect 52733 12733 52745 12736
rect 52779 12733 52791 12767
rect 52733 12727 52791 12733
rect 52822 12724 52828 12776
rect 52880 12764 52886 12776
rect 53024 12773 53052 12804
rect 54294 12792 54300 12804
rect 54352 12792 54358 12844
rect 54938 12792 54944 12844
rect 54996 12832 55002 12844
rect 55033 12835 55091 12841
rect 55033 12832 55045 12835
rect 54996 12804 55045 12832
rect 54996 12792 55002 12804
rect 55033 12801 55045 12804
rect 55079 12801 55091 12835
rect 57514 12832 57520 12844
rect 55033 12795 55091 12801
rect 56060 12804 57520 12832
rect 53009 12767 53067 12773
rect 52880 12736 52925 12764
rect 52880 12724 52886 12736
rect 53009 12733 53021 12767
rect 53055 12733 53067 12767
rect 53009 12727 53067 12733
rect 53098 12724 53104 12776
rect 53156 12764 53162 12776
rect 53156 12736 53201 12764
rect 53156 12724 53162 12736
rect 53926 12724 53932 12776
rect 53984 12764 53990 12776
rect 54021 12767 54079 12773
rect 54021 12764 54033 12767
rect 53984 12736 54033 12764
rect 53984 12724 53990 12736
rect 54021 12733 54033 12736
rect 54067 12733 54079 12767
rect 54202 12764 54208 12776
rect 54163 12736 54208 12764
rect 54021 12727 54079 12733
rect 54202 12724 54208 12736
rect 54260 12724 54266 12776
rect 56060 12764 56088 12804
rect 57514 12792 57520 12804
rect 57572 12792 57578 12844
rect 57238 12764 57244 12776
rect 55140 12736 56088 12764
rect 57199 12736 57244 12764
rect 55140 12696 55168 12736
rect 57238 12724 57244 12736
rect 57296 12724 57302 12776
rect 49344 12668 55168 12696
rect 55300 12699 55358 12705
rect 55300 12665 55312 12699
rect 55346 12696 55358 12699
rect 55582 12696 55588 12708
rect 55346 12668 55588 12696
rect 55346 12665 55358 12668
rect 55300 12659 55358 12665
rect 55582 12656 55588 12668
rect 55640 12656 55646 12708
rect 57974 12696 57980 12708
rect 57935 12668 57980 12696
rect 57974 12656 57980 12668
rect 58032 12656 58038 12708
rect 1946 12628 1952 12640
rect 1907 12600 1952 12628
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 51166 12628 51172 12640
rect 51127 12600 51172 12628
rect 51166 12588 51172 12600
rect 51224 12588 51230 12640
rect 51721 12631 51779 12637
rect 51721 12597 51733 12631
rect 51767 12628 51779 12631
rect 51810 12628 51816 12640
rect 51767 12600 51816 12628
rect 51767 12597 51779 12600
rect 51721 12591 51779 12597
rect 51810 12588 51816 12600
rect 51868 12588 51874 12640
rect 52454 12588 52460 12640
rect 52512 12628 52518 12640
rect 52549 12631 52607 12637
rect 52549 12628 52561 12631
rect 52512 12600 52561 12628
rect 52512 12588 52518 12600
rect 52549 12597 52561 12600
rect 52595 12597 52607 12631
rect 52549 12591 52607 12597
rect 52638 12588 52644 12640
rect 52696 12628 52702 12640
rect 53098 12628 53104 12640
rect 52696 12600 53104 12628
rect 52696 12588 52702 12600
rect 53098 12588 53104 12600
rect 53156 12628 53162 12640
rect 53558 12628 53564 12640
rect 53156 12600 53564 12628
rect 53156 12588 53162 12600
rect 53558 12588 53564 12600
rect 53616 12588 53622 12640
rect 53650 12588 53656 12640
rect 53708 12628 53714 12640
rect 54113 12631 54171 12637
rect 54113 12628 54125 12631
rect 53708 12600 54125 12628
rect 53708 12588 53714 12600
rect 54113 12597 54125 12600
rect 54159 12597 54171 12631
rect 54113 12591 54171 12597
rect 54846 12588 54852 12640
rect 54904 12628 54910 12640
rect 56413 12631 56471 12637
rect 56413 12628 56425 12631
rect 54904 12600 56425 12628
rect 54904 12588 54910 12600
rect 56413 12597 56425 12600
rect 56459 12628 56471 12631
rect 56686 12628 56692 12640
rect 56459 12600 56692 12628
rect 56459 12597 56471 12600
rect 56413 12591 56471 12597
rect 56686 12588 56692 12600
rect 56744 12588 56750 12640
rect 57882 12588 57888 12640
rect 57940 12628 57946 12640
rect 58069 12631 58127 12637
rect 58069 12628 58081 12631
rect 57940 12600 58081 12628
rect 57940 12588 57946 12600
rect 58069 12597 58081 12600
rect 58115 12597 58127 12631
rect 58069 12591 58127 12597
rect 1104 12538 58880 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 50326 12538
rect 50378 12486 50390 12538
rect 50442 12486 50454 12538
rect 50506 12486 50518 12538
rect 50570 12486 58880 12538
rect 1104 12464 58880 12486
rect 51445 12427 51503 12433
rect 51445 12393 51457 12427
rect 51491 12424 51503 12427
rect 51994 12424 52000 12436
rect 51491 12396 52000 12424
rect 51491 12393 51503 12396
rect 51445 12387 51503 12393
rect 51994 12384 52000 12396
rect 52052 12384 52058 12436
rect 52362 12384 52368 12436
rect 52420 12424 52426 12436
rect 52420 12396 54064 12424
rect 52420 12384 52426 12396
rect 50433 12359 50491 12365
rect 50433 12325 50445 12359
rect 50479 12356 50491 12359
rect 52549 12359 52607 12365
rect 50479 12328 52224 12356
rect 50479 12325 50491 12328
rect 50433 12319 50491 12325
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 2685 12291 2743 12297
rect 1627 12260 2636 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 1762 12220 1768 12232
rect 1723 12192 1768 12220
rect 1762 12180 1768 12192
rect 1820 12180 1826 12232
rect 2608 12220 2636 12260
rect 2685 12257 2697 12291
rect 2731 12288 2743 12291
rect 2958 12288 2964 12300
rect 2731 12260 2964 12288
rect 2731 12257 2743 12260
rect 2685 12251 2743 12257
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 49878 12288 49884 12300
rect 49839 12260 49884 12288
rect 49878 12248 49884 12260
rect 49936 12248 49942 12300
rect 50341 12291 50399 12297
rect 50341 12257 50353 12291
rect 50387 12257 50399 12291
rect 50522 12288 50528 12300
rect 50483 12260 50528 12288
rect 50341 12251 50399 12257
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 2608 12192 4445 12220
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 50356 12220 50384 12251
rect 50522 12248 50528 12260
rect 50580 12248 50586 12300
rect 51166 12248 51172 12300
rect 51224 12288 51230 12300
rect 51629 12291 51687 12297
rect 51629 12288 51641 12291
rect 51224 12260 51641 12288
rect 51224 12248 51230 12260
rect 51629 12257 51641 12260
rect 51675 12257 51687 12291
rect 51629 12251 51687 12257
rect 51718 12248 51724 12300
rect 51776 12288 51782 12300
rect 51994 12288 52000 12300
rect 51776 12260 51821 12288
rect 51955 12260 52000 12288
rect 51776 12248 51782 12260
rect 51994 12248 52000 12260
rect 52052 12248 52058 12300
rect 50890 12220 50896 12232
rect 50356 12192 50896 12220
rect 4433 12183 4491 12189
rect 50890 12180 50896 12192
rect 50948 12180 50954 12232
rect 51074 12180 51080 12232
rect 51132 12220 51138 12232
rect 51810 12220 51816 12232
rect 51132 12192 51816 12220
rect 51132 12180 51138 12192
rect 51810 12180 51816 12192
rect 51868 12220 51874 12232
rect 51905 12223 51963 12229
rect 51905 12220 51917 12223
rect 51868 12192 51917 12220
rect 51868 12180 51874 12192
rect 51905 12189 51917 12192
rect 51951 12189 51963 12223
rect 52196 12220 52224 12328
rect 52549 12325 52561 12359
rect 52595 12356 52607 12359
rect 53898 12359 53956 12365
rect 53898 12356 53910 12359
rect 52595 12328 53910 12356
rect 52595 12325 52607 12328
rect 52549 12319 52607 12325
rect 53898 12325 53910 12328
rect 53944 12325 53956 12359
rect 54036 12356 54064 12396
rect 54294 12384 54300 12436
rect 54352 12424 54358 12436
rect 55122 12424 55128 12436
rect 54352 12396 55128 12424
rect 54352 12384 54358 12396
rect 55122 12384 55128 12396
rect 55180 12424 55186 12436
rect 55585 12427 55643 12433
rect 55585 12424 55597 12427
rect 55180 12396 55597 12424
rect 55180 12384 55186 12396
rect 55585 12393 55597 12396
rect 55631 12393 55643 12427
rect 55585 12387 55643 12393
rect 57974 12384 57980 12436
rect 58032 12424 58038 12436
rect 58161 12427 58219 12433
rect 58161 12424 58173 12427
rect 58032 12396 58173 12424
rect 58032 12384 58038 12396
rect 58161 12393 58173 12396
rect 58207 12393 58219 12427
rect 58161 12387 58219 12393
rect 54036 12328 57560 12356
rect 53898 12319 53956 12325
rect 52270 12248 52276 12300
rect 52328 12288 52334 12300
rect 52779 12291 52837 12297
rect 52779 12288 52791 12291
rect 52328 12260 52791 12288
rect 52328 12248 52334 12260
rect 52779 12257 52791 12260
rect 52825 12257 52837 12291
rect 52914 12288 52920 12300
rect 52875 12260 52920 12288
rect 52779 12251 52837 12257
rect 52914 12248 52920 12260
rect 52972 12248 52978 12300
rect 53006 12248 53012 12300
rect 53064 12288 53070 12300
rect 53064 12260 53109 12288
rect 53064 12248 53070 12260
rect 53190 12248 53196 12300
rect 53248 12288 53254 12300
rect 53653 12291 53711 12297
rect 53248 12260 53341 12288
rect 53248 12248 53254 12260
rect 53653 12257 53665 12291
rect 53699 12288 53711 12291
rect 54202 12288 54208 12300
rect 53699 12260 54208 12288
rect 53699 12257 53711 12260
rect 53653 12251 53711 12257
rect 54202 12248 54208 12260
rect 54260 12288 54266 12300
rect 54938 12288 54944 12300
rect 54260 12260 54944 12288
rect 54260 12248 54266 12260
rect 54938 12248 54944 12260
rect 54996 12248 55002 12300
rect 55493 12291 55551 12297
rect 55493 12257 55505 12291
rect 55539 12257 55551 12291
rect 56686 12288 56692 12300
rect 56647 12260 56692 12288
rect 55493 12251 55551 12257
rect 53208 12220 53236 12248
rect 52196 12192 53236 12220
rect 51905 12183 51963 12189
rect 1854 12112 1860 12164
rect 1912 12152 1918 12164
rect 1949 12155 2007 12161
rect 1949 12152 1961 12155
rect 1912 12124 1961 12152
rect 1912 12112 1918 12124
rect 1949 12121 1961 12124
rect 1995 12121 2007 12155
rect 1949 12115 2007 12121
rect 49697 12155 49755 12161
rect 49697 12121 49709 12155
rect 49743 12152 49755 12155
rect 53466 12152 53472 12164
rect 49743 12124 53472 12152
rect 49743 12121 49755 12124
rect 49697 12115 49755 12121
rect 53466 12112 53472 12124
rect 53524 12112 53530 12164
rect 54754 12112 54760 12164
rect 54812 12152 54818 12164
rect 55033 12155 55091 12161
rect 55033 12152 55045 12155
rect 54812 12124 55045 12152
rect 54812 12112 54818 12124
rect 55033 12121 55045 12124
rect 55079 12152 55091 12155
rect 55508 12152 55536 12251
rect 56686 12248 56692 12260
rect 56744 12248 56750 12300
rect 57532 12297 57560 12328
rect 57517 12291 57575 12297
rect 57517 12257 57529 12291
rect 57563 12257 57575 12291
rect 57517 12251 57575 12257
rect 57606 12180 57612 12232
rect 57664 12220 57670 12232
rect 57701 12223 57759 12229
rect 57701 12220 57713 12223
rect 57664 12192 57713 12220
rect 57664 12180 57670 12192
rect 57701 12189 57713 12192
rect 57747 12189 57759 12223
rect 57701 12183 57759 12189
rect 55079 12124 55536 12152
rect 55079 12121 55091 12124
rect 55033 12115 55091 12121
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 49878 12044 49884 12096
rect 49936 12084 49942 12096
rect 50798 12084 50804 12096
rect 49936 12056 50804 12084
rect 49936 12044 49942 12056
rect 50798 12044 50804 12056
rect 50856 12044 50862 12096
rect 50890 12044 50896 12096
rect 50948 12084 50954 12096
rect 52914 12084 52920 12096
rect 50948 12056 52920 12084
rect 50948 12044 50954 12056
rect 52914 12044 52920 12056
rect 52972 12084 52978 12096
rect 54570 12084 54576 12096
rect 52972 12056 54576 12084
rect 52972 12044 52978 12056
rect 54570 12044 54576 12056
rect 54628 12044 54634 12096
rect 55398 12044 55404 12096
rect 55456 12084 55462 12096
rect 56781 12087 56839 12093
rect 56781 12084 56793 12087
rect 55456 12056 56793 12084
rect 55456 12044 55462 12056
rect 56781 12053 56793 12056
rect 56827 12053 56839 12087
rect 56781 12047 56839 12053
rect 1104 11994 58880 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 58880 11994
rect 1104 11920 58880 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 1820 11852 3249 11880
rect 1820 11840 1826 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 51074 11880 51080 11892
rect 3237 11843 3295 11849
rect 49252 11852 51080 11880
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 2924 11648 3433 11676
rect 2924 11636 2930 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 3421 11639 3479 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 49252 11685 49280 11852
rect 51074 11840 51080 11852
rect 51132 11840 51138 11892
rect 51261 11883 51319 11889
rect 51261 11849 51273 11883
rect 51307 11880 51319 11883
rect 51718 11880 51724 11892
rect 51307 11852 51724 11880
rect 51307 11849 51319 11852
rect 51261 11843 51319 11849
rect 51718 11840 51724 11852
rect 51776 11840 51782 11892
rect 51813 11883 51871 11889
rect 51813 11849 51825 11883
rect 51859 11880 51871 11883
rect 51994 11880 52000 11892
rect 51859 11852 52000 11880
rect 51859 11849 51871 11852
rect 51813 11843 51871 11849
rect 51994 11840 52000 11852
rect 52052 11880 52058 11892
rect 52822 11880 52828 11892
rect 52052 11852 52828 11880
rect 52052 11840 52058 11852
rect 52822 11840 52828 11852
rect 52880 11840 52886 11892
rect 53558 11840 53564 11892
rect 53616 11880 53622 11892
rect 55033 11883 55091 11889
rect 55033 11880 55045 11883
rect 53616 11852 55045 11880
rect 53616 11840 53622 11852
rect 55033 11849 55045 11852
rect 55079 11880 55091 11883
rect 55398 11880 55404 11892
rect 55079 11852 55404 11880
rect 55079 11849 55091 11852
rect 55033 11843 55091 11849
rect 55398 11840 55404 11852
rect 55456 11840 55462 11892
rect 55582 11880 55588 11892
rect 55543 11852 55588 11880
rect 55582 11840 55588 11852
rect 55640 11840 55646 11892
rect 51092 11812 51120 11840
rect 51092 11784 52776 11812
rect 52748 11753 52776 11784
rect 53926 11772 53932 11824
rect 53984 11812 53990 11824
rect 54573 11815 54631 11821
rect 54573 11812 54585 11815
rect 53984 11784 54585 11812
rect 53984 11772 53990 11784
rect 54573 11781 54585 11784
rect 54619 11781 54631 11815
rect 56686 11812 56692 11824
rect 56647 11784 56692 11812
rect 54573 11775 54631 11781
rect 56686 11772 56692 11784
rect 56744 11772 56750 11824
rect 52733 11747 52791 11753
rect 52733 11713 52745 11747
rect 52779 11713 52791 11747
rect 52733 11707 52791 11713
rect 53466 11704 53472 11756
rect 53524 11744 53530 11756
rect 57333 11747 57391 11753
rect 57333 11744 57345 11747
rect 53524 11716 57345 11744
rect 53524 11704 53530 11716
rect 57333 11713 57345 11716
rect 57379 11713 57391 11747
rect 57333 11707 57391 11713
rect 49237 11679 49295 11685
rect 49237 11645 49249 11679
rect 49283 11645 49295 11679
rect 49418 11676 49424 11688
rect 49379 11648 49424 11676
rect 49237 11639 49295 11645
rect 49418 11636 49424 11648
rect 49476 11636 49482 11688
rect 49786 11636 49792 11688
rect 49844 11676 49850 11688
rect 49881 11679 49939 11685
rect 49881 11676 49893 11679
rect 49844 11648 49893 11676
rect 49844 11636 49850 11648
rect 49881 11645 49893 11648
rect 49927 11645 49939 11679
rect 50614 11676 50620 11688
rect 49881 11639 49939 11645
rect 50080 11648 50620 11676
rect 1854 11608 1860 11620
rect 1815 11580 1860 11608
rect 1854 11568 1860 11580
rect 1912 11568 1918 11620
rect 2590 11608 2596 11620
rect 2551 11580 2596 11608
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 2774 11608 2780 11620
rect 2735 11580 2780 11608
rect 2774 11568 2780 11580
rect 2832 11568 2838 11620
rect 49326 11608 49332 11620
rect 49287 11580 49332 11608
rect 49326 11568 49332 11580
rect 49384 11568 49390 11620
rect 49436 11608 49464 11636
rect 50080 11608 50108 11648
rect 50614 11636 50620 11648
rect 50672 11636 50678 11688
rect 51166 11636 51172 11688
rect 51224 11676 51230 11688
rect 51721 11679 51779 11685
rect 51721 11676 51733 11679
rect 51224 11648 51733 11676
rect 51224 11636 51230 11648
rect 51721 11645 51733 11648
rect 51767 11645 51779 11679
rect 51721 11639 51779 11645
rect 52365 11679 52423 11685
rect 52365 11645 52377 11679
rect 52411 11645 52423 11679
rect 52365 11639 52423 11645
rect 52537 11679 52595 11685
rect 52537 11645 52549 11679
rect 52583 11645 52595 11679
rect 52537 11639 52595 11645
rect 52641 11679 52699 11685
rect 52641 11645 52653 11679
rect 52687 11645 52699 11679
rect 52641 11639 52699 11645
rect 49436 11580 50108 11608
rect 50148 11611 50206 11617
rect 50148 11577 50160 11611
rect 50194 11608 50206 11611
rect 51534 11608 51540 11620
rect 50194 11580 51540 11608
rect 50194 11577 50206 11580
rect 50148 11571 50206 11577
rect 51534 11568 51540 11580
rect 51592 11568 51598 11620
rect 52380 11608 52408 11639
rect 52380 11580 52500 11608
rect 52472 11552 52500 11580
rect 52564 11552 52592 11639
rect 52656 11608 52684 11639
rect 52822 11636 52828 11688
rect 52880 11676 52886 11688
rect 52917 11679 52975 11685
rect 52917 11676 52929 11679
rect 52880 11648 52929 11676
rect 52880 11636 52886 11648
rect 52917 11645 52929 11648
rect 52963 11645 52975 11679
rect 54754 11676 54760 11688
rect 54715 11648 54760 11676
rect 52917 11639 52975 11645
rect 54754 11636 54760 11648
rect 54812 11636 54818 11688
rect 54846 11636 54852 11688
rect 54904 11676 54910 11688
rect 55122 11676 55128 11688
rect 54904 11648 54949 11676
rect 55083 11648 55128 11676
rect 54904 11636 54910 11648
rect 55122 11636 55128 11648
rect 55180 11636 55186 11688
rect 55582 11676 55588 11688
rect 55543 11648 55588 11676
rect 55582 11636 55588 11648
rect 55640 11636 55646 11688
rect 55769 11679 55827 11685
rect 55769 11645 55781 11679
rect 55815 11645 55827 11679
rect 55769 11639 55827 11645
rect 54662 11608 54668 11620
rect 52656 11580 54668 11608
rect 54662 11568 54668 11580
rect 54720 11568 54726 11620
rect 55140 11608 55168 11636
rect 55784 11608 55812 11639
rect 56318 11636 56324 11688
rect 56376 11676 56382 11688
rect 56505 11679 56563 11685
rect 56505 11676 56517 11679
rect 56376 11648 56517 11676
rect 56376 11636 56382 11648
rect 56505 11645 56517 11648
rect 56551 11645 56563 11679
rect 57146 11676 57152 11688
rect 57107 11648 57152 11676
rect 56505 11639 56563 11645
rect 57146 11636 57152 11648
rect 57204 11636 57210 11688
rect 55140 11580 55812 11608
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 52454 11500 52460 11552
rect 52512 11500 52518 11552
rect 52546 11500 52552 11552
rect 52604 11500 52610 11552
rect 53006 11500 53012 11552
rect 53064 11540 53070 11552
rect 53101 11543 53159 11549
rect 53101 11540 53113 11543
rect 53064 11512 53113 11540
rect 53064 11500 53070 11512
rect 53101 11509 53113 11512
rect 53147 11509 53159 11543
rect 53101 11503 53159 11509
rect 57793 11543 57851 11549
rect 57793 11509 57805 11543
rect 57839 11540 57851 11543
rect 57974 11540 57980 11552
rect 57839 11512 57980 11540
rect 57839 11509 57851 11512
rect 57793 11503 57851 11509
rect 57974 11500 57980 11512
rect 58032 11500 58038 11552
rect 1104 11450 58880 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 50326 11450
rect 50378 11398 50390 11450
rect 50442 11398 50454 11450
rect 50506 11398 50518 11450
rect 50570 11398 58880 11450
rect 1104 11376 58880 11398
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 50433 11339 50491 11345
rect 50433 11305 50445 11339
rect 50479 11336 50491 11339
rect 50706 11336 50712 11348
rect 50479 11308 50712 11336
rect 50479 11305 50491 11308
rect 50433 11299 50491 11305
rect 50706 11296 50712 11308
rect 50764 11296 50770 11348
rect 51534 11336 51540 11348
rect 51495 11308 51540 11336
rect 51534 11296 51540 11308
rect 51592 11296 51598 11348
rect 52641 11339 52699 11345
rect 52641 11305 52653 11339
rect 52687 11336 52699 11339
rect 52730 11336 52736 11348
rect 52687 11308 52736 11336
rect 52687 11305 52699 11308
rect 52641 11299 52699 11305
rect 52730 11296 52736 11308
rect 52788 11296 52794 11348
rect 53006 11296 53012 11348
rect 53064 11336 53070 11348
rect 56686 11336 56692 11348
rect 53064 11308 54340 11336
rect 53064 11296 53070 11308
rect 4062 11268 4068 11280
rect 1872 11240 4068 11268
rect 1872 11209 1900 11240
rect 4062 11228 4068 11240
rect 4120 11228 4126 11280
rect 52362 11268 52368 11280
rect 49896 11240 52368 11268
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 49896 11209 49924 11240
rect 52362 11228 52368 11240
rect 52420 11228 52426 11280
rect 52546 11228 52552 11280
rect 52604 11268 52610 11280
rect 53650 11268 53656 11280
rect 52604 11240 53656 11268
rect 52604 11228 52610 11240
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 2924 11172 3157 11200
rect 2924 11160 2930 11172
rect 3145 11169 3157 11172
rect 3191 11169 3203 11203
rect 3145 11163 3203 11169
rect 49053 11203 49111 11209
rect 49053 11169 49065 11203
rect 49099 11169 49111 11203
rect 49053 11163 49111 11169
rect 49881 11203 49939 11209
rect 49881 11169 49893 11203
rect 49927 11169 49939 11203
rect 49881 11163 49939 11169
rect 50341 11203 50399 11209
rect 50341 11169 50353 11203
rect 50387 11169 50399 11203
rect 50341 11163 50399 11169
rect 50525 11203 50583 11209
rect 50525 11169 50537 11203
rect 50571 11200 50583 11203
rect 50614 11200 50620 11212
rect 50571 11172 50620 11200
rect 50571 11169 50583 11172
rect 50525 11163 50583 11169
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2056 11064 2084 11095
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2056 11036 2973 11064
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 49068 11064 49096 11163
rect 50356 11132 50384 11163
rect 50614 11160 50620 11172
rect 50672 11160 50678 11212
rect 51442 11200 51448 11212
rect 51403 11172 51448 11200
rect 51442 11160 51448 11172
rect 51500 11160 51506 11212
rect 51629 11203 51687 11209
rect 51629 11169 51641 11203
rect 51675 11200 51687 11203
rect 51994 11200 52000 11212
rect 51675 11172 52000 11200
rect 51675 11169 51687 11172
rect 51629 11163 51687 11169
rect 51994 11160 52000 11172
rect 52052 11160 52058 11212
rect 52822 11160 52828 11212
rect 52880 11209 52886 11212
rect 52880 11203 52933 11209
rect 52880 11169 52887 11203
rect 52921 11169 52933 11203
rect 53006 11200 53012 11212
rect 52967 11172 53012 11200
rect 52880 11163 52933 11169
rect 52880 11160 52886 11163
rect 53006 11160 53012 11172
rect 53064 11160 53070 11212
rect 53116 11209 53144 11240
rect 53650 11228 53656 11240
rect 53708 11228 53714 11280
rect 54202 11268 54208 11280
rect 54036 11240 54208 11268
rect 54036 11209 54064 11240
rect 54202 11228 54208 11240
rect 54260 11228 54266 11280
rect 54312 11209 54340 11308
rect 54496 11308 56692 11336
rect 53101 11203 53159 11209
rect 53101 11169 53113 11203
rect 53147 11169 53159 11203
rect 53101 11163 53159 11169
rect 53377 11203 53435 11209
rect 53377 11169 53389 11203
rect 53423 11200 53435 11203
rect 54021 11203 54079 11209
rect 54021 11200 54033 11203
rect 53423 11172 54033 11200
rect 53423 11169 53435 11172
rect 53377 11163 53435 11169
rect 54021 11169 54033 11172
rect 54067 11169 54079 11203
rect 54021 11163 54079 11169
rect 54113 11203 54171 11209
rect 54113 11169 54125 11203
rect 54159 11169 54171 11203
rect 54113 11163 54171 11169
rect 54297 11203 54355 11209
rect 54297 11169 54309 11203
rect 54343 11169 54355 11203
rect 54297 11163 54355 11169
rect 52638 11132 52644 11144
rect 50356 11104 52644 11132
rect 52638 11092 52644 11104
rect 52696 11092 52702 11144
rect 53190 11132 53196 11144
rect 53151 11104 53196 11132
rect 53190 11092 53196 11104
rect 53248 11132 53254 11144
rect 54128 11132 54156 11163
rect 54496 11132 54524 11308
rect 56686 11296 56692 11308
rect 56744 11296 56750 11348
rect 54662 11268 54668 11280
rect 54623 11240 54668 11268
rect 54662 11228 54668 11240
rect 54720 11228 54726 11280
rect 55582 11228 55588 11280
rect 55640 11268 55646 11280
rect 57974 11268 57980 11280
rect 55640 11240 56732 11268
rect 57935 11240 57980 11268
rect 55640 11228 55646 11240
rect 54570 11160 54576 11212
rect 54628 11200 54634 11212
rect 55309 11203 55367 11209
rect 54628 11172 54673 11200
rect 54628 11160 54634 11172
rect 55309 11169 55321 11203
rect 55355 11169 55367 11203
rect 55490 11200 55496 11212
rect 55451 11172 55496 11200
rect 55309 11163 55367 11169
rect 53248 11104 54156 11132
rect 54312 11104 54524 11132
rect 55324 11132 55352 11163
rect 55490 11160 55496 11172
rect 55548 11160 55554 11212
rect 55674 11200 55680 11212
rect 55635 11172 55680 11200
rect 55674 11160 55680 11172
rect 55732 11160 55738 11212
rect 56704 11209 56732 11240
rect 57974 11228 57980 11240
rect 58032 11228 58038 11280
rect 58158 11268 58164 11280
rect 58119 11240 58164 11268
rect 58158 11228 58164 11240
rect 58216 11228 58222 11280
rect 56689 11203 56747 11209
rect 56689 11169 56701 11203
rect 56735 11169 56747 11203
rect 56689 11163 56747 11169
rect 56873 11203 56931 11209
rect 56873 11169 56885 11203
rect 56919 11169 56931 11203
rect 56873 11163 56931 11169
rect 55582 11132 55588 11144
rect 55324 11104 55588 11132
rect 53248 11092 53254 11104
rect 49068 11036 51074 11064
rect 2961 11027 3019 11033
rect 51046 10996 51074 11036
rect 52086 11024 52092 11076
rect 52144 11064 52150 11076
rect 54312 11064 54340 11104
rect 55582 11092 55588 11104
rect 55640 11092 55646 11144
rect 55766 11092 55772 11144
rect 55824 11132 55830 11144
rect 56888 11132 56916 11163
rect 55824 11104 56916 11132
rect 55824 11092 55830 11104
rect 52144 11036 54340 11064
rect 52144 11024 52150 11036
rect 54662 11024 54668 11076
rect 54720 11064 54726 11076
rect 55309 11067 55367 11073
rect 55309 11064 55321 11067
rect 54720 11036 55321 11064
rect 54720 11024 54726 11036
rect 55309 11033 55321 11036
rect 55355 11033 55367 11067
rect 55309 11027 55367 11033
rect 55214 10996 55220 11008
rect 51046 10968 55220 10996
rect 55214 10956 55220 10968
rect 55272 10956 55278 11008
rect 56686 10996 56692 11008
rect 56647 10968 56692 10996
rect 56686 10956 56692 10968
rect 56744 10956 56750 11008
rect 1104 10906 58880 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 58880 10906
rect 1104 10832 58880 10854
rect 1854 10752 1860 10804
rect 1912 10792 1918 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1912 10764 2053 10792
rect 1912 10752 1918 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 54018 10752 54024 10804
rect 54076 10792 54082 10804
rect 54938 10792 54944 10804
rect 54076 10764 54944 10792
rect 54076 10752 54082 10764
rect 54938 10752 54944 10764
rect 54996 10752 55002 10804
rect 55033 10795 55091 10801
rect 55033 10761 55045 10795
rect 55079 10792 55091 10795
rect 55674 10792 55680 10804
rect 55079 10764 55680 10792
rect 55079 10761 55091 10764
rect 55033 10755 55091 10761
rect 55674 10752 55680 10764
rect 55732 10752 55738 10804
rect 52181 10727 52239 10733
rect 52181 10693 52193 10727
rect 52227 10724 52239 10727
rect 53098 10724 53104 10736
rect 52227 10696 53104 10724
rect 52227 10693 52239 10696
rect 52181 10687 52239 10693
rect 53098 10684 53104 10696
rect 53156 10724 53162 10736
rect 53834 10724 53840 10736
rect 53156 10696 53840 10724
rect 53156 10684 53162 10696
rect 53834 10684 53840 10696
rect 53892 10684 53898 10736
rect 54294 10684 54300 10736
rect 54352 10724 54358 10736
rect 54352 10696 55536 10724
rect 54352 10684 54358 10696
rect 50157 10659 50215 10665
rect 50157 10625 50169 10659
rect 50203 10656 50215 10659
rect 54386 10656 54392 10668
rect 50203 10628 54392 10656
rect 50203 10625 50215 10628
rect 50157 10619 50215 10625
rect 54386 10616 54392 10628
rect 54444 10616 54450 10668
rect 54754 10656 54760 10668
rect 54496 10628 54760 10656
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 2498 10588 2504 10600
rect 1903 10560 2504 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 1688 10520 1716 10551
rect 2498 10548 2504 10560
rect 2556 10548 2562 10600
rect 50798 10588 50804 10600
rect 50759 10560 50804 10588
rect 50798 10548 50804 10560
rect 50856 10548 50862 10600
rect 51445 10591 51503 10597
rect 51445 10557 51457 10591
rect 51491 10588 51503 10591
rect 51902 10588 51908 10600
rect 51491 10560 51908 10588
rect 51491 10557 51503 10560
rect 51445 10551 51503 10557
rect 51902 10548 51908 10560
rect 51960 10548 51966 10600
rect 51997 10591 52055 10597
rect 51997 10557 52009 10591
rect 52043 10588 52055 10591
rect 52086 10588 52092 10600
rect 52043 10560 52092 10588
rect 52043 10557 52055 10560
rect 51997 10551 52055 10557
rect 52086 10548 52092 10560
rect 52144 10548 52150 10600
rect 54496 10597 54524 10628
rect 54754 10616 54760 10628
rect 54812 10616 54818 10668
rect 55508 10656 55536 10696
rect 55508 10628 55628 10656
rect 52917 10591 52975 10597
rect 52917 10557 52929 10591
rect 52963 10557 52975 10591
rect 52917 10551 52975 10557
rect 54481 10591 54539 10597
rect 54481 10557 54493 10591
rect 54527 10557 54539 10591
rect 54481 10551 54539 10557
rect 54849 10591 54907 10597
rect 54849 10557 54861 10591
rect 54895 10557 54907 10591
rect 54849 10551 54907 10557
rect 3326 10520 3332 10532
rect 1688 10492 3332 10520
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 52932 10520 52960 10551
rect 54662 10520 54668 10532
rect 52932 10492 54524 10520
rect 54623 10492 54668 10520
rect 54496 10464 54524 10492
rect 54662 10480 54668 10492
rect 54720 10480 54726 10532
rect 54757 10523 54815 10529
rect 54757 10489 54769 10523
rect 54803 10489 54815 10523
rect 54757 10483 54815 10489
rect 51258 10452 51264 10464
rect 51219 10424 51264 10452
rect 51258 10412 51264 10424
rect 51316 10412 51322 10464
rect 52914 10412 52920 10464
rect 52972 10452 52978 10464
rect 53009 10455 53067 10461
rect 53009 10452 53021 10455
rect 52972 10424 53021 10452
rect 52972 10412 52978 10424
rect 53009 10421 53021 10424
rect 53055 10452 53067 10455
rect 53190 10452 53196 10464
rect 53055 10424 53196 10452
rect 53055 10421 53067 10424
rect 53009 10415 53067 10421
rect 53190 10412 53196 10424
rect 53248 10412 53254 10464
rect 54478 10412 54484 10464
rect 54536 10412 54542 10464
rect 54570 10412 54576 10464
rect 54628 10452 54634 10464
rect 54772 10452 54800 10483
rect 54628 10424 54800 10452
rect 54864 10452 54892 10551
rect 54938 10548 54944 10600
rect 54996 10588 55002 10600
rect 55493 10591 55551 10597
rect 55493 10588 55505 10591
rect 54996 10560 55505 10588
rect 54996 10548 55002 10560
rect 55493 10557 55505 10560
rect 55539 10557 55551 10591
rect 55600 10588 55628 10628
rect 55760 10591 55818 10597
rect 55600 10560 55720 10588
rect 55493 10551 55551 10557
rect 55692 10520 55720 10560
rect 55760 10557 55772 10591
rect 55806 10588 55818 10591
rect 56686 10588 56692 10600
rect 55806 10560 56692 10588
rect 55806 10557 55818 10560
rect 55760 10551 55818 10557
rect 56686 10548 56692 10560
rect 56744 10548 56750 10600
rect 57514 10520 57520 10532
rect 55692 10492 57520 10520
rect 57514 10480 57520 10492
rect 57572 10480 57578 10532
rect 57974 10520 57980 10532
rect 57935 10492 57980 10520
rect 57974 10480 57980 10492
rect 58032 10480 58038 10532
rect 58158 10520 58164 10532
rect 58119 10492 58164 10520
rect 58158 10480 58164 10492
rect 58216 10480 58222 10532
rect 55674 10452 55680 10464
rect 54864 10424 55680 10452
rect 54628 10412 54634 10424
rect 55674 10412 55680 10424
rect 55732 10452 55738 10464
rect 56873 10455 56931 10461
rect 56873 10452 56885 10455
rect 55732 10424 56885 10452
rect 55732 10412 55738 10424
rect 56873 10421 56885 10424
rect 56919 10421 56931 10455
rect 56873 10415 56931 10421
rect 1104 10362 58880 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 50326 10362
rect 50378 10310 50390 10362
rect 50442 10310 50454 10362
rect 50506 10310 50518 10362
rect 50570 10310 58880 10362
rect 1104 10288 58880 10310
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 50798 10208 50804 10260
rect 50856 10248 50862 10260
rect 54294 10248 54300 10260
rect 50856 10220 54300 10248
rect 50856 10208 50862 10220
rect 54294 10208 54300 10220
rect 54352 10208 54358 10260
rect 54386 10208 54392 10260
rect 54444 10248 54450 10260
rect 56689 10251 56747 10257
rect 56689 10248 56701 10251
rect 54444 10220 56701 10248
rect 54444 10208 54450 10220
rect 56689 10217 56701 10220
rect 56735 10217 56747 10251
rect 56689 10211 56747 10217
rect 57974 10208 57980 10260
rect 58032 10248 58038 10260
rect 58161 10251 58219 10257
rect 58161 10248 58173 10251
rect 58032 10220 58173 10248
rect 58032 10208 58038 10220
rect 58161 10217 58173 10220
rect 58207 10217 58219 10251
rect 58161 10211 58219 10217
rect 50062 10140 50068 10192
rect 50120 10180 50126 10192
rect 50157 10183 50215 10189
rect 50157 10180 50169 10183
rect 50120 10152 50169 10180
rect 50120 10140 50126 10152
rect 50157 10149 50169 10152
rect 50203 10149 50215 10183
rect 50157 10143 50215 10149
rect 51258 10140 51264 10192
rect 51316 10180 51322 10192
rect 51316 10152 57744 10180
rect 51316 10140 51322 10152
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 2866 10112 2872 10124
rect 2731 10084 2872 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3326 10112 3332 10124
rect 3287 10084 3332 10112
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 49329 10115 49387 10121
rect 49329 10081 49341 10115
rect 49375 10081 49387 10115
rect 49970 10112 49976 10124
rect 49931 10084 49976 10112
rect 49329 10075 49387 10081
rect 49344 10044 49372 10075
rect 49970 10072 49976 10084
rect 50028 10072 50034 10124
rect 51166 10072 51172 10124
rect 51224 10112 51230 10124
rect 51701 10115 51759 10121
rect 51701 10112 51713 10115
rect 51224 10084 51713 10112
rect 51224 10072 51230 10084
rect 51701 10081 51713 10084
rect 51747 10081 51759 10115
rect 51701 10075 51759 10081
rect 52454 10072 52460 10124
rect 52512 10112 52518 10124
rect 53515 10115 53573 10121
rect 53515 10112 53527 10115
rect 52512 10084 53527 10112
rect 52512 10072 52518 10084
rect 53515 10081 53527 10084
rect 53561 10081 53573 10115
rect 53515 10075 53573 10081
rect 53653 10115 53711 10121
rect 53653 10081 53665 10115
rect 53699 10081 53711 10115
rect 53653 10075 53711 10081
rect 53745 10115 53803 10121
rect 53745 10081 53757 10115
rect 53791 10112 53803 10115
rect 53834 10112 53840 10124
rect 53791 10084 53840 10112
rect 53791 10081 53803 10084
rect 53745 10075 53803 10081
rect 50154 10044 50160 10056
rect 49344 10016 50160 10044
rect 50154 10004 50160 10016
rect 50212 10004 50218 10056
rect 50982 10004 50988 10056
rect 51040 10044 51046 10056
rect 51445 10047 51503 10053
rect 51445 10044 51457 10047
rect 51040 10016 51457 10044
rect 51040 10004 51046 10016
rect 51445 10013 51457 10016
rect 51491 10013 51503 10047
rect 53668 10044 53696 10075
rect 53834 10072 53840 10084
rect 53892 10072 53898 10124
rect 53926 10072 53932 10124
rect 53984 10112 53990 10124
rect 54570 10112 54576 10124
rect 53984 10084 54029 10112
rect 54483 10084 54576 10112
rect 53984 10072 53990 10084
rect 54570 10072 54576 10084
rect 54628 10072 54634 10124
rect 55214 10112 55220 10124
rect 55175 10084 55220 10112
rect 55214 10072 55220 10084
rect 55272 10072 55278 10124
rect 55355 10115 55413 10121
rect 55355 10081 55367 10115
rect 55401 10081 55413 10115
rect 55355 10075 55413 10081
rect 54478 10044 54484 10056
rect 53668 10016 54484 10044
rect 51445 10007 51503 10013
rect 54478 10004 54484 10016
rect 54536 10004 54542 10056
rect 52825 9979 52883 9985
rect 52825 9945 52837 9979
rect 52871 9976 52883 9979
rect 54588 9976 54616 10072
rect 54665 10047 54723 10053
rect 54665 10013 54677 10047
rect 54711 10044 54723 10047
rect 55385 10044 55413 10075
rect 55490 10072 55496 10124
rect 55548 10112 55554 10124
rect 55674 10121 55680 10124
rect 55631 10115 55680 10121
rect 55548 10084 55593 10112
rect 55548 10072 55554 10084
rect 55631 10081 55643 10115
rect 55677 10081 55680 10115
rect 55631 10075 55680 10081
rect 55674 10072 55680 10075
rect 55732 10072 55738 10124
rect 56870 10112 56876 10124
rect 56831 10084 56876 10112
rect 56870 10072 56876 10084
rect 56928 10072 56934 10124
rect 57716 10121 57744 10152
rect 57701 10115 57759 10121
rect 57701 10081 57713 10115
rect 57747 10081 57759 10115
rect 57701 10075 57759 10081
rect 55766 10044 55772 10056
rect 54711 10016 55772 10044
rect 54711 10013 54723 10016
rect 54665 10007 54723 10013
rect 55766 10004 55772 10016
rect 55824 10004 55830 10056
rect 56689 10047 56747 10053
rect 56689 10013 56701 10047
rect 56735 10044 56747 10047
rect 57517 10047 57575 10053
rect 57517 10044 57529 10047
rect 56735 10016 57529 10044
rect 56735 10013 56747 10016
rect 56689 10007 56747 10013
rect 57517 10013 57529 10016
rect 57563 10013 57575 10047
rect 57517 10007 57575 10013
rect 55490 9976 55496 9988
rect 52871 9948 55496 9976
rect 52871 9945 52883 9948
rect 52825 9939 52883 9945
rect 55490 9936 55496 9948
rect 55548 9936 55554 9988
rect 57054 9976 57060 9988
rect 57015 9948 57060 9976
rect 57054 9936 57060 9948
rect 57112 9936 57118 9988
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 50338 9908 50344 9920
rect 50299 9880 50344 9908
rect 50338 9868 50344 9880
rect 50396 9868 50402 9920
rect 53285 9911 53343 9917
rect 53285 9877 53297 9911
rect 53331 9908 53343 9911
rect 54110 9908 54116 9920
rect 53331 9880 54116 9908
rect 53331 9877 53343 9880
rect 53285 9871 53343 9877
rect 54110 9868 54116 9880
rect 54168 9868 54174 9920
rect 54202 9868 54208 9920
rect 54260 9908 54266 9920
rect 55769 9911 55827 9917
rect 55769 9908 55781 9911
rect 54260 9880 55781 9908
rect 54260 9868 54266 9880
rect 55769 9877 55781 9880
rect 55815 9877 55827 9911
rect 55769 9871 55827 9877
rect 1104 9818 58880 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 58880 9818
rect 1104 9744 58880 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 2133 9707 2191 9713
rect 2133 9704 2145 9707
rect 1912 9676 2145 9704
rect 1912 9664 1918 9676
rect 2133 9673 2145 9676
rect 2179 9673 2191 9707
rect 51166 9704 51172 9716
rect 51127 9676 51172 9704
rect 2133 9667 2191 9673
rect 51166 9664 51172 9676
rect 51224 9664 51230 9716
rect 54036 9676 54984 9704
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 1964 9608 2881 9636
rect 1964 9577 1992 9608
rect 2869 9605 2881 9608
rect 2915 9605 2927 9639
rect 2869 9599 2927 9605
rect 50706 9596 50712 9648
rect 50764 9636 50770 9648
rect 54036 9636 54064 9676
rect 50764 9608 54064 9636
rect 54956 9636 54984 9676
rect 56870 9664 56876 9716
rect 56928 9704 56934 9716
rect 57149 9707 57207 9713
rect 57149 9704 57161 9707
rect 56928 9676 57161 9704
rect 56928 9664 56934 9676
rect 57149 9673 57161 9676
rect 57195 9673 57207 9707
rect 57149 9667 57207 9673
rect 54956 9608 56824 9636
rect 50764 9596 50770 9608
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 3697 9571 3755 9577
rect 3697 9568 3709 9571
rect 1949 9531 2007 9537
rect 2700 9540 3709 9568
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2700 9500 2728 9540
rect 3697 9537 3709 9540
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 50154 9528 50160 9580
rect 50212 9568 50218 9580
rect 56796 9577 56824 9608
rect 56781 9571 56839 9577
rect 50212 9540 52040 9568
rect 50212 9528 50218 9540
rect 1811 9472 2728 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2866 9460 2872 9512
rect 2924 9500 2930 9512
rect 3053 9503 3111 9509
rect 3053 9500 3065 9503
rect 2924 9472 3065 9500
rect 2924 9460 2930 9472
rect 3053 9469 3065 9472
rect 3099 9469 3111 9503
rect 3053 9463 3111 9469
rect 49053 9503 49111 9509
rect 49053 9469 49065 9503
rect 49099 9469 49111 9503
rect 49053 9463 49111 9469
rect 49320 9503 49378 9509
rect 49320 9469 49332 9503
rect 49366 9500 49378 9503
rect 50338 9500 50344 9512
rect 49366 9472 50344 9500
rect 49366 9469 49378 9472
rect 49320 9463 49378 9469
rect 48866 9392 48872 9444
rect 48924 9432 48930 9444
rect 49068 9432 49096 9463
rect 50338 9460 50344 9472
rect 50396 9460 50402 9512
rect 51169 9503 51227 9509
rect 51169 9469 51181 9503
rect 51215 9469 51227 9503
rect 51350 9500 51356 9512
rect 51311 9472 51356 9500
rect 51169 9463 51227 9469
rect 50982 9432 50988 9444
rect 48924 9404 50988 9432
rect 48924 9392 48930 9404
rect 50982 9392 50988 9404
rect 51040 9392 51046 9444
rect 51184 9432 51212 9463
rect 51350 9460 51356 9472
rect 51408 9500 51414 9512
rect 51810 9500 51816 9512
rect 51408 9472 51816 9500
rect 51408 9460 51414 9472
rect 51810 9460 51816 9472
rect 51868 9460 51874 9512
rect 52012 9432 52040 9540
rect 52288 9540 52592 9568
rect 52086 9503 52144 9509
rect 52086 9469 52098 9503
rect 52132 9500 52144 9503
rect 52288 9500 52316 9540
rect 52454 9500 52460 9512
rect 52132 9472 52316 9500
rect 52415 9472 52460 9500
rect 52132 9469 52144 9472
rect 52086 9463 52144 9469
rect 52454 9460 52460 9472
rect 52512 9460 52518 9512
rect 52564 9509 52592 9540
rect 56781 9537 56793 9571
rect 56827 9537 56839 9571
rect 56781 9531 56839 9537
rect 52549 9503 52607 9509
rect 52549 9469 52561 9503
rect 52595 9500 52607 9503
rect 53377 9503 53435 9509
rect 53377 9500 53389 9503
rect 52595 9472 53389 9500
rect 52595 9469 52607 9472
rect 52549 9463 52607 9469
rect 53377 9469 53389 9472
rect 53423 9469 53435 9503
rect 53377 9463 53435 9469
rect 53834 9460 53840 9512
rect 53892 9500 53898 9512
rect 54018 9500 54024 9512
rect 53892 9472 54024 9500
rect 53892 9460 53898 9472
rect 54018 9460 54024 9472
rect 54076 9460 54082 9512
rect 54110 9460 54116 9512
rect 54168 9500 54174 9512
rect 54277 9503 54335 9509
rect 54277 9500 54289 9503
rect 54168 9472 54289 9500
rect 54168 9460 54174 9472
rect 54277 9469 54289 9472
rect 54323 9469 54335 9503
rect 54277 9463 54335 9469
rect 55582 9460 55588 9512
rect 55640 9500 55646 9512
rect 55861 9503 55919 9509
rect 55861 9500 55873 9503
rect 55640 9472 55873 9500
rect 55640 9460 55646 9472
rect 55861 9469 55873 9472
rect 55907 9469 55919 9503
rect 56962 9500 56968 9512
rect 56923 9472 56968 9500
rect 55861 9463 55919 9469
rect 56962 9460 56968 9472
rect 57020 9460 57026 9512
rect 55214 9432 55220 9444
rect 51184 9404 51948 9432
rect 52012 9404 55220 9432
rect 50154 9324 50160 9376
rect 50212 9364 50218 9376
rect 51920 9373 51948 9404
rect 55214 9392 55220 9404
rect 55272 9392 55278 9444
rect 55306 9392 55312 9444
rect 55364 9432 55370 9444
rect 57974 9432 57980 9444
rect 55364 9404 55996 9432
rect 57935 9404 57980 9432
rect 55364 9392 55370 9404
rect 55968 9376 55996 9404
rect 57974 9392 57980 9404
rect 58032 9392 58038 9444
rect 58158 9432 58164 9444
rect 58119 9404 58164 9432
rect 58158 9392 58164 9404
rect 58216 9392 58222 9444
rect 50433 9367 50491 9373
rect 50433 9364 50445 9367
rect 50212 9336 50445 9364
rect 50212 9324 50218 9336
rect 50433 9333 50445 9336
rect 50479 9333 50491 9367
rect 50433 9327 50491 9333
rect 51905 9367 51963 9373
rect 51905 9333 51917 9367
rect 51951 9333 51963 9367
rect 51905 9327 51963 9333
rect 52089 9367 52147 9373
rect 52089 9333 52101 9367
rect 52135 9364 52147 9367
rect 52454 9364 52460 9376
rect 52135 9336 52460 9364
rect 52135 9333 52147 9336
rect 52089 9327 52147 9333
rect 52454 9324 52460 9336
rect 52512 9324 52518 9376
rect 53377 9367 53435 9373
rect 53377 9333 53389 9367
rect 53423 9364 53435 9367
rect 54202 9364 54208 9376
rect 53423 9336 54208 9364
rect 53423 9333 53435 9336
rect 53377 9327 53435 9333
rect 54202 9324 54208 9336
rect 54260 9324 54266 9376
rect 54662 9324 54668 9376
rect 54720 9364 54726 9376
rect 55401 9367 55459 9373
rect 55401 9364 55413 9367
rect 54720 9336 55413 9364
rect 54720 9324 54726 9336
rect 55401 9333 55413 9336
rect 55447 9333 55459 9367
rect 55950 9364 55956 9376
rect 55911 9336 55956 9364
rect 55401 9327 55459 9333
rect 55950 9324 55956 9336
rect 56008 9324 56014 9376
rect 1104 9274 58880 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 50326 9274
rect 50378 9222 50390 9274
rect 50442 9222 50454 9274
rect 50506 9222 50518 9274
rect 50570 9222 58880 9274
rect 1104 9200 58880 9222
rect 49970 9160 49976 9172
rect 49931 9132 49976 9160
rect 49970 9120 49976 9132
rect 50028 9120 50034 9172
rect 50706 9120 50712 9172
rect 50764 9160 50770 9172
rect 51994 9160 52000 9172
rect 50764 9132 52000 9160
rect 50764 9120 50770 9132
rect 51994 9120 52000 9132
rect 52052 9120 52058 9172
rect 52365 9163 52423 9169
rect 52365 9129 52377 9163
rect 52411 9160 52423 9163
rect 53285 9163 53343 9169
rect 52411 9132 53052 9160
rect 52411 9129 52423 9132
rect 52365 9123 52423 9129
rect 53024 9104 53052 9132
rect 53285 9129 53297 9163
rect 53331 9160 53343 9163
rect 53926 9160 53932 9172
rect 53331 9132 53932 9160
rect 53331 9129 53343 9132
rect 53285 9123 53343 9129
rect 53926 9120 53932 9132
rect 53984 9120 53990 9172
rect 54478 9160 54484 9172
rect 54439 9132 54484 9160
rect 54478 9120 54484 9132
rect 54536 9120 54542 9172
rect 56873 9163 56931 9169
rect 56873 9129 56885 9163
rect 56919 9160 56931 9163
rect 57698 9160 57704 9172
rect 56919 9132 57704 9160
rect 56919 9129 56931 9132
rect 56873 9123 56931 9129
rect 57698 9120 57704 9132
rect 57756 9120 57762 9172
rect 57974 9120 57980 9172
rect 58032 9160 58038 9172
rect 58161 9163 58219 9169
rect 58161 9160 58173 9163
rect 58032 9132 58173 9160
rect 58032 9120 58038 9132
rect 58161 9129 58173 9132
rect 58207 9129 58219 9163
rect 58161 9123 58219 9129
rect 50890 9092 50896 9104
rect 48700 9064 50896 9092
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 2961 9027 3019 9033
rect 2961 9024 2973 9027
rect 2924 8996 2973 9024
rect 2924 8984 2930 8996
rect 2961 8993 2973 8996
rect 3007 8993 3019 9027
rect 48038 9024 48044 9036
rect 47999 8996 48044 9024
rect 2961 8987 3019 8993
rect 48038 8984 48044 8996
rect 48096 8984 48102 9036
rect 48700 9033 48728 9064
rect 50890 9052 50896 9064
rect 50948 9052 50954 9104
rect 51537 9095 51595 9101
rect 51537 9061 51549 9095
rect 51583 9092 51595 9095
rect 51626 9092 51632 9104
rect 51583 9064 51632 9092
rect 51583 9061 51595 9064
rect 51537 9055 51595 9061
rect 51626 9052 51632 9064
rect 51684 9052 51690 9104
rect 52914 9092 52920 9104
rect 52875 9064 52920 9092
rect 52914 9052 52920 9064
rect 52972 9052 52978 9104
rect 53006 9052 53012 9104
rect 53064 9092 53070 9104
rect 53101 9095 53159 9101
rect 53101 9092 53113 9095
rect 53064 9064 53113 9092
rect 53064 9052 53070 9064
rect 53101 9061 53113 9064
rect 53147 9061 53159 9095
rect 54386 9092 54392 9104
rect 53101 9055 53159 9061
rect 53760 9064 54392 9092
rect 48685 9027 48743 9033
rect 48685 8993 48697 9027
rect 48731 8993 48743 9027
rect 48685 8987 48743 8993
rect 48869 9027 48927 9033
rect 48869 8993 48881 9027
rect 48915 8993 48927 9027
rect 49510 9024 49516 9036
rect 49471 8996 49516 9024
rect 48869 8987 48927 8993
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 1857 8959 1915 8965
rect 1857 8925 1869 8959
rect 1903 8925 1915 8959
rect 48884 8956 48912 8987
rect 49510 8984 49516 8996
rect 49568 8984 49574 9036
rect 50154 9024 50160 9036
rect 50115 8996 50160 9024
rect 50154 8984 50160 8996
rect 50212 8984 50218 9036
rect 50246 8984 50252 9036
rect 50304 9024 50310 9036
rect 50525 9027 50583 9033
rect 50304 8996 50349 9024
rect 50304 8984 50310 8996
rect 50525 8993 50537 9027
rect 50571 9024 50583 9027
rect 50798 9024 50804 9036
rect 50571 8996 50804 9024
rect 50571 8993 50583 8996
rect 50525 8987 50583 8993
rect 50798 8984 50804 8996
rect 50856 8984 50862 9036
rect 52273 9027 52331 9033
rect 51644 8996 51856 9024
rect 49602 8956 49608 8968
rect 48884 8928 49608 8956
rect 1857 8919 1915 8925
rect 1872 8888 1900 8919
rect 49602 8916 49608 8928
rect 49660 8956 49666 8968
rect 50433 8959 50491 8965
rect 50433 8956 50445 8959
rect 49660 8928 50445 8956
rect 49660 8916 49666 8928
rect 50433 8925 50445 8928
rect 50479 8956 50491 8959
rect 51442 8956 51448 8968
rect 50479 8928 51448 8956
rect 50479 8925 50491 8928
rect 50433 8919 50491 8925
rect 51442 8916 51448 8928
rect 51500 8916 51506 8968
rect 2777 8891 2835 8897
rect 2777 8888 2789 8891
rect 1872 8860 2789 8888
rect 2777 8857 2789 8860
rect 2823 8857 2835 8891
rect 2777 8851 2835 8857
rect 49329 8891 49387 8897
rect 49329 8857 49341 8891
rect 49375 8888 49387 8891
rect 51644 8888 51672 8996
rect 49375 8860 51672 8888
rect 51828 8888 51856 8996
rect 52273 8993 52285 9027
rect 52319 9024 52331 9027
rect 52362 9024 52368 9036
rect 52319 8996 52368 9024
rect 52319 8993 52331 8996
rect 52273 8987 52331 8993
rect 52362 8984 52368 8996
rect 52420 8984 52426 9036
rect 53760 9033 53788 9064
rect 54386 9052 54392 9064
rect 54444 9052 54450 9104
rect 54680 9064 55536 9092
rect 54680 9036 54708 9064
rect 53745 9027 53803 9033
rect 53745 9024 53757 9027
rect 52472 8996 53757 9024
rect 52181 8959 52239 8965
rect 52181 8925 52193 8959
rect 52227 8956 52239 8959
rect 52472 8956 52500 8996
rect 53745 8993 53757 8996
rect 53791 8993 53803 9027
rect 53745 8987 53803 8993
rect 53929 9027 53987 9033
rect 53929 8993 53941 9027
rect 53975 8993 53987 9027
rect 54662 9024 54668 9036
rect 54623 8996 54668 9024
rect 53929 8987 53987 8993
rect 52227 8928 52500 8956
rect 52227 8925 52239 8928
rect 52181 8919 52239 8925
rect 52822 8916 52828 8968
rect 52880 8956 52886 8968
rect 53944 8956 53972 8987
rect 54662 8984 54668 8996
rect 54720 8984 54726 9036
rect 54754 8984 54760 9036
rect 54812 9024 54818 9036
rect 55508 9033 55536 9064
rect 55033 9027 55091 9033
rect 54812 8996 54857 9024
rect 54812 8984 54818 8996
rect 55033 8993 55045 9027
rect 55079 8993 55091 9027
rect 55033 8987 55091 8993
rect 55493 9027 55551 9033
rect 55493 8993 55505 9027
rect 55539 8993 55551 9027
rect 55493 8987 55551 8993
rect 55048 8956 55076 8987
rect 56778 8984 56784 9036
rect 56836 9024 56842 9036
rect 57057 9027 57115 9033
rect 57057 9024 57069 9027
rect 56836 8996 57069 9024
rect 56836 8984 56842 8996
rect 57057 8993 57069 8996
rect 57103 8993 57115 9027
rect 57514 9024 57520 9036
rect 57475 8996 57520 9024
rect 57057 8987 57115 8993
rect 57514 8984 57520 8996
rect 57572 8984 57578 9036
rect 55585 8959 55643 8965
rect 55585 8956 55597 8959
rect 52880 8928 55597 8956
rect 52880 8916 52886 8928
rect 55585 8925 55597 8928
rect 55631 8925 55643 8959
rect 57698 8956 57704 8968
rect 57659 8928 57704 8956
rect 55585 8919 55643 8925
rect 57698 8916 57704 8928
rect 57756 8916 57762 8968
rect 56962 8888 56968 8900
rect 51828 8860 56968 8888
rect 49375 8857 49387 8860
rect 49329 8851 49387 8857
rect 56962 8848 56968 8860
rect 57020 8848 57026 8900
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 2590 8820 2596 8832
rect 2363 8792 2596 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 48682 8820 48688 8832
rect 48643 8792 48688 8820
rect 48682 8780 48688 8792
rect 48740 8780 48746 8832
rect 49878 8780 49884 8832
rect 49936 8820 49942 8832
rect 51629 8823 51687 8829
rect 51629 8820 51641 8823
rect 49936 8792 51641 8820
rect 49936 8780 49942 8792
rect 51629 8789 51641 8792
rect 51675 8820 51687 8823
rect 52181 8823 52239 8829
rect 52181 8820 52193 8823
rect 51675 8792 52193 8820
rect 51675 8789 51687 8792
rect 51629 8783 51687 8789
rect 52181 8789 52193 8792
rect 52227 8789 52239 8823
rect 52181 8783 52239 8789
rect 53745 8823 53803 8829
rect 53745 8789 53757 8823
rect 53791 8820 53803 8823
rect 54110 8820 54116 8832
rect 53791 8792 54116 8820
rect 53791 8789 53803 8792
rect 53745 8783 53803 8789
rect 54110 8780 54116 8792
rect 54168 8780 54174 8832
rect 54938 8820 54944 8832
rect 54899 8792 54944 8820
rect 54938 8780 54944 8792
rect 54996 8780 55002 8832
rect 1104 8730 58880 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 58880 8730
rect 1104 8656 58880 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 1728 8588 4353 8616
rect 1728 8576 1734 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 4341 8579 4399 8585
rect 47673 8619 47731 8625
rect 47673 8585 47685 8619
rect 47719 8616 47731 8619
rect 47719 8588 56456 8616
rect 47719 8585 47731 8588
rect 47673 8579 47731 8585
rect 2774 8548 2780 8560
rect 2735 8520 2780 8548
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 3694 8548 3700 8560
rect 3651 8520 3700 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 3694 8508 3700 8520
rect 3752 8508 3758 8560
rect 50246 8548 50252 8560
rect 50159 8520 50252 8548
rect 50246 8508 50252 8520
rect 50304 8548 50310 8560
rect 51442 8548 51448 8560
rect 50304 8520 51074 8548
rect 51403 8520 51448 8548
rect 50304 8508 50310 8520
rect 48866 8480 48872 8492
rect 3344 8452 26234 8480
rect 48827 8452 48872 8480
rect 2590 8412 2596 8424
rect 2551 8384 2596 8412
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 3142 8412 3148 8424
rect 3055 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8412 3206 8424
rect 3344 8421 3372 8452
rect 3329 8415 3387 8421
rect 3329 8412 3341 8415
rect 3200 8384 3341 8412
rect 3200 8372 3206 8384
rect 3329 8381 3341 8384
rect 3375 8381 3387 8415
rect 3329 8375 3387 8381
rect 1854 8344 1860 8356
rect 1815 8316 1860 8344
rect 1854 8304 1860 8316
rect 1912 8304 1918 8356
rect 2038 8344 2044 8356
rect 1999 8316 2044 8344
rect 2038 8304 2044 8316
rect 2096 8304 2102 8356
rect 26206 8344 26234 8452
rect 48866 8440 48872 8452
rect 48924 8440 48930 8492
rect 50154 8440 50160 8492
rect 50212 8480 50218 8492
rect 51046 8480 51074 8520
rect 51442 8508 51448 8520
rect 51500 8508 51506 8560
rect 51736 8520 52408 8548
rect 50212 8452 50752 8480
rect 51046 8452 51396 8480
rect 50212 8440 50218 8452
rect 47026 8412 47032 8424
rect 46987 8384 47032 8412
rect 47026 8372 47032 8384
rect 47084 8372 47090 8424
rect 47673 8415 47731 8421
rect 47673 8381 47685 8415
rect 47719 8381 47731 8415
rect 47673 8375 47731 8381
rect 47578 8344 47584 8356
rect 26206 8316 47584 8344
rect 47578 8304 47584 8316
rect 47636 8304 47642 8356
rect 47688 8344 47716 8375
rect 47762 8372 47768 8424
rect 47820 8412 47826 8424
rect 50724 8421 50752 8452
rect 51368 8421 51396 8452
rect 47857 8415 47915 8421
rect 47857 8412 47869 8415
rect 47820 8384 47869 8412
rect 47820 8372 47826 8384
rect 47857 8381 47869 8384
rect 47903 8381 47915 8415
rect 50709 8415 50767 8421
rect 47857 8375 47915 8381
rect 49068 8384 50200 8412
rect 49068 8344 49096 8384
rect 47688 8316 49096 8344
rect 49136 8347 49194 8353
rect 49136 8313 49148 8347
rect 49182 8344 49194 8347
rect 50062 8344 50068 8356
rect 49182 8316 50068 8344
rect 49182 8313 49194 8316
rect 49136 8307 49194 8313
rect 50062 8304 50068 8316
rect 50120 8304 50126 8356
rect 50172 8344 50200 8384
rect 50709 8381 50721 8415
rect 50755 8381 50767 8415
rect 50709 8375 50767 8381
rect 51353 8415 51411 8421
rect 51353 8381 51365 8415
rect 51399 8381 51411 8415
rect 51353 8375 51411 8381
rect 51736 8344 51764 8520
rect 51810 8440 51816 8492
rect 51868 8480 51874 8492
rect 51868 8452 52224 8480
rect 51868 8440 51874 8452
rect 51902 8372 51908 8424
rect 51960 8412 51966 8424
rect 52196 8421 52224 8452
rect 51997 8415 52055 8421
rect 51997 8412 52009 8415
rect 51960 8384 52009 8412
rect 51960 8372 51966 8384
rect 51997 8381 52009 8384
rect 52043 8381 52055 8415
rect 51997 8375 52055 8381
rect 52181 8415 52239 8421
rect 52181 8381 52193 8415
rect 52227 8381 52239 8415
rect 52181 8375 52239 8381
rect 52380 8344 52408 8520
rect 52454 8508 52460 8560
rect 52512 8548 52518 8560
rect 53009 8551 53067 8557
rect 53009 8548 53021 8551
rect 52512 8520 53021 8548
rect 52512 8508 52518 8520
rect 53009 8517 53021 8520
rect 53055 8517 53067 8551
rect 53009 8511 53067 8517
rect 55401 8551 55459 8557
rect 55401 8517 55413 8551
rect 55447 8517 55459 8551
rect 55401 8511 55459 8517
rect 53101 8483 53159 8489
rect 53101 8449 53113 8483
rect 53147 8480 53159 8483
rect 53926 8480 53932 8492
rect 53147 8452 53932 8480
rect 53147 8449 53159 8452
rect 53101 8443 53159 8449
rect 53926 8440 53932 8452
rect 53984 8440 53990 8492
rect 52822 8412 52828 8424
rect 52783 8384 52828 8412
rect 52822 8372 52828 8384
rect 52880 8372 52886 8424
rect 52914 8372 52920 8424
rect 52972 8412 52978 8424
rect 52972 8384 53017 8412
rect 52972 8372 52978 8384
rect 53834 8372 53840 8424
rect 53892 8412 53898 8424
rect 54021 8415 54079 8421
rect 54021 8412 54033 8415
rect 53892 8384 54033 8412
rect 53892 8372 53898 8384
rect 54021 8381 54033 8384
rect 54067 8381 54079 8415
rect 54021 8375 54079 8381
rect 54110 8372 54116 8424
rect 54168 8412 54174 8424
rect 54277 8415 54335 8421
rect 54277 8412 54289 8415
rect 54168 8384 54289 8412
rect 54168 8372 54174 8384
rect 54277 8381 54289 8384
rect 54323 8381 54335 8415
rect 54277 8375 54335 8381
rect 54754 8372 54760 8424
rect 54812 8412 54818 8424
rect 55122 8412 55128 8424
rect 54812 8384 55128 8412
rect 54812 8372 54818 8384
rect 55122 8372 55128 8384
rect 55180 8412 55186 8424
rect 55416 8412 55444 8511
rect 56428 8489 56456 8588
rect 56413 8483 56471 8489
rect 56413 8449 56425 8483
rect 56459 8449 56471 8483
rect 56413 8443 56471 8449
rect 56594 8412 56600 8424
rect 55180 8384 55444 8412
rect 56555 8384 56600 8412
rect 55180 8372 55186 8384
rect 56594 8372 56600 8384
rect 56652 8372 56658 8424
rect 55950 8344 55956 8356
rect 50172 8316 51764 8344
rect 51920 8316 52224 8344
rect 52380 8316 55956 8344
rect 46934 8236 46940 8288
rect 46992 8276 46998 8288
rect 50614 8276 50620 8288
rect 46992 8248 50620 8276
rect 46992 8236 46998 8248
rect 50614 8236 50620 8248
rect 50672 8236 50678 8288
rect 50798 8276 50804 8288
rect 50759 8248 50804 8276
rect 50798 8236 50804 8248
rect 50856 8236 50862 8288
rect 51258 8236 51264 8288
rect 51316 8276 51322 8288
rect 51920 8276 51948 8316
rect 52086 8276 52092 8288
rect 51316 8248 51948 8276
rect 52047 8248 52092 8276
rect 51316 8236 51322 8248
rect 52086 8236 52092 8248
rect 52144 8236 52150 8288
rect 52196 8276 52224 8316
rect 55950 8304 55956 8316
rect 56008 8304 56014 8356
rect 57057 8347 57115 8353
rect 57057 8313 57069 8347
rect 57103 8344 57115 8347
rect 57977 8347 58035 8353
rect 57977 8344 57989 8347
rect 57103 8316 57989 8344
rect 57103 8313 57115 8316
rect 57057 8307 57115 8313
rect 57977 8313 57989 8316
rect 58023 8313 58035 8347
rect 58158 8344 58164 8356
rect 58119 8316 58164 8344
rect 57977 8307 58035 8313
rect 58158 8304 58164 8316
rect 58216 8304 58222 8356
rect 57422 8276 57428 8288
rect 52196 8248 57428 8276
rect 57422 8236 57428 8248
rect 57480 8236 57486 8288
rect 1104 8186 58880 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 50326 8186
rect 50378 8134 50390 8186
rect 50442 8134 50454 8186
rect 50506 8134 50518 8186
rect 50570 8134 58880 8186
rect 1104 8112 58880 8134
rect 49326 8072 49332 8084
rect 49287 8044 49332 8072
rect 49326 8032 49332 8044
rect 49384 8032 49390 8084
rect 50062 8072 50068 8084
rect 50023 8044 50068 8072
rect 50062 8032 50068 8044
rect 50120 8032 50126 8084
rect 55214 8072 55220 8084
rect 50172 8044 55220 8072
rect 3142 8004 3148 8016
rect 2516 7976 3148 8004
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2314 7936 2320 7948
rect 1903 7908 2320 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 2516 7945 2544 7976
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 47026 7964 47032 8016
rect 47084 8004 47090 8016
rect 50172 8004 50200 8044
rect 55214 8032 55220 8044
rect 55272 8032 55278 8084
rect 56689 8075 56747 8081
rect 56689 8041 56701 8075
rect 56735 8072 56747 8075
rect 57606 8072 57612 8084
rect 56735 8044 57612 8072
rect 56735 8041 56747 8044
rect 56689 8035 56747 8041
rect 57606 8032 57612 8044
rect 57664 8032 57670 8084
rect 47084 7976 50200 8004
rect 47084 7964 47090 7976
rect 50614 7964 50620 8016
rect 50672 8004 50678 8016
rect 51258 8004 51264 8016
rect 50672 7976 51264 8004
rect 50672 7964 50678 7976
rect 51258 7964 51264 7976
rect 51316 7964 51322 8016
rect 51350 7964 51356 8016
rect 51408 8004 51414 8016
rect 51896 8007 51954 8013
rect 51408 7976 51856 8004
rect 51408 7964 51414 7976
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7905 2559 7939
rect 2501 7899 2559 7905
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 3329 7939 3387 7945
rect 3329 7936 3341 7939
rect 2832 7908 3341 7936
rect 2832 7896 2838 7908
rect 3329 7905 3341 7908
rect 3375 7905 3387 7939
rect 46934 7936 46940 7948
rect 46895 7908 46940 7936
rect 3329 7899 3387 7905
rect 46934 7896 46940 7908
rect 46992 7896 46998 7948
rect 47397 7939 47455 7945
rect 47397 7905 47409 7939
rect 47443 7905 47455 7939
rect 47397 7899 47455 7905
rect 47581 7939 47639 7945
rect 47581 7905 47593 7939
rect 47627 7936 47639 7939
rect 47762 7936 47768 7948
rect 47627 7908 47768 7936
rect 47627 7905 47639 7908
rect 47581 7899 47639 7905
rect 47412 7800 47440 7899
rect 47762 7896 47768 7908
rect 47820 7896 47826 7948
rect 47946 7896 47952 7948
rect 48004 7936 48010 7948
rect 48041 7939 48099 7945
rect 48041 7936 48053 7939
rect 48004 7908 48053 7936
rect 48004 7896 48010 7908
rect 48041 7905 48053 7908
rect 48087 7905 48099 7939
rect 48041 7899 48099 7905
rect 48406 7896 48412 7948
rect 48464 7936 48470 7948
rect 48869 7939 48927 7945
rect 48869 7936 48881 7939
rect 48464 7908 48881 7936
rect 48464 7896 48470 7908
rect 48869 7905 48881 7908
rect 48915 7905 48927 7939
rect 48869 7899 48927 7905
rect 48958 7896 48964 7948
rect 49016 7936 49022 7948
rect 49510 7936 49516 7948
rect 49016 7908 49516 7936
rect 49016 7896 49022 7908
rect 49510 7896 49516 7908
rect 49568 7896 49574 7948
rect 49878 7896 49884 7948
rect 49936 7936 49942 7948
rect 49973 7939 50031 7945
rect 49973 7936 49985 7939
rect 49936 7908 49985 7936
rect 49936 7896 49942 7908
rect 49973 7905 49985 7908
rect 50019 7905 50031 7939
rect 49973 7899 50031 7905
rect 50157 7939 50215 7945
rect 50157 7905 50169 7939
rect 50203 7936 50215 7939
rect 50798 7936 50804 7948
rect 50203 7908 50804 7936
rect 50203 7905 50215 7908
rect 50157 7899 50215 7905
rect 50798 7896 50804 7908
rect 50856 7896 50862 7948
rect 50982 7896 50988 7948
rect 51040 7936 51046 7948
rect 51629 7939 51687 7945
rect 51629 7936 51641 7939
rect 51040 7908 51641 7936
rect 51040 7896 51046 7908
rect 51629 7905 51641 7908
rect 51675 7905 51687 7939
rect 51828 7936 51856 7976
rect 51896 7973 51908 8007
rect 51942 8004 51954 8007
rect 52086 8004 52092 8016
rect 51942 7976 52092 8004
rect 51942 7973 51954 7976
rect 51896 7967 51954 7973
rect 52086 7964 52092 7976
rect 52144 7964 52150 8016
rect 54938 8004 54944 8016
rect 52932 7976 54944 8004
rect 52932 7948 52960 7976
rect 54938 7964 54944 7976
rect 54996 8004 55002 8016
rect 54996 7976 55260 8004
rect 54996 7964 55002 7976
rect 52914 7936 52920 7948
rect 51828 7908 52920 7936
rect 51629 7899 51687 7905
rect 52914 7896 52920 7908
rect 52972 7896 52978 7948
rect 53190 7896 53196 7948
rect 53248 7936 53254 7948
rect 53561 7939 53619 7945
rect 53561 7936 53573 7939
rect 53248 7908 53573 7936
rect 53248 7896 53254 7908
rect 53561 7905 53573 7908
rect 53607 7905 53619 7939
rect 53721 7939 53779 7945
rect 53721 7936 53733 7939
rect 53561 7899 53619 7905
rect 53659 7908 53733 7936
rect 47489 7871 47547 7877
rect 47489 7837 47501 7871
rect 47535 7868 47547 7871
rect 51534 7868 51540 7880
rect 47535 7840 51540 7868
rect 47535 7837 47547 7840
rect 47489 7831 47547 7837
rect 51534 7828 51540 7840
rect 51592 7828 51598 7880
rect 53469 7871 53527 7877
rect 53469 7837 53481 7871
rect 53515 7868 53527 7871
rect 53659 7868 53687 7908
rect 53721 7905 53733 7908
rect 53767 7905 53779 7939
rect 53721 7899 53779 7905
rect 54665 7939 54723 7945
rect 54665 7905 54677 7939
rect 54711 7936 54723 7939
rect 54754 7936 54760 7948
rect 54711 7908 54760 7936
rect 54711 7905 54723 7908
rect 54665 7899 54723 7905
rect 54754 7896 54760 7908
rect 54812 7896 54818 7948
rect 55122 7936 55128 7948
rect 55083 7908 55128 7936
rect 55122 7896 55128 7908
rect 55180 7896 55186 7948
rect 55232 7945 55260 7976
rect 55217 7939 55275 7945
rect 55217 7905 55229 7939
rect 55263 7905 55275 7939
rect 55217 7899 55275 7905
rect 56778 7896 56784 7948
rect 56836 7936 56842 7948
rect 56873 7939 56931 7945
rect 56873 7936 56885 7939
rect 56836 7908 56885 7936
rect 56836 7896 56842 7908
rect 56873 7905 56885 7908
rect 56919 7905 56931 7939
rect 56873 7899 56931 7905
rect 53515 7840 53687 7868
rect 54389 7871 54447 7877
rect 53515 7837 53527 7840
rect 53469 7831 53527 7837
rect 54389 7837 54401 7871
rect 54435 7868 54447 7871
rect 56962 7868 56968 7880
rect 54435 7840 56968 7868
rect 54435 7837 54447 7840
rect 54389 7831 54447 7837
rect 56962 7828 56968 7840
rect 57020 7828 57026 7880
rect 57330 7868 57336 7880
rect 57291 7840 57336 7868
rect 57330 7828 57336 7840
rect 57388 7828 57394 7880
rect 57517 7871 57575 7877
rect 57517 7837 57529 7871
rect 57563 7837 57575 7871
rect 57517 7831 57575 7837
rect 48685 7803 48743 7809
rect 47412 7772 48636 7800
rect 1946 7732 1952 7744
rect 1907 7704 1952 7732
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2685 7735 2743 7741
rect 2685 7701 2697 7735
rect 2731 7732 2743 7735
rect 2774 7732 2780 7744
rect 2731 7704 2780 7732
rect 2731 7701 2743 7704
rect 2685 7695 2743 7701
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3142 7732 3148 7744
rect 3103 7704 3148 7732
rect 3142 7692 3148 7704
rect 3200 7692 3206 7744
rect 47762 7692 47768 7744
rect 47820 7732 47826 7744
rect 48225 7735 48283 7741
rect 48225 7732 48237 7735
rect 47820 7704 48237 7732
rect 47820 7692 47826 7704
rect 48225 7701 48237 7704
rect 48271 7701 48283 7735
rect 48608 7732 48636 7772
rect 48685 7769 48697 7803
rect 48731 7800 48743 7803
rect 57532 7800 57560 7831
rect 48731 7772 51672 7800
rect 48731 7769 48743 7772
rect 48685 7763 48743 7769
rect 51350 7732 51356 7744
rect 48608 7704 51356 7732
rect 48225 7695 48283 7701
rect 51350 7692 51356 7704
rect 51408 7692 51414 7744
rect 51644 7732 51672 7772
rect 52656 7772 57560 7800
rect 52656 7732 52684 7772
rect 51644 7704 52684 7732
rect 53009 7735 53067 7741
rect 53009 7701 53021 7735
rect 53055 7732 53067 7735
rect 53466 7732 53472 7744
rect 53055 7704 53472 7732
rect 53055 7701 53067 7704
rect 53009 7695 53067 7701
rect 53466 7692 53472 7704
rect 53524 7692 53530 7744
rect 53558 7692 53564 7744
rect 53616 7732 53622 7744
rect 54389 7735 54447 7741
rect 53616 7704 53661 7732
rect 53616 7692 53622 7704
rect 54389 7701 54401 7735
rect 54435 7732 54447 7735
rect 54481 7735 54539 7741
rect 54481 7732 54493 7735
rect 54435 7704 54493 7732
rect 54435 7701 54447 7704
rect 54389 7695 54447 7701
rect 54481 7701 54493 7704
rect 54527 7701 54539 7735
rect 54481 7695 54539 7701
rect 54754 7692 54760 7744
rect 54812 7732 54818 7744
rect 55490 7732 55496 7744
rect 54812 7704 55496 7732
rect 54812 7692 54818 7704
rect 55490 7692 55496 7704
rect 55548 7732 55554 7744
rect 55858 7732 55864 7744
rect 55548 7704 55864 7732
rect 55548 7692 55554 7704
rect 55858 7692 55864 7704
rect 55916 7692 55922 7744
rect 56870 7692 56876 7744
rect 56928 7732 56934 7744
rect 57701 7735 57759 7741
rect 57701 7732 57713 7735
rect 56928 7704 57713 7732
rect 56928 7692 56934 7704
rect 57701 7701 57713 7704
rect 57747 7701 57759 7735
rect 57701 7695 57759 7701
rect 1104 7642 58880 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 58880 7642
rect 1104 7568 58880 7590
rect 1854 7488 1860 7540
rect 1912 7528 1918 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1912 7500 2053 7528
rect 1912 7488 1918 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 47578 7488 47584 7540
rect 47636 7528 47642 7540
rect 47946 7528 47952 7540
rect 47636 7500 47952 7528
rect 47636 7488 47642 7500
rect 47946 7488 47952 7500
rect 48004 7528 48010 7540
rect 49694 7528 49700 7540
rect 48004 7500 49700 7528
rect 48004 7488 48010 7500
rect 49694 7488 49700 7500
rect 49752 7488 49758 7540
rect 50709 7531 50767 7537
rect 50709 7497 50721 7531
rect 50755 7528 50767 7531
rect 51442 7528 51448 7540
rect 50755 7500 51304 7528
rect 51403 7500 51448 7528
rect 50755 7497 50767 7500
rect 50709 7491 50767 7497
rect 49602 7420 49608 7472
rect 49660 7460 49666 7472
rect 49789 7463 49847 7469
rect 49789 7460 49801 7463
rect 49660 7432 49801 7460
rect 49660 7420 49666 7432
rect 49789 7429 49801 7432
rect 49835 7429 49847 7463
rect 51276 7460 51304 7500
rect 51442 7488 51448 7500
rect 51500 7488 51506 7540
rect 51534 7488 51540 7540
rect 51592 7528 51598 7540
rect 55769 7531 55827 7537
rect 51592 7500 54984 7528
rect 51592 7488 51598 7500
rect 51718 7460 51724 7472
rect 49789 7423 49847 7429
rect 49896 7432 50476 7460
rect 51276 7432 51724 7460
rect 49896 7401 49924 7432
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 1719 7364 2973 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2961 7361 2973 7364
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 49881 7395 49939 7401
rect 49881 7361 49893 7395
rect 49927 7361 49939 7395
rect 49881 7355 49939 7361
rect 50154 7352 50160 7404
rect 50212 7392 50218 7404
rect 50341 7395 50399 7401
rect 50341 7392 50353 7395
rect 50212 7364 50353 7392
rect 50212 7352 50218 7364
rect 50341 7361 50353 7364
rect 50387 7361 50399 7395
rect 50448 7392 50476 7432
rect 51718 7420 51724 7432
rect 51776 7420 51782 7472
rect 52733 7463 52791 7469
rect 52733 7429 52745 7463
rect 52779 7460 52791 7463
rect 52822 7460 52828 7472
rect 52779 7432 52828 7460
rect 52779 7429 52791 7432
rect 52733 7423 52791 7429
rect 52822 7420 52828 7432
rect 52880 7420 52886 7472
rect 50798 7392 50804 7404
rect 50448 7364 50804 7392
rect 50341 7355 50399 7361
rect 50798 7352 50804 7364
rect 50856 7392 50862 7404
rect 51445 7395 51503 7401
rect 51445 7392 51457 7395
rect 50856 7364 51457 7392
rect 50856 7352 50862 7364
rect 51445 7361 51457 7364
rect 51491 7361 51503 7395
rect 51445 7355 51503 7361
rect 51626 7352 51632 7404
rect 51684 7392 51690 7404
rect 53650 7392 53656 7404
rect 51684 7364 53656 7392
rect 51684 7352 51690 7364
rect 53650 7352 53656 7364
rect 53708 7352 53714 7404
rect 54113 7395 54171 7401
rect 54113 7361 54125 7395
rect 54159 7392 54171 7395
rect 54570 7392 54576 7404
rect 54159 7364 54576 7392
rect 54159 7361 54171 7364
rect 54113 7355 54171 7361
rect 54570 7352 54576 7364
rect 54628 7392 54634 7404
rect 54956 7392 54984 7500
rect 55769 7497 55781 7531
rect 55815 7528 55827 7531
rect 57698 7528 57704 7540
rect 55815 7500 57704 7528
rect 55815 7497 55827 7500
rect 55769 7491 55827 7497
rect 57698 7488 57704 7500
rect 57756 7488 57762 7540
rect 56413 7395 56471 7401
rect 56413 7392 56425 7395
rect 54628 7364 54892 7392
rect 54956 7364 56425 7392
rect 54628 7352 54634 7364
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 3142 7324 3148 7336
rect 1903 7296 3148 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 3142 7284 3148 7296
rect 3200 7284 3206 7336
rect 46566 7324 46572 7336
rect 46527 7296 46572 7324
rect 46566 7284 46572 7296
rect 46624 7284 46630 7336
rect 46937 7327 46995 7333
rect 46937 7293 46949 7327
rect 46983 7324 46995 7327
rect 47210 7324 47216 7336
rect 46983 7296 47216 7324
rect 46983 7293 46995 7296
rect 46937 7287 46995 7293
rect 47210 7284 47216 7296
rect 47268 7284 47274 7336
rect 47854 7324 47860 7336
rect 47815 7296 47860 7324
rect 47854 7284 47860 7296
rect 47912 7284 47918 7336
rect 48958 7324 48964 7336
rect 48919 7296 48964 7324
rect 48958 7284 48964 7296
rect 49016 7284 49022 7336
rect 49605 7327 49663 7333
rect 49605 7293 49617 7327
rect 49651 7324 49663 7327
rect 50614 7324 50620 7336
rect 49651 7296 50620 7324
rect 49651 7293 49663 7296
rect 49605 7287 49663 7293
rect 50614 7284 50620 7296
rect 50672 7324 50678 7336
rect 51353 7327 51411 7333
rect 51353 7324 51365 7327
rect 50672 7296 51365 7324
rect 50672 7284 50678 7296
rect 51353 7293 51365 7296
rect 51399 7293 51411 7327
rect 51353 7287 51411 7293
rect 52178 7284 52184 7336
rect 52236 7324 52242 7336
rect 52549 7327 52607 7333
rect 52549 7324 52561 7327
rect 52236 7296 52561 7324
rect 52236 7284 52242 7296
rect 52549 7293 52561 7296
rect 52595 7293 52607 7327
rect 52549 7287 52607 7293
rect 52825 7327 52883 7333
rect 52825 7293 52837 7327
rect 52871 7324 52883 7327
rect 53282 7324 53288 7336
rect 52871 7296 53288 7324
rect 52871 7293 52883 7296
rect 52825 7287 52883 7293
rect 53282 7284 53288 7296
rect 53340 7284 53346 7336
rect 53466 7284 53472 7336
rect 53524 7324 53530 7336
rect 54021 7327 54079 7333
rect 54021 7324 54033 7327
rect 53524 7296 54033 7324
rect 53524 7284 53530 7296
rect 54021 7293 54033 7296
rect 54067 7293 54079 7327
rect 54021 7287 54079 7293
rect 54386 7284 54392 7336
rect 54444 7324 54450 7336
rect 54864 7333 54892 7364
rect 56413 7361 56425 7364
rect 56459 7361 56471 7395
rect 56778 7392 56784 7404
rect 56413 7355 56471 7361
rect 56520 7364 56784 7392
rect 54665 7327 54723 7333
rect 54665 7324 54677 7327
rect 54444 7296 54677 7324
rect 54444 7284 54450 7296
rect 54665 7293 54677 7296
rect 54711 7293 54723 7327
rect 54665 7287 54723 7293
rect 54849 7327 54907 7333
rect 54849 7293 54861 7327
rect 54895 7293 54907 7327
rect 54849 7287 54907 7293
rect 55953 7327 56011 7333
rect 55953 7293 55965 7327
rect 55999 7324 56011 7327
rect 56520 7324 56548 7364
rect 56778 7352 56784 7364
rect 56836 7352 56842 7404
rect 58158 7392 58164 7404
rect 58119 7364 58164 7392
rect 58158 7352 58164 7364
rect 58216 7352 58222 7404
rect 55999 7296 56548 7324
rect 56597 7327 56655 7333
rect 55999 7293 56011 7296
rect 55953 7287 56011 7293
rect 56597 7293 56609 7327
rect 56643 7293 56655 7327
rect 56597 7287 56655 7293
rect 56612 7256 56640 7287
rect 57974 7256 57980 7268
rect 48792 7228 56640 7256
rect 57935 7228 57980 7256
rect 48792 7197 48820 7228
rect 57974 7216 57980 7228
rect 58032 7216 58038 7268
rect 48777 7191 48835 7197
rect 48777 7157 48789 7191
rect 48823 7157 48835 7191
rect 48777 7151 48835 7157
rect 49421 7191 49479 7197
rect 49421 7157 49433 7191
rect 49467 7188 49479 7191
rect 50154 7188 50160 7200
rect 49467 7160 50160 7188
rect 49467 7157 49479 7160
rect 49421 7151 49479 7157
rect 50154 7148 50160 7160
rect 50212 7148 50218 7200
rect 50706 7188 50712 7200
rect 50667 7160 50712 7188
rect 50706 7148 50712 7160
rect 50764 7148 50770 7200
rect 50890 7188 50896 7200
rect 50851 7160 50896 7188
rect 50890 7148 50896 7160
rect 50948 7148 50954 7200
rect 52086 7148 52092 7200
rect 52144 7188 52150 7200
rect 52365 7191 52423 7197
rect 52365 7188 52377 7191
rect 52144 7160 52377 7188
rect 52144 7148 52150 7160
rect 52365 7157 52377 7160
rect 52411 7157 52423 7191
rect 54754 7188 54760 7200
rect 54715 7160 54760 7188
rect 52365 7151 52423 7157
rect 54754 7148 54760 7160
rect 54812 7148 54818 7200
rect 57054 7188 57060 7200
rect 57015 7160 57060 7188
rect 57054 7148 57060 7160
rect 57112 7148 57118 7200
rect 1104 7098 58880 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 50326 7098
rect 50378 7046 50390 7098
rect 50442 7046 50454 7098
rect 50506 7046 50518 7098
rect 50570 7046 58880 7098
rect 1104 7024 58880 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 46566 6944 46572 6996
rect 46624 6984 46630 6996
rect 52086 6984 52092 6996
rect 46624 6956 51948 6984
rect 52047 6956 52092 6984
rect 46624 6944 46630 6956
rect 47854 6876 47860 6928
rect 47912 6916 47918 6928
rect 51626 6916 51632 6928
rect 47912 6888 51632 6916
rect 47912 6876 47918 6888
rect 51626 6876 51632 6888
rect 51684 6876 51690 6928
rect 51920 6916 51948 6956
rect 52086 6944 52092 6956
rect 52144 6944 52150 6996
rect 52730 6944 52736 6996
rect 52788 6984 52794 6996
rect 53377 6987 53435 6993
rect 53377 6984 53389 6987
rect 52788 6956 53389 6984
rect 52788 6944 52794 6956
rect 53377 6953 53389 6956
rect 53423 6953 53435 6987
rect 57514 6984 57520 6996
rect 53377 6947 53435 6953
rect 53484 6956 57520 6984
rect 53484 6916 53512 6956
rect 57514 6944 57520 6956
rect 57572 6944 57578 6996
rect 57974 6944 57980 6996
rect 58032 6984 58038 6996
rect 58161 6987 58219 6993
rect 58161 6984 58173 6987
rect 58032 6956 58173 6984
rect 58032 6944 58038 6956
rect 58161 6953 58173 6956
rect 58207 6953 58219 6987
rect 58161 6947 58219 6953
rect 51920 6888 53512 6916
rect 54472 6919 54530 6925
rect 54472 6885 54484 6919
rect 54518 6916 54530 6919
rect 54754 6916 54760 6928
rect 54518 6888 54760 6916
rect 54518 6885 54530 6888
rect 54472 6879 54530 6885
rect 54754 6876 54760 6888
rect 54812 6876 54818 6928
rect 56873 6919 56931 6925
rect 56873 6885 56885 6919
rect 56919 6916 56931 6919
rect 57054 6916 57060 6928
rect 56919 6888 57060 6916
rect 56919 6885 56931 6888
rect 56873 6879 56931 6885
rect 57054 6876 57060 6888
rect 57112 6876 57118 6928
rect 1673 6851 1731 6857
rect 1673 6817 1685 6851
rect 1719 6848 1731 6851
rect 2961 6851 3019 6857
rect 2961 6848 2973 6851
rect 1719 6820 2973 6848
rect 1719 6817 1731 6820
rect 1673 6811 1731 6817
rect 2961 6817 2973 6820
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 45097 6851 45155 6857
rect 45097 6817 45109 6851
rect 45143 6848 45155 6851
rect 45186 6848 45192 6860
rect 45143 6820 45192 6848
rect 45143 6817 45155 6820
rect 45097 6811 45155 6817
rect 45186 6808 45192 6820
rect 45244 6808 45250 6860
rect 47581 6851 47639 6857
rect 47581 6817 47593 6851
rect 47627 6848 47639 6851
rect 48774 6848 48780 6860
rect 47627 6820 48780 6848
rect 47627 6817 47639 6820
rect 47581 6811 47639 6817
rect 48774 6808 48780 6820
rect 48832 6808 48838 6860
rect 48952 6851 49010 6857
rect 48952 6817 48964 6851
rect 48998 6848 49010 6851
rect 50890 6848 50896 6860
rect 48998 6820 50896 6848
rect 48998 6817 49010 6820
rect 48952 6811 49010 6817
rect 50890 6808 50896 6820
rect 50948 6808 50954 6860
rect 51813 6851 51871 6857
rect 51813 6817 51825 6851
rect 51859 6848 51871 6851
rect 52086 6848 52092 6860
rect 51859 6820 52092 6848
rect 51859 6817 51871 6820
rect 51813 6811 51871 6817
rect 52086 6808 52092 6820
rect 52144 6808 52150 6860
rect 53190 6848 53196 6860
rect 53151 6820 53196 6848
rect 53190 6808 53196 6820
rect 53248 6808 53254 6860
rect 53374 6848 53380 6860
rect 53335 6820 53380 6848
rect 53374 6808 53380 6820
rect 53432 6808 53438 6860
rect 55306 6848 55312 6860
rect 53484 6820 55312 6848
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6780 1915 6783
rect 2498 6780 2504 6792
rect 1903 6752 2504 6780
rect 1903 6749 1915 6752
rect 1857 6743 1915 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 48682 6780 48688 6792
rect 48643 6752 48688 6780
rect 48682 6740 48688 6752
rect 48740 6740 48746 6792
rect 49694 6740 49700 6792
rect 49752 6780 49758 6792
rect 50798 6780 50804 6792
rect 49752 6752 50804 6780
rect 49752 6740 49758 6752
rect 50798 6740 50804 6752
rect 50856 6740 50862 6792
rect 51629 6783 51687 6789
rect 51629 6749 51641 6783
rect 51675 6780 51687 6783
rect 52181 6783 52239 6789
rect 52181 6780 52193 6783
rect 51675 6752 52193 6780
rect 51675 6749 51687 6752
rect 51629 6743 51687 6749
rect 52181 6749 52193 6752
rect 52227 6780 52239 6783
rect 52730 6780 52736 6792
rect 52227 6752 52736 6780
rect 52227 6749 52239 6752
rect 52181 6743 52239 6749
rect 52730 6740 52736 6752
rect 52788 6740 52794 6792
rect 46937 6715 46995 6721
rect 46937 6681 46949 6715
rect 46983 6712 46995 6715
rect 51534 6712 51540 6724
rect 46983 6684 48728 6712
rect 46983 6681 46995 6684
rect 46937 6675 46995 6681
rect 48225 6647 48283 6653
rect 48225 6613 48237 6647
rect 48271 6644 48283 6647
rect 48590 6644 48596 6656
rect 48271 6616 48596 6644
rect 48271 6613 48283 6616
rect 48225 6607 48283 6613
rect 48590 6604 48596 6616
rect 48648 6604 48654 6656
rect 48700 6644 48728 6684
rect 49620 6684 51540 6712
rect 49620 6644 49648 6684
rect 51534 6672 51540 6684
rect 51592 6672 51598 6724
rect 51902 6712 51908 6724
rect 51863 6684 51908 6712
rect 51902 6672 51908 6684
rect 51960 6672 51966 6724
rect 53484 6712 53512 6820
rect 55306 6808 55312 6820
rect 55364 6808 55370 6860
rect 56962 6808 56968 6860
rect 57020 6848 57026 6860
rect 57701 6851 57759 6857
rect 57701 6848 57713 6851
rect 57020 6820 57713 6848
rect 57020 6808 57026 6820
rect 57701 6817 57713 6820
rect 57747 6817 57759 6851
rect 57701 6811 57759 6817
rect 53558 6740 53564 6792
rect 53616 6780 53622 6792
rect 53745 6783 53803 6789
rect 53745 6780 53757 6783
rect 53616 6752 53757 6780
rect 53616 6740 53622 6752
rect 53745 6749 53757 6752
rect 53791 6749 53803 6783
rect 53745 6743 53803 6749
rect 53834 6740 53840 6792
rect 53892 6780 53898 6792
rect 54205 6783 54263 6789
rect 54205 6780 54217 6783
rect 53892 6752 54217 6780
rect 53892 6740 53898 6752
rect 54205 6749 54217 6752
rect 54251 6749 54263 6783
rect 54205 6743 54263 6749
rect 57057 6783 57115 6789
rect 57057 6749 57069 6783
rect 57103 6780 57115 6783
rect 57146 6780 57152 6792
rect 57103 6752 57152 6780
rect 57103 6749 57115 6752
rect 57057 6743 57115 6749
rect 57146 6740 57152 6752
rect 57204 6740 57210 6792
rect 57422 6740 57428 6792
rect 57480 6780 57486 6792
rect 57517 6783 57575 6789
rect 57517 6780 57529 6783
rect 57480 6752 57529 6780
rect 57480 6740 57486 6752
rect 57517 6749 57529 6752
rect 57563 6749 57575 6783
rect 57517 6743 57575 6749
rect 52012 6684 53512 6712
rect 48700 6616 49648 6644
rect 49694 6604 49700 6656
rect 49752 6644 49758 6656
rect 49970 6644 49976 6656
rect 49752 6616 49976 6644
rect 49752 6604 49758 6616
rect 49970 6604 49976 6616
rect 50028 6604 50034 6656
rect 50065 6647 50123 6653
rect 50065 6613 50077 6647
rect 50111 6644 50123 6647
rect 50430 6644 50436 6656
rect 50111 6616 50436 6644
rect 50111 6613 50123 6616
rect 50065 6607 50123 6613
rect 50430 6604 50436 6616
rect 50488 6604 50494 6656
rect 51166 6604 51172 6656
rect 51224 6644 51230 6656
rect 52012 6644 52040 6684
rect 51224 6616 52040 6644
rect 51224 6604 51230 6616
rect 53190 6604 53196 6656
rect 53248 6644 53254 6656
rect 55214 6644 55220 6656
rect 53248 6616 55220 6644
rect 53248 6604 53254 6616
rect 55214 6604 55220 6616
rect 55272 6644 55278 6656
rect 55585 6647 55643 6653
rect 55585 6644 55597 6647
rect 55272 6616 55597 6644
rect 55272 6604 55278 6616
rect 55585 6613 55597 6616
rect 55631 6613 55643 6647
rect 55585 6607 55643 6613
rect 1104 6554 58880 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 58880 6554
rect 1104 6480 58880 6502
rect 2498 6440 2504 6452
rect 2459 6412 2504 6440
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 46569 6443 46627 6449
rect 46569 6409 46581 6443
rect 46615 6440 46627 6443
rect 51810 6440 51816 6452
rect 46615 6412 51816 6440
rect 46615 6409 46627 6412
rect 46569 6403 46627 6409
rect 51810 6400 51816 6412
rect 51868 6400 51874 6452
rect 52362 6440 52368 6452
rect 52323 6412 52368 6440
rect 52362 6400 52368 6412
rect 52420 6400 52426 6452
rect 53282 6400 53288 6452
rect 53340 6440 53346 6452
rect 54202 6440 54208 6452
rect 53340 6412 54208 6440
rect 53340 6400 53346 6412
rect 54202 6400 54208 6412
rect 54260 6400 54266 6452
rect 47688 6344 54524 6372
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 2774 6236 2780 6248
rect 2731 6208 2780 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3326 6236 3332 6248
rect 3287 6208 3332 6236
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 44453 6239 44511 6245
rect 44453 6205 44465 6239
rect 44499 6205 44511 6239
rect 44453 6199 44511 6205
rect 45005 6239 45063 6245
rect 45005 6205 45017 6239
rect 45051 6236 45063 6239
rect 45278 6236 45284 6248
rect 45051 6208 45284 6236
rect 45051 6205 45063 6208
rect 45005 6199 45063 6205
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 2314 6168 2320 6180
rect 1903 6140 2320 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 2314 6128 2320 6140
rect 2372 6128 2378 6180
rect 44468 6168 44496 6199
rect 45278 6196 45284 6208
rect 45336 6196 45342 6248
rect 45649 6239 45707 6245
rect 45649 6205 45661 6239
rect 45695 6236 45707 6239
rect 45925 6239 45983 6245
rect 45925 6236 45937 6239
rect 45695 6208 45937 6236
rect 45695 6205 45707 6208
rect 45649 6199 45707 6205
rect 45925 6205 45937 6208
rect 45971 6236 45983 6239
rect 46474 6236 46480 6248
rect 45971 6208 46480 6236
rect 45971 6205 45983 6208
rect 45925 6199 45983 6205
rect 46474 6196 46480 6208
rect 46532 6196 46538 6248
rect 47688 6245 47716 6344
rect 47765 6307 47823 6313
rect 47765 6273 47777 6307
rect 47811 6304 47823 6307
rect 50890 6304 50896 6316
rect 47811 6276 50896 6304
rect 47811 6273 47823 6276
rect 47765 6267 47823 6273
rect 50890 6264 50896 6276
rect 50948 6264 50954 6316
rect 51534 6264 51540 6316
rect 51592 6304 51598 6316
rect 52454 6304 52460 6316
rect 51592 6276 52460 6304
rect 51592 6264 51598 6276
rect 52454 6264 52460 6276
rect 52512 6264 52518 6316
rect 52730 6304 52736 6316
rect 52691 6276 52736 6304
rect 52730 6264 52736 6276
rect 52788 6264 52794 6316
rect 53558 6264 53564 6316
rect 53616 6304 53622 6316
rect 54496 6313 54524 6344
rect 54389 6307 54447 6313
rect 54389 6304 54401 6307
rect 53616 6276 54401 6304
rect 53616 6264 53622 6276
rect 54389 6273 54401 6276
rect 54435 6273 54447 6307
rect 54389 6267 54447 6273
rect 54481 6307 54539 6313
rect 54481 6273 54493 6307
rect 54527 6304 54539 6307
rect 55309 6307 55367 6313
rect 55309 6304 55321 6307
rect 54527 6276 55321 6304
rect 54527 6273 54539 6276
rect 54481 6267 54539 6273
rect 55309 6273 55321 6276
rect 55355 6273 55367 6307
rect 57514 6304 57520 6316
rect 57475 6276 57520 6304
rect 55309 6267 55367 6273
rect 57514 6264 57520 6276
rect 57572 6264 57578 6316
rect 47213 6239 47271 6245
rect 47213 6205 47225 6239
rect 47259 6205 47271 6239
rect 47213 6199 47271 6205
rect 47673 6239 47731 6245
rect 47673 6205 47685 6239
rect 47719 6205 47731 6239
rect 47673 6199 47731 6205
rect 47857 6239 47915 6245
rect 47857 6205 47869 6239
rect 47903 6205 47915 6239
rect 47857 6199 47915 6205
rect 45370 6168 45376 6180
rect 44468 6140 45376 6168
rect 45370 6128 45376 6140
rect 45428 6128 45434 6180
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 47228 6100 47256 6199
rect 47762 6128 47768 6180
rect 47820 6168 47826 6180
rect 47872 6168 47900 6199
rect 48314 6196 48320 6248
rect 48372 6236 48378 6248
rect 49053 6239 49111 6245
rect 49053 6236 49065 6239
rect 48372 6208 49065 6236
rect 48372 6196 48378 6208
rect 49053 6205 49065 6208
rect 49099 6205 49111 6239
rect 49510 6236 49516 6248
rect 49471 6208 49516 6236
rect 49053 6199 49111 6205
rect 49510 6196 49516 6208
rect 49568 6196 49574 6248
rect 50157 6239 50215 6245
rect 50157 6236 50169 6239
rect 49988 6208 50169 6236
rect 47820 6140 47900 6168
rect 47820 6128 47826 6140
rect 49418 6128 49424 6180
rect 49476 6168 49482 6180
rect 49988 6168 50016 6208
rect 50157 6205 50169 6208
rect 50203 6205 50215 6239
rect 50430 6236 50436 6248
rect 50391 6208 50436 6236
rect 50157 6199 50215 6205
rect 50430 6196 50436 6208
rect 50488 6196 50494 6248
rect 50525 6239 50583 6245
rect 50525 6205 50537 6239
rect 50571 6236 50583 6239
rect 50706 6236 50712 6248
rect 50571 6208 50712 6236
rect 50571 6205 50583 6208
rect 50525 6199 50583 6205
rect 50706 6196 50712 6208
rect 50764 6196 50770 6248
rect 51169 6239 51227 6245
rect 51169 6205 51181 6239
rect 51215 6205 51227 6239
rect 51169 6199 51227 6205
rect 49476 6140 50016 6168
rect 49476 6128 49482 6140
rect 50062 6128 50068 6180
rect 50120 6168 50126 6180
rect 50341 6171 50399 6177
rect 50341 6168 50353 6171
rect 50120 6140 50353 6168
rect 50120 6128 50126 6140
rect 50341 6137 50353 6140
rect 50387 6168 50399 6171
rect 51184 6168 51212 6199
rect 51258 6196 51264 6248
rect 51316 6236 51322 6248
rect 51353 6239 51411 6245
rect 51353 6236 51365 6239
rect 51316 6208 51365 6236
rect 51316 6196 51322 6208
rect 51353 6205 51365 6208
rect 51399 6205 51411 6239
rect 51353 6199 51411 6205
rect 51629 6239 51687 6245
rect 51629 6205 51641 6239
rect 51675 6236 51687 6239
rect 52086 6236 52092 6248
rect 51675 6208 52092 6236
rect 51675 6205 51687 6208
rect 51629 6199 51687 6205
rect 52086 6196 52092 6208
rect 52144 6236 52150 6248
rect 52549 6239 52607 6245
rect 52549 6236 52561 6239
rect 52144 6208 52561 6236
rect 52144 6196 52150 6208
rect 52549 6205 52561 6208
rect 52595 6205 52607 6239
rect 52549 6199 52607 6205
rect 52638 6196 52644 6248
rect 52696 6236 52702 6248
rect 52825 6239 52883 6245
rect 52696 6208 52741 6236
rect 52696 6196 52702 6208
rect 52825 6205 52837 6239
rect 52871 6236 52883 6239
rect 54018 6236 54024 6248
rect 52871 6208 54024 6236
rect 52871 6205 52883 6208
rect 52825 6199 52883 6205
rect 54018 6196 54024 6208
rect 54076 6196 54082 6248
rect 54202 6236 54208 6248
rect 54163 6208 54208 6236
rect 54202 6196 54208 6208
rect 54260 6196 54266 6248
rect 54294 6196 54300 6248
rect 54352 6236 54358 6248
rect 54352 6208 54397 6236
rect 54352 6196 54358 6208
rect 54570 6196 54576 6248
rect 54628 6236 54634 6248
rect 54665 6239 54723 6245
rect 54665 6236 54677 6239
rect 54628 6208 54677 6236
rect 54628 6196 54634 6208
rect 54665 6205 54677 6208
rect 54711 6205 54723 6239
rect 55214 6236 55220 6248
rect 55175 6208 55220 6236
rect 54665 6199 54723 6205
rect 55214 6196 55220 6208
rect 55272 6196 55278 6248
rect 56413 6239 56471 6245
rect 56413 6205 56425 6239
rect 56459 6205 56471 6239
rect 56413 6199 56471 6205
rect 51718 6168 51724 6180
rect 50387 6140 51212 6168
rect 51679 6140 51724 6168
rect 50387 6137 50399 6140
rect 50341 6131 50399 6137
rect 51718 6128 51724 6140
rect 51776 6128 51782 6180
rect 56428 6168 56456 6199
rect 56502 6196 56508 6248
rect 56560 6236 56566 6248
rect 56597 6239 56655 6245
rect 56597 6236 56609 6239
rect 56560 6208 56609 6236
rect 56560 6196 56566 6208
rect 56597 6205 56609 6208
rect 56643 6205 56655 6239
rect 56597 6199 56655 6205
rect 57701 6239 57759 6245
rect 57701 6205 57713 6239
rect 57747 6236 57759 6239
rect 58066 6236 58072 6248
rect 57747 6208 58072 6236
rect 57747 6205 57759 6208
rect 57701 6199 57759 6205
rect 58066 6196 58072 6208
rect 58124 6196 58130 6248
rect 52380 6140 56456 6168
rect 48682 6100 48688 6112
rect 47228 6072 48688 6100
rect 48682 6060 48688 6072
rect 48740 6060 48746 6112
rect 48866 6100 48872 6112
rect 48827 6072 48872 6100
rect 48866 6060 48872 6072
rect 48924 6060 48930 6112
rect 48958 6060 48964 6112
rect 49016 6100 49022 6112
rect 49602 6100 49608 6112
rect 49016 6072 49608 6100
rect 49016 6060 49022 6072
rect 49602 6060 49608 6072
rect 49660 6100 49666 6112
rect 49697 6103 49755 6109
rect 49697 6100 49709 6103
rect 49660 6072 49709 6100
rect 49660 6060 49666 6072
rect 49697 6069 49709 6072
rect 49743 6069 49755 6103
rect 49697 6063 49755 6069
rect 50614 6060 50620 6112
rect 50672 6100 50678 6112
rect 50709 6103 50767 6109
rect 50709 6100 50721 6103
rect 50672 6072 50721 6100
rect 50672 6060 50678 6072
rect 50709 6069 50721 6072
rect 50755 6069 50767 6103
rect 50709 6063 50767 6069
rect 50890 6060 50896 6112
rect 50948 6100 50954 6112
rect 52380 6100 52408 6140
rect 50948 6072 52408 6100
rect 50948 6060 50954 6072
rect 52454 6060 52460 6112
rect 52512 6100 52518 6112
rect 53190 6100 53196 6112
rect 52512 6072 53196 6100
rect 52512 6060 52518 6072
rect 53190 6060 53196 6072
rect 53248 6060 53254 6112
rect 53742 6060 53748 6112
rect 53800 6100 53806 6112
rect 54021 6103 54079 6109
rect 54021 6100 54033 6103
rect 53800 6072 54033 6100
rect 53800 6060 53806 6072
rect 54021 6069 54033 6072
rect 54067 6069 54079 6103
rect 57054 6100 57060 6112
rect 57015 6072 57060 6100
rect 54021 6063 54079 6069
rect 57054 6060 57060 6072
rect 57112 6060 57118 6112
rect 57974 6060 57980 6112
rect 58032 6100 58038 6112
rect 58161 6103 58219 6109
rect 58161 6100 58173 6103
rect 58032 6072 58173 6100
rect 58032 6060 58038 6072
rect 58161 6069 58173 6072
rect 58207 6069 58219 6103
rect 58161 6063 58219 6069
rect 1104 6010 58880 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 50326 6010
rect 50378 5958 50390 6010
rect 50442 5958 50454 6010
rect 50506 5958 50518 6010
rect 50570 5958 58880 6010
rect 1104 5936 58880 5958
rect 2314 5896 2320 5908
rect 2275 5868 2320 5896
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 46492 5868 51028 5896
rect 2774 5788 2780 5840
rect 2832 5828 2838 5840
rect 2832 5800 3004 5828
rect 2832 5788 2838 5800
rect 2976 5769 3004 5800
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 2961 5763 3019 5769
rect 1719 5732 2912 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 2884 5692 2912 5732
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3418 5760 3424 5772
rect 3007 5732 3424 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 43806 5760 43812 5772
rect 43767 5732 43812 5760
rect 43806 5720 43812 5732
rect 43864 5720 43870 5772
rect 46492 5769 46520 5868
rect 47673 5831 47731 5837
rect 47673 5797 47685 5831
rect 47719 5828 47731 5831
rect 49970 5828 49976 5840
rect 47719 5800 49976 5828
rect 47719 5797 47731 5800
rect 47673 5791 47731 5797
rect 49970 5788 49976 5800
rect 50028 5788 50034 5840
rect 50062 5788 50068 5840
rect 50120 5828 50126 5840
rect 50249 5831 50307 5837
rect 50249 5828 50261 5831
rect 50120 5800 50261 5828
rect 50120 5788 50126 5800
rect 50249 5797 50261 5800
rect 50295 5797 50307 5831
rect 51000 5828 51028 5868
rect 51902 5856 51908 5908
rect 51960 5856 51966 5908
rect 51994 5856 52000 5908
rect 52052 5856 52058 5908
rect 52638 5856 52644 5908
rect 52696 5896 52702 5908
rect 52733 5899 52791 5905
rect 52733 5896 52745 5899
rect 52696 5868 52745 5896
rect 52696 5856 52702 5868
rect 52733 5865 52745 5868
rect 52779 5865 52791 5899
rect 52733 5859 52791 5865
rect 53190 5856 53196 5908
rect 53248 5896 53254 5908
rect 55398 5896 55404 5908
rect 53248 5868 55404 5896
rect 53248 5856 53254 5868
rect 55398 5856 55404 5868
rect 55456 5856 55462 5908
rect 51350 5828 51356 5840
rect 51000 5800 51356 5828
rect 50249 5791 50307 5797
rect 51350 5788 51356 5800
rect 51408 5788 51414 5840
rect 51920 5828 51948 5856
rect 51911 5800 51948 5828
rect 46477 5763 46535 5769
rect 46477 5729 46489 5763
rect 46523 5729 46535 5763
rect 46477 5723 46535 5729
rect 47581 5763 47639 5769
rect 47581 5729 47593 5763
rect 47627 5729 47639 5763
rect 47762 5760 47768 5772
rect 47723 5732 47768 5760
rect 47581 5723 47639 5729
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 2884 5664 4445 5692
rect 1857 5655 1915 5661
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 47596 5692 47624 5723
rect 47762 5720 47768 5732
rect 47820 5720 47826 5772
rect 48406 5760 48412 5772
rect 48367 5732 48412 5760
rect 48406 5720 48412 5732
rect 48464 5720 48470 5772
rect 49050 5760 49056 5772
rect 49011 5732 49056 5760
rect 49050 5720 49056 5732
rect 49108 5720 49114 5772
rect 49602 5720 49608 5772
rect 49660 5760 49666 5772
rect 49697 5763 49755 5769
rect 49697 5760 49709 5763
rect 49660 5732 49709 5760
rect 49660 5720 49666 5732
rect 49697 5729 49709 5732
rect 49743 5729 49755 5763
rect 50154 5760 50160 5772
rect 50115 5732 50160 5760
rect 49697 5723 49755 5729
rect 50154 5720 50160 5732
rect 50212 5720 50218 5772
rect 51911 5769 51939 5800
rect 52012 5769 52040 5856
rect 57974 5828 57980 5840
rect 57935 5800 57980 5828
rect 57974 5788 57980 5800
rect 58032 5788 58038 5840
rect 51767 5763 51825 5769
rect 51767 5729 51779 5763
rect 51813 5729 51825 5763
rect 51767 5723 51825 5729
rect 51886 5763 51944 5769
rect 51886 5729 51898 5763
rect 51932 5729 51944 5763
rect 51886 5723 51944 5729
rect 51986 5763 52044 5769
rect 51986 5729 51998 5763
rect 52032 5729 52044 5763
rect 52178 5760 52184 5772
rect 52139 5732 52184 5760
rect 51986 5723 52044 5729
rect 50890 5692 50896 5704
rect 47596 5664 50896 5692
rect 4433 5655 4491 5661
rect 1872 5624 1900 5655
rect 50890 5652 50896 5664
rect 50948 5652 50954 5704
rect 50982 5652 50988 5704
rect 51040 5692 51046 5704
rect 51626 5692 51632 5704
rect 51040 5664 51632 5692
rect 51040 5652 51046 5664
rect 51626 5652 51632 5664
rect 51684 5652 51690 5704
rect 51797 5692 51825 5723
rect 52178 5720 52184 5732
rect 52236 5720 52242 5772
rect 52914 5760 52920 5772
rect 52875 5732 52920 5760
rect 52914 5720 52920 5732
rect 52972 5720 52978 5772
rect 53009 5763 53067 5769
rect 53009 5729 53021 5763
rect 53055 5729 53067 5763
rect 53282 5760 53288 5772
rect 53243 5732 53288 5760
rect 53009 5723 53067 5729
rect 52086 5692 52092 5704
rect 51797 5664 52092 5692
rect 52086 5652 52092 5664
rect 52144 5652 52150 5704
rect 53024 5692 53052 5723
rect 53282 5720 53288 5732
rect 53340 5720 53346 5772
rect 53742 5760 53748 5772
rect 53703 5732 53748 5760
rect 53742 5720 53748 5732
rect 53800 5720 53806 5772
rect 53837 5763 53895 5769
rect 53837 5729 53849 5763
rect 53883 5760 53895 5763
rect 54018 5760 54024 5772
rect 53883 5732 54024 5760
rect 53883 5729 53895 5732
rect 53837 5723 53895 5729
rect 54018 5720 54024 5732
rect 54076 5720 54082 5772
rect 54481 5763 54539 5769
rect 54481 5729 54493 5763
rect 54527 5760 54539 5763
rect 54754 5760 54760 5772
rect 54527 5732 54760 5760
rect 54527 5729 54539 5732
rect 54481 5723 54539 5729
rect 54496 5692 54524 5723
rect 54754 5720 54760 5732
rect 54812 5720 54818 5772
rect 55585 5763 55643 5769
rect 55585 5729 55597 5763
rect 55631 5760 55643 5763
rect 56318 5760 56324 5772
rect 55631 5732 56324 5760
rect 55631 5729 55643 5732
rect 55585 5723 55643 5729
rect 56318 5720 56324 5732
rect 56376 5720 56382 5772
rect 58158 5760 58164 5772
rect 58119 5732 58164 5760
rect 58158 5720 58164 5732
rect 58216 5720 58222 5772
rect 56686 5692 56692 5704
rect 53024 5664 54524 5692
rect 56647 5664 56692 5692
rect 56686 5652 56692 5664
rect 56744 5652 56750 5704
rect 56778 5652 56784 5704
rect 56836 5692 56842 5704
rect 56873 5695 56931 5701
rect 56873 5692 56885 5695
rect 56836 5664 56885 5692
rect 56836 5652 56842 5664
rect 56873 5661 56885 5664
rect 56919 5661 56931 5695
rect 56873 5655 56931 5661
rect 2777 5627 2835 5633
rect 2777 5624 2789 5627
rect 1872 5596 2789 5624
rect 2777 5593 2789 5596
rect 2823 5593 2835 5627
rect 2777 5587 2835 5593
rect 48038 5584 48044 5636
rect 48096 5624 48102 5636
rect 49513 5627 49571 5633
rect 48096 5596 49464 5624
rect 48096 5584 48102 5596
rect 44361 5559 44419 5565
rect 44361 5525 44373 5559
rect 44407 5556 44419 5559
rect 44634 5556 44640 5568
rect 44407 5528 44640 5556
rect 44407 5525 44419 5528
rect 44361 5519 44419 5525
rect 44634 5516 44640 5528
rect 44692 5516 44698 5568
rect 44910 5556 44916 5568
rect 44871 5528 44916 5556
rect 44910 5516 44916 5528
rect 44968 5556 44974 5568
rect 45281 5559 45339 5565
rect 45281 5556 45293 5559
rect 44968 5528 45293 5556
rect 44968 5516 44974 5528
rect 45281 5525 45293 5528
rect 45327 5525 45339 5559
rect 47118 5556 47124 5568
rect 47079 5528 47124 5556
rect 45281 5519 45339 5525
rect 47118 5516 47124 5528
rect 47176 5516 47182 5568
rect 48130 5516 48136 5568
rect 48188 5556 48194 5568
rect 48225 5559 48283 5565
rect 48225 5556 48237 5559
rect 48188 5528 48237 5556
rect 48188 5516 48194 5528
rect 48225 5525 48237 5528
rect 48271 5525 48283 5559
rect 48225 5519 48283 5525
rect 48869 5559 48927 5565
rect 48869 5525 48881 5559
rect 48915 5556 48927 5559
rect 49326 5556 49332 5568
rect 48915 5528 49332 5556
rect 48915 5525 48927 5528
rect 48869 5519 48927 5525
rect 49326 5516 49332 5528
rect 49384 5516 49390 5568
rect 49436 5556 49464 5596
rect 49513 5593 49525 5627
rect 49559 5624 49571 5627
rect 56502 5624 56508 5636
rect 49559 5596 56508 5624
rect 49559 5593 49571 5596
rect 49513 5587 49571 5593
rect 56502 5584 56508 5596
rect 56560 5584 56566 5636
rect 51166 5556 51172 5568
rect 49436 5528 51172 5556
rect 51166 5516 51172 5528
rect 51224 5516 51230 5568
rect 51534 5556 51540 5568
rect 51495 5528 51540 5556
rect 51534 5516 51540 5528
rect 51592 5516 51598 5568
rect 51902 5516 51908 5568
rect 51960 5556 51966 5568
rect 52638 5556 52644 5568
rect 51960 5528 52644 5556
rect 51960 5516 51966 5528
rect 52638 5516 52644 5528
rect 52696 5516 52702 5568
rect 52822 5516 52828 5568
rect 52880 5556 52886 5568
rect 53193 5559 53251 5565
rect 53193 5556 53205 5559
rect 52880 5528 53205 5556
rect 52880 5516 52886 5528
rect 53193 5525 53205 5528
rect 53239 5556 53251 5559
rect 54294 5556 54300 5568
rect 53239 5528 54300 5556
rect 53239 5525 53251 5528
rect 53193 5519 53251 5525
rect 54294 5516 54300 5528
rect 54352 5556 54358 5568
rect 54573 5559 54631 5565
rect 54573 5556 54585 5559
rect 54352 5528 54585 5556
rect 54352 5516 54358 5528
rect 54573 5525 54585 5528
rect 54619 5525 54631 5559
rect 54573 5519 54631 5525
rect 55677 5559 55735 5565
rect 55677 5525 55689 5559
rect 55723 5556 55735 5559
rect 56410 5556 56416 5568
rect 55723 5528 56416 5556
rect 55723 5525 55735 5528
rect 55677 5519 55735 5525
rect 56410 5516 56416 5528
rect 56468 5516 56474 5568
rect 56594 5516 56600 5568
rect 56652 5556 56658 5568
rect 57057 5559 57115 5565
rect 57057 5556 57069 5559
rect 56652 5528 57069 5556
rect 56652 5516 56658 5528
rect 57057 5525 57069 5528
rect 57103 5525 57115 5559
rect 57057 5519 57115 5525
rect 1104 5466 58880 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 58880 5466
rect 1104 5392 58880 5414
rect 47673 5355 47731 5361
rect 47673 5321 47685 5355
rect 47719 5352 47731 5355
rect 49694 5352 49700 5364
rect 47719 5324 49700 5352
rect 47719 5321 47731 5324
rect 47673 5315 47731 5321
rect 49694 5312 49700 5324
rect 49752 5312 49758 5364
rect 50706 5352 50712 5364
rect 50667 5324 50712 5352
rect 50706 5312 50712 5324
rect 50764 5312 50770 5364
rect 51166 5312 51172 5364
rect 51224 5352 51230 5364
rect 51261 5355 51319 5361
rect 51261 5352 51273 5355
rect 51224 5324 51273 5352
rect 51224 5312 51230 5324
rect 51261 5321 51273 5324
rect 51307 5321 51319 5355
rect 51261 5315 51319 5321
rect 51997 5355 52055 5361
rect 51997 5321 52009 5355
rect 52043 5352 52055 5355
rect 52178 5352 52184 5364
rect 52043 5324 52184 5352
rect 52043 5321 52055 5324
rect 51997 5315 52055 5321
rect 52178 5312 52184 5324
rect 52236 5312 52242 5364
rect 53009 5355 53067 5361
rect 53009 5321 53021 5355
rect 53055 5352 53067 5355
rect 53282 5352 53288 5364
rect 53055 5324 53288 5352
rect 53055 5321 53067 5324
rect 53009 5315 53067 5321
rect 53282 5312 53288 5324
rect 53340 5312 53346 5364
rect 53374 5312 53380 5364
rect 53432 5352 53438 5364
rect 55490 5352 55496 5364
rect 53432 5324 55496 5352
rect 53432 5312 53438 5324
rect 55490 5312 55496 5324
rect 55548 5312 55554 5364
rect 56962 5352 56968 5364
rect 56923 5324 56968 5352
rect 56962 5312 56968 5324
rect 57020 5312 57026 5364
rect 43806 5244 43812 5296
rect 43864 5284 43870 5296
rect 55766 5284 55772 5296
rect 43864 5256 49372 5284
rect 55727 5256 55772 5284
rect 43864 5244 43870 5256
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2866 5216 2872 5228
rect 2087 5188 2872 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2866 5176 2872 5188
rect 2924 5176 2930 5228
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3016 5188 4077 5216
rect 3016 5176 3022 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 44361 5219 44419 5225
rect 44361 5185 44373 5219
rect 44407 5216 44419 5219
rect 49142 5216 49148 5228
rect 44407 5188 49148 5216
rect 44407 5185 44419 5188
rect 44361 5179 44419 5185
rect 49142 5176 49148 5188
rect 49200 5176 49206 5228
rect 49344 5216 49372 5256
rect 55766 5244 55772 5256
rect 55824 5244 55830 5296
rect 57146 5244 57152 5296
rect 57204 5284 57210 5296
rect 57885 5287 57943 5293
rect 57885 5284 57897 5287
rect 57204 5256 57897 5284
rect 57204 5244 57210 5256
rect 57885 5253 57897 5256
rect 57931 5253 57943 5287
rect 57885 5247 57943 5253
rect 49344 5188 49464 5216
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3418 5148 3424 5160
rect 3379 5120 3424 5148
rect 3418 5108 3424 5120
rect 3476 5108 3482 5160
rect 43533 5151 43591 5157
rect 43533 5117 43545 5151
rect 43579 5148 43591 5151
rect 44082 5148 44088 5160
rect 43579 5120 44088 5148
rect 43579 5117 43591 5120
rect 43533 5111 43591 5117
rect 44082 5108 44088 5120
rect 44140 5108 44146 5160
rect 45002 5148 45008 5160
rect 44963 5120 45008 5148
rect 45002 5108 45008 5120
rect 45060 5108 45066 5160
rect 45646 5148 45652 5160
rect 45607 5120 45652 5148
rect 45646 5108 45652 5120
rect 45704 5108 45710 5160
rect 46569 5151 46627 5157
rect 46569 5117 46581 5151
rect 46615 5148 46627 5151
rect 46934 5148 46940 5160
rect 46615 5120 46940 5148
rect 46615 5117 46627 5120
rect 46569 5111 46627 5117
rect 46934 5108 46940 5120
rect 46992 5108 46998 5160
rect 47029 5151 47087 5157
rect 47029 5117 47041 5151
rect 47075 5117 47087 5151
rect 47029 5111 47087 5117
rect 47213 5151 47271 5157
rect 47213 5117 47225 5151
rect 47259 5148 47271 5151
rect 47762 5148 47768 5160
rect 47259 5120 47768 5148
rect 47259 5117 47271 5120
rect 47213 5111 47271 5117
rect 1857 5083 1915 5089
rect 1857 5049 1869 5083
rect 1903 5080 1915 5083
rect 2314 5080 2320 5092
rect 1903 5052 2320 5080
rect 1903 5049 1915 5052
rect 1857 5043 1915 5049
rect 2314 5040 2320 5052
rect 2372 5040 2378 5092
rect 2590 5080 2596 5092
rect 2551 5052 2596 5080
rect 2590 5040 2596 5052
rect 2648 5040 2654 5092
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3237 5015 3295 5021
rect 3237 5012 3249 5015
rect 2832 4984 3249 5012
rect 2832 4972 2838 4984
rect 3237 4981 3249 4984
rect 3283 4981 3295 5015
rect 47044 5012 47072 5111
rect 47762 5108 47768 5120
rect 47820 5108 47826 5160
rect 47854 5108 47860 5160
rect 47912 5148 47918 5160
rect 48314 5148 48320 5160
rect 47912 5120 48320 5148
rect 47912 5108 47918 5120
rect 48314 5108 48320 5120
rect 48372 5108 48378 5160
rect 48774 5108 48780 5160
rect 48832 5148 48838 5160
rect 49234 5148 49240 5160
rect 48832 5120 49240 5148
rect 48832 5108 48838 5120
rect 49234 5108 49240 5120
rect 49292 5148 49298 5160
rect 49329 5151 49387 5157
rect 49329 5148 49341 5151
rect 49292 5120 49341 5148
rect 49292 5108 49298 5120
rect 49329 5117 49341 5120
rect 49375 5117 49387 5151
rect 49436 5148 49464 5188
rect 55306 5176 55312 5228
rect 55364 5216 55370 5228
rect 57701 5219 57759 5225
rect 57701 5216 57713 5219
rect 55364 5188 57713 5216
rect 55364 5176 55370 5188
rect 57701 5185 57713 5188
rect 57747 5185 57759 5219
rect 57701 5179 57759 5185
rect 50154 5148 50160 5160
rect 49436 5120 50160 5148
rect 49329 5111 49387 5117
rect 50154 5108 50160 5120
rect 50212 5108 50218 5160
rect 50706 5108 50712 5160
rect 50764 5148 50770 5160
rect 51169 5151 51227 5157
rect 51169 5148 51181 5151
rect 50764 5120 51181 5148
rect 50764 5108 50770 5120
rect 51169 5117 51181 5120
rect 51215 5117 51227 5151
rect 51902 5148 51908 5160
rect 51863 5120 51908 5148
rect 51169 5111 51227 5117
rect 51902 5108 51908 5120
rect 51960 5108 51966 5160
rect 52086 5148 52092 5160
rect 52047 5120 52092 5148
rect 52086 5108 52092 5120
rect 52144 5108 52150 5160
rect 52914 5148 52920 5160
rect 52875 5120 52920 5148
rect 52914 5108 52920 5120
rect 52972 5108 52978 5160
rect 54018 5108 54024 5160
rect 54076 5157 54082 5160
rect 54076 5148 54085 5157
rect 54202 5148 54208 5160
rect 54076 5120 54121 5148
rect 54163 5120 54208 5148
rect 54076 5111 54085 5120
rect 54076 5108 54082 5111
rect 54202 5108 54208 5120
rect 54260 5108 54266 5160
rect 54386 5108 54392 5160
rect 54444 5148 54450 5160
rect 55401 5151 55459 5157
rect 55401 5148 55413 5151
rect 54444 5120 55413 5148
rect 54444 5108 54450 5120
rect 55401 5117 55413 5120
rect 55447 5117 55459 5151
rect 55401 5111 55459 5117
rect 55490 5108 55496 5160
rect 55548 5148 55554 5160
rect 55585 5151 55643 5157
rect 55585 5148 55597 5151
rect 55548 5120 55597 5148
rect 55548 5108 55554 5120
rect 55585 5117 55597 5120
rect 55631 5117 55643 5151
rect 55585 5111 55643 5117
rect 56873 5151 56931 5157
rect 56873 5117 56885 5151
rect 56919 5148 56931 5151
rect 57054 5148 57060 5160
rect 56919 5120 57060 5148
rect 56919 5117 56931 5120
rect 56873 5111 56931 5117
rect 57054 5108 57060 5120
rect 57112 5108 57118 5160
rect 57517 5151 57575 5157
rect 57517 5117 57529 5151
rect 57563 5117 57575 5151
rect 57517 5111 57575 5117
rect 47121 5083 47179 5089
rect 47121 5049 47133 5083
rect 47167 5080 47179 5083
rect 49596 5083 49654 5089
rect 47167 5052 49556 5080
rect 47167 5049 47179 5052
rect 47121 5043 47179 5049
rect 49418 5012 49424 5024
rect 47044 4984 49424 5012
rect 3237 4975 3295 4981
rect 49418 4972 49424 4984
rect 49476 4972 49482 5024
rect 49528 5012 49556 5052
rect 49596 5049 49608 5083
rect 49642 5080 49654 5083
rect 49970 5080 49976 5092
rect 49642 5052 49976 5080
rect 49642 5049 49654 5052
rect 49596 5043 49654 5049
rect 49970 5040 49976 5052
rect 50028 5040 50034 5092
rect 54757 5083 54815 5089
rect 54757 5049 54769 5083
rect 54803 5080 54815 5083
rect 56502 5080 56508 5092
rect 54803 5052 56508 5080
rect 54803 5049 54815 5052
rect 54757 5043 54815 5049
rect 56502 5040 56508 5052
rect 56560 5040 56566 5092
rect 51074 5012 51080 5024
rect 49528 4984 51080 5012
rect 51074 4972 51080 4984
rect 51132 4972 51138 5024
rect 51166 4972 51172 5024
rect 51224 5012 51230 5024
rect 53374 5012 53380 5024
rect 51224 4984 53380 5012
rect 51224 4972 51230 4984
rect 53374 4972 53380 4984
rect 53432 4972 53438 5024
rect 53466 4972 53472 5024
rect 53524 5012 53530 5024
rect 53834 5012 53840 5024
rect 53524 4984 53840 5012
rect 53524 4972 53530 4984
rect 53834 4972 53840 4984
rect 53892 4972 53898 5024
rect 54110 5012 54116 5024
rect 54071 4984 54116 5012
rect 54110 4972 54116 4984
rect 54168 4972 54174 5024
rect 54849 5015 54907 5021
rect 54849 4981 54861 5015
rect 54895 5012 54907 5015
rect 56226 5012 56232 5024
rect 54895 4984 56232 5012
rect 54895 4981 54907 4984
rect 54849 4975 54907 4981
rect 56226 4972 56232 4984
rect 56284 4972 56290 5024
rect 57330 5012 57336 5024
rect 57291 4984 57336 5012
rect 57330 4972 57336 4984
rect 57388 5012 57394 5024
rect 57532 5012 57560 5111
rect 57388 4984 57560 5012
rect 57388 4972 57394 4984
rect 1104 4922 58880 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 50326 4922
rect 50378 4870 50390 4922
rect 50442 4870 50454 4922
rect 50506 4870 50518 4922
rect 50570 4870 58880 4922
rect 1104 4848 58880 4870
rect 2590 4808 2596 4820
rect 2551 4780 2596 4808
rect 2590 4768 2596 4780
rect 2648 4768 2654 4820
rect 45278 4768 45284 4820
rect 45336 4808 45342 4820
rect 47762 4808 47768 4820
rect 45336 4780 47768 4808
rect 45336 4768 45342 4780
rect 47762 4768 47768 4780
rect 47820 4768 47826 4820
rect 47946 4768 47952 4820
rect 48004 4808 48010 4820
rect 48777 4811 48835 4817
rect 48777 4808 48789 4811
rect 48004 4780 48789 4808
rect 48004 4768 48010 4780
rect 48777 4777 48789 4780
rect 48823 4808 48835 4811
rect 49050 4808 49056 4820
rect 48823 4780 49056 4808
rect 48823 4777 48835 4780
rect 48777 4771 48835 4777
rect 49050 4768 49056 4780
rect 49108 4768 49114 4820
rect 49970 4808 49976 4820
rect 49931 4780 49976 4808
rect 49970 4768 49976 4780
rect 50028 4768 50034 4820
rect 50154 4768 50160 4820
rect 50212 4808 50218 4820
rect 55214 4808 55220 4820
rect 50212 4780 55220 4808
rect 50212 4768 50218 4780
rect 55214 4768 55220 4780
rect 55272 4768 55278 4820
rect 47854 4740 47860 4752
rect 46860 4712 47860 4740
rect 2133 4675 2191 4681
rect 2133 4641 2145 4675
rect 2179 4672 2191 4675
rect 2774 4672 2780 4684
rect 2179 4644 2780 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 3237 4675 3295 4681
rect 3237 4641 3249 4675
rect 3283 4672 3295 4675
rect 3418 4672 3424 4684
rect 3283 4644 3424 4672
rect 3283 4641 3295 4644
rect 3237 4635 3295 4641
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 38102 4672 38108 4684
rect 38063 4644 38108 4672
rect 38102 4632 38108 4644
rect 38160 4632 38166 4684
rect 46566 4632 46572 4684
rect 46624 4672 46630 4684
rect 46860 4681 46888 4712
rect 47854 4700 47860 4712
rect 47912 4700 47918 4752
rect 50246 4700 50252 4752
rect 50304 4740 50310 4752
rect 50304 4712 51488 4740
rect 50304 4700 50310 4712
rect 46845 4675 46903 4681
rect 46845 4672 46857 4675
rect 46624 4644 46857 4672
rect 46624 4632 46630 4644
rect 46845 4641 46857 4644
rect 46891 4641 46903 4675
rect 46845 4635 46903 4641
rect 47302 4632 47308 4684
rect 47360 4672 47366 4684
rect 47489 4675 47547 4681
rect 47489 4672 47501 4675
rect 47360 4644 47501 4672
rect 47360 4632 47366 4644
rect 47489 4641 47501 4644
rect 47535 4672 47547 4675
rect 47946 4672 47952 4684
rect 47535 4644 47952 4672
rect 47535 4641 47547 4644
rect 47489 4635 47547 4641
rect 47946 4632 47952 4644
rect 48004 4672 48010 4684
rect 48133 4675 48191 4681
rect 48133 4672 48145 4675
rect 48004 4644 48145 4672
rect 48004 4632 48010 4644
rect 48133 4641 48145 4644
rect 48179 4641 48191 4675
rect 48133 4635 48191 4641
rect 48593 4675 48651 4681
rect 48593 4641 48605 4675
rect 48639 4672 48651 4675
rect 48774 4672 48780 4684
rect 48639 4644 48780 4672
rect 48639 4641 48651 4644
rect 48593 4635 48651 4641
rect 48774 4632 48780 4644
rect 48832 4632 48838 4684
rect 49421 4675 49479 4681
rect 49421 4641 49433 4675
rect 49467 4672 49479 4675
rect 49602 4672 49608 4684
rect 49467 4644 49608 4672
rect 49467 4641 49479 4644
rect 49421 4635 49479 4641
rect 49602 4632 49608 4644
rect 49660 4632 49666 4684
rect 49878 4672 49884 4684
rect 49839 4644 49884 4672
rect 49878 4632 49884 4644
rect 49936 4632 49942 4684
rect 50062 4672 50068 4684
rect 50023 4644 50068 4672
rect 50062 4632 50068 4644
rect 50120 4632 50126 4684
rect 51460 4672 51488 4712
rect 51534 4700 51540 4752
rect 51592 4740 51598 4752
rect 51782 4743 51840 4749
rect 51782 4740 51794 4743
rect 51592 4712 51794 4740
rect 51592 4700 51598 4712
rect 51782 4709 51794 4712
rect 51828 4709 51840 4743
rect 51782 4703 51840 4709
rect 53644 4743 53702 4749
rect 53644 4709 53656 4743
rect 53690 4740 53702 4743
rect 54110 4740 54116 4752
rect 53690 4712 54116 4740
rect 53690 4709 53702 4712
rect 53644 4703 53702 4709
rect 54110 4700 54116 4712
rect 54168 4700 54174 4752
rect 56873 4743 56931 4749
rect 56873 4709 56885 4743
rect 56919 4740 56931 4743
rect 57146 4740 57152 4752
rect 56919 4712 57152 4740
rect 56919 4709 56931 4712
rect 56873 4703 56931 4709
rect 57146 4700 57152 4712
rect 57204 4700 57210 4752
rect 55309 4675 55367 4681
rect 55309 4672 55321 4675
rect 51460 4644 55321 4672
rect 55309 4641 55321 4644
rect 55355 4641 55367 4675
rect 55309 4635 55367 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 3326 4604 3332 4616
rect 1995 4576 3332 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 50706 4604 50712 4616
rect 48056 4576 50712 4604
rect 46661 4539 46719 4545
rect 46661 4505 46673 4539
rect 46707 4536 46719 4539
rect 47394 4536 47400 4548
rect 46707 4508 47400 4536
rect 46707 4505 46719 4508
rect 46661 4499 46719 4505
rect 47394 4496 47400 4508
rect 47452 4496 47458 4548
rect 47762 4496 47768 4548
rect 47820 4536 47826 4548
rect 48056 4536 48084 4576
rect 50706 4564 50712 4576
rect 50764 4564 50770 4616
rect 50890 4564 50896 4616
rect 50948 4604 50954 4616
rect 51537 4607 51595 4613
rect 51537 4604 51549 4607
rect 50948 4576 51549 4604
rect 50948 4564 50954 4576
rect 51537 4573 51549 4576
rect 51583 4573 51595 4607
rect 53374 4604 53380 4616
rect 53335 4576 53380 4604
rect 51537 4567 51595 4573
rect 53374 4564 53380 4576
rect 53432 4564 53438 4616
rect 57238 4564 57244 4616
rect 57296 4604 57302 4616
rect 57333 4607 57391 4613
rect 57333 4604 57345 4607
rect 57296 4576 57345 4604
rect 57296 4564 57302 4576
rect 57333 4573 57345 4576
rect 57379 4604 57391 4607
rect 57517 4607 57575 4613
rect 57517 4604 57529 4607
rect 57379 4576 57529 4604
rect 57379 4573 57391 4576
rect 57333 4567 57391 4573
rect 57517 4573 57529 4576
rect 57563 4573 57575 4607
rect 57517 4567 57575 4573
rect 57701 4607 57759 4613
rect 57701 4573 57713 4607
rect 57747 4573 57759 4607
rect 57701 4567 57759 4573
rect 47820 4508 48084 4536
rect 47820 4496 47826 4508
rect 48130 4496 48136 4548
rect 48188 4536 48194 4548
rect 51442 4536 51448 4548
rect 48188 4508 51448 4536
rect 48188 4496 48194 4508
rect 51442 4496 51448 4508
rect 51500 4496 51506 4548
rect 52914 4536 52920 4548
rect 52875 4508 52920 4536
rect 52914 4496 52920 4508
rect 52972 4496 52978 4548
rect 55493 4539 55551 4545
rect 55493 4536 55505 4539
rect 54312 4508 55505 4536
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4468 4491 4471
rect 4614 4468 4620 4480
rect 4479 4440 4620 4468
rect 4479 4437 4491 4440
rect 4433 4431 4491 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 34514 4468 34520 4480
rect 34475 4440 34520 4468
rect 34514 4428 34520 4440
rect 34572 4428 34578 4480
rect 35894 4428 35900 4480
rect 35952 4468 35958 4480
rect 35952 4440 35997 4468
rect 35952 4428 35958 4440
rect 36262 4428 36268 4480
rect 36320 4468 36326 4480
rect 36725 4471 36783 4477
rect 36725 4468 36737 4471
rect 36320 4440 36737 4468
rect 36320 4428 36326 4440
rect 36725 4437 36737 4440
rect 36771 4437 36783 4471
rect 36725 4431 36783 4437
rect 37921 4471 37979 4477
rect 37921 4437 37933 4471
rect 37967 4468 37979 4471
rect 38470 4468 38476 4480
rect 37967 4440 38476 4468
rect 37967 4437 37979 4440
rect 37921 4431 37979 4437
rect 38470 4428 38476 4440
rect 38528 4428 38534 4480
rect 38746 4468 38752 4480
rect 38707 4440 38752 4468
rect 38746 4428 38752 4440
rect 38804 4428 38810 4480
rect 42794 4468 42800 4480
rect 42755 4440 42800 4468
rect 42794 4428 42800 4440
rect 42852 4428 42858 4480
rect 43530 4468 43536 4480
rect 43491 4440 43536 4468
rect 43530 4428 43536 4440
rect 43588 4428 43594 4480
rect 44174 4468 44180 4480
rect 44135 4440 44180 4468
rect 44174 4428 44180 4440
rect 44232 4428 44238 4480
rect 45094 4468 45100 4480
rect 45055 4440 45100 4468
rect 45094 4428 45100 4440
rect 45152 4428 45158 4480
rect 47305 4471 47363 4477
rect 47305 4437 47317 4471
rect 47351 4468 47363 4471
rect 47670 4468 47676 4480
rect 47351 4440 47676 4468
rect 47351 4437 47363 4440
rect 47305 4431 47363 4437
rect 47670 4428 47676 4440
rect 47728 4428 47734 4480
rect 47946 4468 47952 4480
rect 47907 4440 47952 4468
rect 47946 4428 47952 4440
rect 48004 4428 48010 4480
rect 49234 4468 49240 4480
rect 49195 4440 49240 4468
rect 49234 4428 49240 4440
rect 49292 4428 49298 4480
rect 49786 4428 49792 4480
rect 49844 4468 49850 4480
rect 50890 4468 50896 4480
rect 49844 4440 50896 4468
rect 49844 4428 49850 4440
rect 50890 4428 50896 4440
rect 50948 4428 50954 4480
rect 51074 4428 51080 4480
rect 51132 4468 51138 4480
rect 54312 4468 54340 4508
rect 55493 4505 55505 4508
rect 55539 4505 55551 4539
rect 55493 4499 55551 4505
rect 55582 4496 55588 4548
rect 55640 4536 55646 4548
rect 57716 4536 57744 4567
rect 55640 4508 57744 4536
rect 55640 4496 55646 4508
rect 54754 4468 54760 4480
rect 51132 4440 54340 4468
rect 54715 4440 54760 4468
rect 51132 4428 51138 4440
rect 54754 4428 54760 4440
rect 54812 4428 54818 4480
rect 56962 4468 56968 4480
rect 56923 4440 56968 4468
rect 56962 4428 56968 4440
rect 57020 4428 57026 4480
rect 57974 4468 57980 4480
rect 57935 4440 57980 4468
rect 57974 4428 57980 4440
rect 58032 4428 58038 4480
rect 1104 4378 58880 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 58880 4378
rect 1104 4304 58880 4326
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 44634 4224 44640 4276
rect 44692 4264 44698 4276
rect 52181 4267 52239 4273
rect 44692 4236 52132 4264
rect 44692 4224 44698 4236
rect 39761 4199 39819 4205
rect 39761 4165 39773 4199
rect 39807 4196 39819 4199
rect 40034 4196 40040 4208
rect 39807 4168 40040 4196
rect 39807 4165 39819 4168
rect 39761 4159 39819 4165
rect 40034 4156 40040 4168
rect 40092 4156 40098 4208
rect 41141 4199 41199 4205
rect 41141 4165 41153 4199
rect 41187 4196 41199 4199
rect 41598 4196 41604 4208
rect 41187 4168 41604 4196
rect 41187 4165 41199 4168
rect 41141 4159 41199 4165
rect 41598 4156 41604 4168
rect 41656 4156 41662 4208
rect 41969 4199 42027 4205
rect 41969 4165 41981 4199
rect 42015 4196 42027 4199
rect 42702 4196 42708 4208
rect 42015 4168 42708 4196
rect 42015 4165 42027 4168
rect 41969 4159 42027 4165
rect 42702 4156 42708 4168
rect 42760 4156 42766 4208
rect 46382 4196 46388 4208
rect 43364 4168 46388 4196
rect 43364 4140 43392 4168
rect 46382 4156 46388 4168
rect 46440 4156 46446 4208
rect 46566 4196 46572 4208
rect 46527 4168 46572 4196
rect 46566 4156 46572 4168
rect 46624 4156 46630 4208
rect 47029 4199 47087 4205
rect 47029 4165 47041 4199
rect 47075 4165 47087 4199
rect 47029 4159 47087 4165
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 3050 4128 3056 4140
rect 1811 4100 3056 4128
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 3050 4088 3056 4100
rect 3108 4088 3114 4140
rect 4614 4128 4620 4140
rect 3160 4100 4620 4128
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4060 1639 4063
rect 3160 4060 3188 4100
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 37182 4128 37188 4140
rect 36832 4100 37188 4128
rect 1627 4032 3188 4060
rect 3605 4063 3663 4069
rect 1627 4029 1639 4032
rect 1581 4023 1639 4029
rect 3605 4029 3617 4063
rect 3651 4060 3663 4063
rect 3694 4060 3700 4072
rect 3651 4032 3700 4060
rect 3651 4029 3663 4032
rect 3605 4023 3663 4029
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 4154 4020 4160 4072
rect 4212 4060 4218 4072
rect 4249 4063 4307 4069
rect 4249 4060 4261 4063
rect 4212 4032 4261 4060
rect 4212 4020 4218 4032
rect 4249 4029 4261 4032
rect 4295 4029 4307 4063
rect 4249 4023 4307 4029
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 33321 4063 33379 4069
rect 33321 4029 33333 4063
rect 33367 4060 33379 4063
rect 33410 4060 33416 4072
rect 33367 4032 33416 4060
rect 33367 4029 33379 4032
rect 33321 4023 33379 4029
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 2777 3995 2835 4001
rect 2777 3992 2789 3995
rect 2271 3964 2789 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 2777 3961 2789 3964
rect 2823 3961 2835 3995
rect 4724 3992 4752 4023
rect 33410 4020 33416 4032
rect 33468 4020 33474 4072
rect 33962 4060 33968 4072
rect 33923 4032 33968 4060
rect 33962 4020 33968 4032
rect 34020 4020 34026 4072
rect 36832 4069 36860 4100
rect 37182 4088 37188 4100
rect 37240 4128 37246 4140
rect 43346 4128 43352 4140
rect 37240 4100 43352 4128
rect 37240 4088 37246 4100
rect 43346 4088 43352 4100
rect 43404 4088 43410 4140
rect 46584 4128 46612 4156
rect 45940 4100 46612 4128
rect 47044 4128 47072 4159
rect 47486 4156 47492 4208
rect 47544 4196 47550 4208
rect 50246 4196 50252 4208
rect 47544 4168 50252 4196
rect 47544 4156 47550 4168
rect 50246 4156 50252 4168
rect 50304 4156 50310 4208
rect 52104 4196 52132 4236
rect 52181 4233 52193 4267
rect 52227 4264 52239 4267
rect 55582 4264 55588 4276
rect 52227 4236 55588 4264
rect 52227 4233 52239 4236
rect 52181 4227 52239 4233
rect 55582 4224 55588 4236
rect 55640 4224 55646 4276
rect 56502 4224 56508 4276
rect 56560 4264 56566 4276
rect 56873 4267 56931 4273
rect 56873 4264 56885 4267
rect 56560 4236 56885 4264
rect 56560 4224 56566 4236
rect 56873 4233 56885 4236
rect 56919 4233 56931 4267
rect 56873 4227 56931 4233
rect 57330 4196 57336 4208
rect 52104 4168 57336 4196
rect 57330 4156 57336 4168
rect 57388 4156 57394 4208
rect 49510 4128 49516 4140
rect 47044 4100 49516 4128
rect 34609 4063 34667 4069
rect 34609 4029 34621 4063
rect 34655 4060 34667 4063
rect 35713 4063 35771 4069
rect 35713 4060 35725 4063
rect 34655 4032 35725 4060
rect 34655 4029 34667 4032
rect 34609 4023 34667 4029
rect 35713 4029 35725 4032
rect 35759 4060 35771 4063
rect 36357 4063 36415 4069
rect 36357 4060 36369 4063
rect 35759 4032 36369 4060
rect 35759 4029 35771 4032
rect 35713 4023 35771 4029
rect 36357 4029 36369 4032
rect 36403 4029 36415 4063
rect 36357 4023 36415 4029
rect 36817 4063 36875 4069
rect 36817 4029 36829 4063
rect 36863 4029 36875 4063
rect 36817 4023 36875 4029
rect 2777 3955 2835 3961
rect 2884 3964 4752 3992
rect 33428 3992 33456 4020
rect 34624 3992 34652 4023
rect 33428 3964 34652 3992
rect 36372 3992 36400 4023
rect 37366 4020 37372 4072
rect 37424 4060 37430 4072
rect 38102 4060 38108 4072
rect 37424 4032 38108 4060
rect 37424 4020 37430 4032
rect 38102 4020 38108 4032
rect 38160 4060 38166 4072
rect 38473 4063 38531 4069
rect 38473 4060 38485 4063
rect 38160 4032 38485 4060
rect 38160 4020 38166 4032
rect 38473 4029 38485 4032
rect 38519 4029 38531 4063
rect 39114 4060 39120 4072
rect 39075 4032 39120 4060
rect 38473 4023 38531 4029
rect 39114 4020 39120 4032
rect 39172 4020 39178 4072
rect 40494 4060 40500 4072
rect 40455 4032 40500 4060
rect 40494 4020 40500 4032
rect 40552 4020 40558 4072
rect 42613 4063 42671 4069
rect 42613 4029 42625 4063
rect 42659 4060 42671 4063
rect 44177 4063 44235 4069
rect 44177 4060 44189 4063
rect 42659 4032 44189 4060
rect 42659 4029 42671 4032
rect 42613 4023 42671 4029
rect 44177 4029 44189 4032
rect 44223 4060 44235 4063
rect 44634 4060 44640 4072
rect 44223 4032 44640 4060
rect 44223 4029 44235 4032
rect 44177 4023 44235 4029
rect 44634 4020 44640 4032
rect 44692 4060 44698 4072
rect 45281 4063 45339 4069
rect 45281 4060 45293 4063
rect 44692 4032 45293 4060
rect 44692 4020 44698 4032
rect 45281 4029 45293 4032
rect 45327 4029 45339 4063
rect 45281 4023 45339 4029
rect 45738 4020 45744 4072
rect 45796 4060 45802 4072
rect 45940 4069 45968 4100
rect 49510 4088 49516 4100
rect 49568 4088 49574 4140
rect 50338 4088 50344 4140
rect 50396 4128 50402 4140
rect 56321 4131 56379 4137
rect 56321 4128 56333 4131
rect 50396 4100 56333 4128
rect 50396 4088 50402 4100
rect 56321 4097 56333 4100
rect 56367 4128 56379 4131
rect 56505 4131 56563 4137
rect 56505 4128 56517 4131
rect 56367 4100 56517 4128
rect 56367 4097 56379 4100
rect 56321 4091 56379 4097
rect 56505 4097 56517 4100
rect 56551 4097 56563 4131
rect 56686 4128 56692 4140
rect 56647 4100 56692 4128
rect 56505 4091 56563 4097
rect 56686 4088 56692 4100
rect 56744 4088 56750 4140
rect 45925 4063 45983 4069
rect 45925 4060 45937 4063
rect 45796 4032 45937 4060
rect 45796 4020 45802 4032
rect 45925 4029 45937 4032
rect 45971 4029 45983 4063
rect 46382 4060 46388 4072
rect 46343 4032 46388 4060
rect 45925 4023 45983 4029
rect 46382 4020 46388 4032
rect 46440 4020 46446 4072
rect 46474 4020 46480 4072
rect 46532 4060 46538 4072
rect 47213 4063 47271 4069
rect 46532 4032 47164 4060
rect 46532 4020 46538 4032
rect 47026 3992 47032 4004
rect 36372 3964 37044 3992
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 2884 3924 2912 3964
rect 1452 3896 2912 3924
rect 1452 3884 1458 3896
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 3016 3896 3433 3924
rect 3016 3884 3022 3896
rect 3421 3893 3433 3896
rect 3467 3893 3479 3927
rect 3421 3887 3479 3893
rect 33137 3927 33195 3933
rect 33137 3893 33149 3927
rect 33183 3924 33195 3927
rect 33778 3924 33784 3936
rect 33183 3896 33784 3924
rect 33183 3893 33195 3896
rect 33137 3887 33195 3893
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 34425 3927 34483 3933
rect 34425 3893 34437 3927
rect 34471 3924 34483 3927
rect 34790 3924 34796 3936
rect 34471 3896 34796 3924
rect 34471 3893 34483 3896
rect 34425 3887 34483 3893
rect 34790 3884 34796 3896
rect 34848 3884 34854 3936
rect 35526 3924 35532 3936
rect 35487 3896 35532 3924
rect 35526 3884 35532 3896
rect 35584 3884 35590 3936
rect 36170 3924 36176 3936
rect 36131 3896 36176 3924
rect 36170 3884 36176 3896
rect 36228 3884 36234 3936
rect 37016 3933 37044 3964
rect 45756 3964 47032 3992
rect 37001 3927 37059 3933
rect 37001 3893 37013 3927
rect 37047 3893 37059 3927
rect 37001 3887 37059 3893
rect 38289 3927 38347 3933
rect 38289 3893 38301 3927
rect 38335 3924 38347 3927
rect 39022 3924 39028 3936
rect 38335 3896 39028 3924
rect 38335 3893 38347 3896
rect 38289 3887 38347 3893
rect 39022 3884 39028 3896
rect 39080 3884 39086 3936
rect 42429 3927 42487 3933
rect 42429 3893 42441 3927
rect 42475 3924 42487 3927
rect 42886 3924 42892 3936
rect 42475 3896 42892 3924
rect 42475 3893 42487 3896
rect 42429 3887 42487 3893
rect 42886 3884 42892 3896
rect 42944 3884 42950 3936
rect 43993 3927 44051 3933
rect 43993 3893 44005 3927
rect 44039 3924 44051 3927
rect 44358 3924 44364 3936
rect 44039 3896 44364 3924
rect 44039 3893 44051 3896
rect 43993 3887 44051 3893
rect 44358 3884 44364 3896
rect 44416 3884 44422 3936
rect 45097 3927 45155 3933
rect 45097 3893 45109 3927
rect 45143 3924 45155 3927
rect 45462 3924 45468 3936
rect 45143 3896 45468 3924
rect 45143 3893 45155 3896
rect 45097 3887 45155 3893
rect 45462 3884 45468 3896
rect 45520 3884 45526 3936
rect 45756 3933 45784 3964
rect 47026 3952 47032 3964
rect 47084 3952 47090 4004
rect 47136 3992 47164 4032
rect 47213 4029 47225 4063
rect 47259 4060 47271 4063
rect 47302 4060 47308 4072
rect 47259 4032 47308 4060
rect 47259 4029 47271 4032
rect 47213 4023 47271 4029
rect 47302 4020 47308 4032
rect 47360 4060 47366 4072
rect 47857 4063 47915 4069
rect 47857 4060 47869 4063
rect 47360 4032 47869 4060
rect 47360 4020 47366 4032
rect 47857 4029 47869 4032
rect 47903 4029 47915 4063
rect 47857 4023 47915 4029
rect 49145 4063 49203 4069
rect 49145 4029 49157 4063
rect 49191 4060 49203 4063
rect 49602 4060 49608 4072
rect 49191 4032 49608 4060
rect 49191 4029 49203 4032
rect 49145 4023 49203 4029
rect 49602 4020 49608 4032
rect 49660 4060 49666 4072
rect 49789 4063 49847 4069
rect 49789 4060 49801 4063
rect 49660 4032 49801 4060
rect 49660 4020 49666 4032
rect 49789 4029 49801 4032
rect 49835 4060 49847 4063
rect 50433 4063 50491 4069
rect 50433 4060 50445 4063
rect 49835 4032 50445 4060
rect 49835 4029 49847 4032
rect 49789 4023 49847 4029
rect 50433 4029 50445 4032
rect 50479 4029 50491 4063
rect 50890 4060 50896 4072
rect 50851 4032 50896 4060
rect 50433 4023 50491 4029
rect 50338 3992 50344 4004
rect 47136 3964 50344 3992
rect 50338 3952 50344 3964
rect 50396 3952 50402 4004
rect 50448 3992 50476 4023
rect 50890 4020 50896 4032
rect 50948 4020 50954 4072
rect 51718 4020 51724 4072
rect 51776 4060 51782 4072
rect 52365 4063 52423 4069
rect 51776 4032 51821 4060
rect 51776 4020 51782 4032
rect 52365 4029 52377 4063
rect 52411 4060 52423 4063
rect 52730 4060 52736 4072
rect 52411 4032 52736 4060
rect 52411 4029 52423 4032
rect 52365 4023 52423 4029
rect 52730 4020 52736 4032
rect 52788 4020 52794 4072
rect 52917 4063 52975 4069
rect 52917 4029 52929 4063
rect 52963 4060 52975 4063
rect 55861 4063 55919 4069
rect 52963 4032 55812 4060
rect 52963 4029 52975 4032
rect 52917 4023 52975 4029
rect 50448 3964 51120 3992
rect 45741 3927 45799 3933
rect 45741 3893 45753 3927
rect 45787 3893 45799 3927
rect 45741 3887 45799 3893
rect 47673 3927 47731 3933
rect 47673 3893 47685 3927
rect 47719 3924 47731 3927
rect 48130 3924 48136 3936
rect 47719 3896 48136 3924
rect 47719 3893 47731 3896
rect 47673 3887 47731 3893
rect 48130 3884 48136 3896
rect 48188 3884 48194 3936
rect 48961 3927 49019 3933
rect 48961 3893 48973 3927
rect 49007 3924 49019 3927
rect 49418 3924 49424 3936
rect 49007 3896 49424 3924
rect 49007 3893 49019 3896
rect 48961 3887 49019 3893
rect 49418 3884 49424 3896
rect 49476 3884 49482 3936
rect 49605 3927 49663 3933
rect 49605 3893 49617 3927
rect 49651 3924 49663 3927
rect 50062 3924 50068 3936
rect 49651 3896 50068 3924
rect 49651 3893 49663 3896
rect 49605 3887 49663 3893
rect 50062 3884 50068 3896
rect 50120 3884 50126 3936
rect 50249 3927 50307 3933
rect 50249 3893 50261 3927
rect 50295 3924 50307 3927
rect 50982 3924 50988 3936
rect 50295 3896 50988 3924
rect 50295 3893 50307 3896
rect 50249 3887 50307 3893
rect 50982 3884 50988 3896
rect 51040 3884 51046 3936
rect 51092 3933 51120 3964
rect 53098 3952 53104 4004
rect 53156 3992 53162 4004
rect 54389 3995 54447 4001
rect 53156 3964 53201 3992
rect 53156 3952 53162 3964
rect 54389 3961 54401 3995
rect 54435 3992 54447 3995
rect 55030 3992 55036 4004
rect 54435 3964 55036 3992
rect 54435 3961 54447 3964
rect 54389 3955 54447 3961
rect 55030 3952 55036 3964
rect 55088 3952 55094 4004
rect 55125 3995 55183 4001
rect 55125 3961 55137 3995
rect 55171 3992 55183 3995
rect 55582 3992 55588 4004
rect 55171 3964 55588 3992
rect 55171 3961 55183 3964
rect 55125 3955 55183 3961
rect 55582 3952 55588 3964
rect 55640 3952 55646 4004
rect 51077 3927 51135 3933
rect 51077 3893 51089 3927
rect 51123 3893 51135 3927
rect 51077 3887 51135 3893
rect 51537 3927 51595 3933
rect 51537 3893 51549 3927
rect 51583 3924 51595 3927
rect 54202 3924 54208 3936
rect 51583 3896 54208 3924
rect 51583 3893 51595 3896
rect 51537 3887 51595 3893
rect 54202 3884 54208 3896
rect 54260 3884 54266 3936
rect 54478 3924 54484 3936
rect 54439 3896 54484 3924
rect 54478 3884 54484 3896
rect 54536 3884 54542 3936
rect 55217 3927 55275 3933
rect 55217 3893 55229 3927
rect 55263 3924 55275 3927
rect 55674 3924 55680 3936
rect 55263 3896 55680 3924
rect 55263 3893 55275 3896
rect 55217 3887 55275 3893
rect 55674 3884 55680 3896
rect 55732 3884 55738 3936
rect 55784 3924 55812 4032
rect 55861 4029 55873 4063
rect 55907 4060 55919 4063
rect 57974 4060 57980 4072
rect 55907 4032 56456 4060
rect 57935 4032 57980 4060
rect 55907 4029 55919 4032
rect 55861 4023 55919 4029
rect 56042 3992 56048 4004
rect 56003 3964 56048 3992
rect 56042 3952 56048 3964
rect 56100 3952 56106 4004
rect 56428 3992 56456 4032
rect 57974 4020 57980 4032
rect 58032 4020 58038 4072
rect 56594 3992 56600 4004
rect 56428 3964 56600 3992
rect 56594 3952 56600 3964
rect 56652 3952 56658 4004
rect 58158 3992 58164 4004
rect 58119 3964 58164 3992
rect 58158 3952 58164 3964
rect 58216 3952 58222 4004
rect 57238 3924 57244 3936
rect 55784 3896 57244 3924
rect 57238 3884 57244 3896
rect 57296 3884 57302 3936
rect 1104 3834 58880 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 50326 3834
rect 50378 3782 50390 3834
rect 50442 3782 50454 3834
rect 50506 3782 50518 3834
rect 50570 3782 58880 3834
rect 1104 3760 58880 3782
rect 44453 3723 44511 3729
rect 44453 3689 44465 3723
rect 44499 3720 44511 3723
rect 45554 3720 45560 3732
rect 44499 3692 45560 3720
rect 44499 3689 44511 3692
rect 44453 3683 44511 3689
rect 45554 3680 45560 3692
rect 45612 3680 45618 3732
rect 47026 3680 47032 3732
rect 47084 3720 47090 3732
rect 47210 3720 47216 3732
rect 47084 3692 47216 3720
rect 47084 3680 47090 3692
rect 47210 3680 47216 3692
rect 47268 3680 47274 3732
rect 48038 3680 48044 3732
rect 48096 3720 48102 3732
rect 48096 3692 57744 3720
rect 48096 3680 48102 3692
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 1728 3624 41414 3652
rect 1728 3612 1734 3624
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2866 3584 2872 3596
rect 1995 3556 2872 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 3142 3584 3148 3596
rect 3103 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 3970 3516 3976 3528
rect 2179 3488 3976 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 2314 3448 2320 3460
rect 2275 3420 2320 3448
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 5552 3448 5580 3547
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 6181 3587 6239 3593
rect 6181 3584 6193 3587
rect 6144 3556 6193 3584
rect 6144 3544 6150 3556
rect 6181 3553 6193 3556
rect 6227 3553 6239 3587
rect 28534 3584 28540 3596
rect 28495 3556 28540 3584
rect 6181 3547 6239 3553
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 29365 3587 29423 3593
rect 29365 3553 29377 3587
rect 29411 3584 29423 3587
rect 29454 3584 29460 3596
rect 29411 3556 29460 3584
rect 29411 3553 29423 3556
rect 29365 3547 29423 3553
rect 29454 3544 29460 3556
rect 29512 3544 29518 3596
rect 30745 3587 30803 3593
rect 30745 3553 30757 3587
rect 30791 3584 30803 3587
rect 31294 3584 31300 3596
rect 30791 3556 31300 3584
rect 30791 3553 30803 3556
rect 30745 3547 30803 3553
rect 31294 3544 31300 3556
rect 31352 3544 31358 3596
rect 33318 3584 33324 3596
rect 33279 3556 33324 3584
rect 33318 3544 33324 3556
rect 33376 3544 33382 3596
rect 34238 3584 34244 3596
rect 34199 3556 34244 3584
rect 34238 3544 34244 3556
rect 34296 3544 34302 3596
rect 35802 3584 35808 3596
rect 35763 3556 35808 3584
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 37090 3584 37096 3596
rect 37051 3556 37096 3584
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 38013 3587 38071 3593
rect 38013 3553 38025 3587
rect 38059 3584 38071 3587
rect 38654 3584 38660 3596
rect 38059 3556 38660 3584
rect 38059 3553 38071 3556
rect 38013 3547 38071 3553
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 38930 3584 38936 3596
rect 38891 3556 38936 3584
rect 38930 3544 38936 3556
rect 38988 3544 38994 3596
rect 39758 3584 39764 3596
rect 39719 3556 39764 3584
rect 39758 3544 39764 3556
rect 39816 3584 39822 3596
rect 41141 3587 41199 3593
rect 41141 3584 41153 3587
rect 39816 3556 41153 3584
rect 39816 3544 39822 3556
rect 41141 3553 41153 3556
rect 41187 3553 41199 3587
rect 41141 3547 41199 3553
rect 2464 3420 5580 3448
rect 41386 3448 41414 3624
rect 46382 3612 46388 3664
rect 46440 3652 46446 3664
rect 48774 3652 48780 3664
rect 46440 3624 48780 3652
rect 46440 3612 46446 3624
rect 48774 3612 48780 3624
rect 48832 3652 48838 3664
rect 50525 3655 50583 3661
rect 50525 3652 50537 3655
rect 48832 3624 50537 3652
rect 48832 3612 48838 3624
rect 50525 3621 50537 3624
rect 50571 3621 50583 3655
rect 50525 3615 50583 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52362 3652 52368 3664
rect 51500 3624 52368 3652
rect 51500 3612 51506 3624
rect 52362 3612 52368 3624
rect 52420 3612 52426 3664
rect 52454 3612 52460 3664
rect 52512 3652 52518 3664
rect 55585 3655 55643 3661
rect 52512 3624 55343 3652
rect 52512 3612 52518 3624
rect 42153 3587 42211 3593
rect 42153 3553 42165 3587
rect 42199 3553 42211 3587
rect 42153 3547 42211 3553
rect 42705 3587 42763 3593
rect 42705 3553 42717 3587
rect 42751 3584 42763 3587
rect 43070 3584 43076 3596
rect 42751 3556 43076 3584
rect 42751 3553 42763 3556
rect 42705 3547 42763 3553
rect 42168 3516 42196 3547
rect 43070 3544 43076 3556
rect 43128 3544 43134 3596
rect 43346 3593 43352 3596
rect 43341 3584 43352 3593
rect 43307 3556 43352 3584
rect 43341 3547 43352 3556
rect 43346 3544 43352 3547
rect 43404 3544 43410 3596
rect 44634 3584 44640 3596
rect 44595 3556 44640 3584
rect 44634 3544 44640 3556
rect 44692 3544 44698 3596
rect 45281 3587 45339 3593
rect 45281 3553 45293 3587
rect 45327 3584 45339 3587
rect 45738 3584 45744 3596
rect 45327 3556 45744 3584
rect 45327 3553 45339 3556
rect 45281 3547 45339 3553
rect 45738 3544 45744 3556
rect 45796 3544 45802 3596
rect 46290 3584 46296 3596
rect 46251 3556 46296 3584
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 47026 3584 47032 3596
rect 46987 3556 47032 3584
rect 47026 3544 47032 3556
rect 47084 3544 47090 3596
rect 47762 3584 47768 3596
rect 47723 3556 47768 3584
rect 47762 3544 47768 3556
rect 47820 3544 47826 3596
rect 47854 3544 47860 3596
rect 47912 3584 47918 3596
rect 48501 3587 48559 3593
rect 48501 3584 48513 3587
rect 47912 3556 48513 3584
rect 47912 3544 47918 3556
rect 48501 3553 48513 3556
rect 48547 3553 48559 3587
rect 48501 3547 48559 3553
rect 49602 3544 49608 3596
rect 49660 3584 49666 3596
rect 49789 3587 49847 3593
rect 49789 3584 49801 3587
rect 49660 3556 49801 3584
rect 49660 3544 49666 3556
rect 49789 3553 49801 3556
rect 49835 3553 49847 3587
rect 49789 3547 49847 3553
rect 50154 3544 50160 3596
rect 50212 3584 50218 3596
rect 50341 3587 50399 3593
rect 50341 3584 50353 3587
rect 50212 3556 50353 3584
rect 50212 3544 50218 3556
rect 50341 3553 50353 3556
rect 50387 3553 50399 3587
rect 50341 3547 50399 3553
rect 52089 3587 52147 3593
rect 52089 3553 52101 3587
rect 52135 3584 52147 3587
rect 52638 3584 52644 3596
rect 52135 3556 52644 3584
rect 52135 3553 52147 3556
rect 52089 3547 52147 3553
rect 52638 3544 52644 3556
rect 52696 3544 52702 3596
rect 53006 3584 53012 3596
rect 52967 3556 53012 3584
rect 53006 3544 53012 3556
rect 53064 3544 53070 3596
rect 53929 3587 53987 3593
rect 53929 3584 53941 3587
rect 53116 3556 53941 3584
rect 42168 3488 43576 3516
rect 43548 3457 43576 3488
rect 43533 3451 43591 3457
rect 41386 3420 43484 3448
rect 2464 3408 2470 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 3237 3383 3295 3389
rect 3237 3380 3249 3383
rect 2924 3352 3249 3380
rect 2924 3340 2930 3352
rect 3237 3349 3249 3352
rect 3283 3349 3295 3383
rect 3237 3343 3295 3349
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4614 3380 4620 3392
rect 4479 3352 4620 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5074 3380 5080 3392
rect 5035 3352 5080 3380
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 30561 3383 30619 3389
rect 30561 3349 30573 3383
rect 30607 3380 30619 3383
rect 31110 3380 31116 3392
rect 30607 3352 31116 3380
rect 30607 3349 30619 3352
rect 30561 3343 30619 3349
rect 31110 3340 31116 3352
rect 31168 3340 31174 3392
rect 31386 3380 31392 3392
rect 31347 3352 31392 3380
rect 31386 3340 31392 3352
rect 31444 3340 31450 3392
rect 32030 3380 32036 3392
rect 31991 3352 32036 3380
rect 32030 3340 32036 3352
rect 32088 3340 32094 3392
rect 32769 3383 32827 3389
rect 32769 3349 32781 3383
rect 32815 3380 32827 3383
rect 33134 3380 33140 3392
rect 32815 3352 33140 3380
rect 32815 3349 32827 3352
rect 32769 3343 32827 3349
rect 33134 3340 33140 3352
rect 33192 3340 33198 3392
rect 33226 3340 33232 3392
rect 33284 3380 33290 3392
rect 33413 3383 33471 3389
rect 33413 3380 33425 3383
rect 33284 3352 33425 3380
rect 33284 3340 33290 3352
rect 33413 3349 33425 3352
rect 33459 3349 33471 3383
rect 33413 3343 33471 3349
rect 34146 3340 34152 3392
rect 34204 3380 34210 3392
rect 34333 3383 34391 3389
rect 34333 3380 34345 3383
rect 34204 3352 34345 3380
rect 34204 3340 34210 3352
rect 34333 3349 34345 3352
rect 34379 3349 34391 3383
rect 34333 3343 34391 3349
rect 35250 3340 35256 3392
rect 35308 3380 35314 3392
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35308 3352 35909 3380
rect 35308 3340 35314 3352
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 36998 3340 37004 3392
rect 37056 3380 37062 3392
rect 37185 3383 37243 3389
rect 37185 3380 37197 3383
rect 37056 3352 37197 3380
rect 37056 3340 37062 3352
rect 37185 3349 37197 3352
rect 37231 3349 37243 3383
rect 37185 3343 37243 3349
rect 37918 3340 37924 3392
rect 37976 3380 37982 3392
rect 38105 3383 38163 3389
rect 38105 3380 38117 3383
rect 37976 3352 38117 3380
rect 37976 3340 37982 3352
rect 38105 3349 38117 3352
rect 38151 3349 38163 3383
rect 38105 3343 38163 3349
rect 38838 3340 38844 3392
rect 38896 3380 38902 3392
rect 39025 3383 39083 3389
rect 39025 3380 39037 3383
rect 38896 3352 39037 3380
rect 38896 3340 38902 3352
rect 39025 3349 39037 3352
rect 39071 3349 39083 3383
rect 39025 3343 39083 3349
rect 39577 3383 39635 3389
rect 39577 3349 39589 3383
rect 39623 3380 39635 3383
rect 40218 3380 40224 3392
rect 39623 3352 40224 3380
rect 39623 3349 39635 3352
rect 39577 3343 39635 3349
rect 40218 3340 40224 3352
rect 40276 3340 40282 3392
rect 40957 3383 41015 3389
rect 40957 3349 40969 3383
rect 41003 3380 41015 3383
rect 41782 3380 41788 3392
rect 41003 3352 41788 3380
rect 41003 3349 41015 3352
rect 40957 3343 41015 3349
rect 41782 3340 41788 3352
rect 41840 3340 41846 3392
rect 41966 3380 41972 3392
rect 41927 3352 41972 3380
rect 41966 3340 41972 3352
rect 42024 3340 42030 3392
rect 42610 3340 42616 3392
rect 42668 3380 42674 3392
rect 42797 3383 42855 3389
rect 42797 3380 42809 3383
rect 42668 3352 42809 3380
rect 42668 3340 42674 3352
rect 42797 3349 42809 3352
rect 42843 3349 42855 3383
rect 43456 3380 43484 3420
rect 43533 3417 43545 3451
rect 43579 3448 43591 3451
rect 44652 3448 44680 3544
rect 47578 3516 47584 3528
rect 43579 3420 44680 3448
rect 45020 3488 47584 3516
rect 43579 3417 43591 3420
rect 43533 3411 43591 3417
rect 45020 3380 45048 3488
rect 47578 3476 47584 3488
rect 47636 3476 47642 3528
rect 47946 3476 47952 3528
rect 48004 3516 48010 3528
rect 53116 3516 53144 3556
rect 53929 3553 53941 3556
rect 53975 3553 53987 3587
rect 53929 3547 53987 3553
rect 55033 3587 55091 3593
rect 55033 3553 55045 3587
rect 55079 3584 55091 3587
rect 55214 3584 55220 3596
rect 55079 3556 55220 3584
rect 55079 3553 55091 3556
rect 55033 3547 55091 3553
rect 55214 3544 55220 3556
rect 55272 3544 55278 3596
rect 55315 3584 55343 3624
rect 55585 3621 55597 3655
rect 55631 3652 55643 3655
rect 55766 3652 55772 3664
rect 55631 3624 55772 3652
rect 55631 3621 55643 3624
rect 55585 3615 55643 3621
rect 55766 3612 55772 3624
rect 55824 3612 55830 3664
rect 56870 3652 56876 3664
rect 56831 3624 56876 3652
rect 56870 3612 56876 3624
rect 56928 3612 56934 3664
rect 55315 3556 56088 3584
rect 48004 3488 53144 3516
rect 48004 3476 48010 3488
rect 53650 3476 53656 3528
rect 53708 3516 53714 3528
rect 53745 3519 53803 3525
rect 53745 3516 53757 3519
rect 53708 3488 53757 3516
rect 53708 3476 53714 3488
rect 53745 3485 53757 3488
rect 53791 3485 53803 3519
rect 56060 3516 56088 3556
rect 56410 3544 56416 3596
rect 56468 3584 56474 3596
rect 57606 3584 57612 3596
rect 56468 3556 57612 3584
rect 56468 3544 56474 3556
rect 57606 3544 57612 3556
rect 57664 3544 57670 3596
rect 57716 3593 57744 3692
rect 57701 3587 57759 3593
rect 57701 3553 57713 3587
rect 57747 3553 57759 3587
rect 57701 3547 57759 3553
rect 57333 3519 57391 3525
rect 57333 3516 57345 3519
rect 56060 3488 57345 3516
rect 53745 3479 53803 3485
rect 57333 3485 57345 3488
rect 57379 3516 57391 3519
rect 57517 3519 57575 3525
rect 57517 3516 57529 3519
rect 57379 3488 57529 3516
rect 57379 3485 57391 3488
rect 57333 3479 57391 3485
rect 57517 3485 57529 3488
rect 57563 3485 57575 3519
rect 57517 3479 57575 3485
rect 45097 3451 45155 3457
rect 45097 3417 45109 3451
rect 45143 3448 45155 3451
rect 48958 3448 48964 3460
rect 45143 3420 48964 3448
rect 45143 3417 45155 3420
rect 45097 3411 45155 3417
rect 48958 3408 48964 3420
rect 49016 3408 49022 3460
rect 49050 3408 49056 3460
rect 49108 3448 49114 3460
rect 55214 3448 55220 3460
rect 49108 3420 55220 3448
rect 49108 3408 49114 3420
rect 55214 3408 55220 3420
rect 55272 3408 55278 3460
rect 55766 3448 55772 3460
rect 55727 3420 55772 3448
rect 55766 3408 55772 3420
rect 55824 3408 55830 3460
rect 43456 3352 45048 3380
rect 42797 3343 42855 3349
rect 45370 3340 45376 3392
rect 45428 3380 45434 3392
rect 46385 3383 46443 3389
rect 46385 3380 46397 3383
rect 45428 3352 46397 3380
rect 45428 3340 45434 3352
rect 46385 3349 46397 3352
rect 46431 3349 46443 3383
rect 46385 3343 46443 3349
rect 46474 3340 46480 3392
rect 46532 3380 46538 3392
rect 47121 3383 47179 3389
rect 47121 3380 47133 3383
rect 46532 3352 47133 3380
rect 46532 3340 46538 3352
rect 47121 3349 47133 3352
rect 47167 3349 47179 3383
rect 47121 3343 47179 3349
rect 47302 3340 47308 3392
rect 47360 3380 47366 3392
rect 47857 3383 47915 3389
rect 47857 3380 47869 3383
rect 47360 3352 47869 3380
rect 47360 3340 47366 3352
rect 47857 3349 47869 3352
rect 47903 3349 47915 3383
rect 47857 3343 47915 3349
rect 48222 3340 48228 3392
rect 48280 3380 48286 3392
rect 48593 3383 48651 3389
rect 48593 3380 48605 3383
rect 48280 3352 48605 3380
rect 48280 3340 48286 3352
rect 48593 3349 48605 3352
rect 48639 3349 48651 3383
rect 49602 3380 49608 3392
rect 49563 3352 49608 3380
rect 48593 3343 48651 3349
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 51994 3340 52000 3392
rect 52052 3380 52058 3392
rect 52181 3383 52239 3389
rect 52181 3380 52193 3383
rect 52052 3352 52193 3380
rect 52052 3340 52058 3352
rect 52181 3349 52193 3352
rect 52227 3349 52239 3383
rect 52181 3343 52239 3349
rect 52914 3340 52920 3392
rect 52972 3380 52978 3392
rect 53101 3383 53159 3389
rect 53101 3380 53113 3383
rect 52972 3352 53113 3380
rect 52972 3340 52978 3352
rect 53101 3349 53113 3352
rect 53147 3349 53159 3383
rect 54386 3380 54392 3392
rect 54347 3352 54392 3380
rect 53101 3343 53159 3349
rect 54386 3340 54392 3352
rect 54444 3340 54450 3392
rect 54849 3383 54907 3389
rect 54849 3349 54861 3383
rect 54895 3380 54907 3383
rect 55306 3380 55312 3392
rect 54895 3352 55312 3380
rect 54895 3349 54907 3352
rect 54849 3343 54907 3349
rect 55306 3340 55312 3352
rect 55364 3340 55370 3392
rect 56410 3340 56416 3392
rect 56468 3380 56474 3392
rect 56965 3383 57023 3389
rect 56965 3380 56977 3383
rect 56468 3352 56977 3380
rect 56468 3340 56474 3352
rect 56965 3349 56977 3352
rect 57011 3349 57023 3383
rect 57974 3380 57980 3392
rect 57935 3352 57980 3380
rect 56965 3343 57023 3349
rect 57974 3340 57980 3352
rect 58032 3340 58038 3392
rect 1104 3290 58880 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 58880 3290
rect 1104 3216 58880 3238
rect 3142 3176 3148 3188
rect 3103 3148 3148 3176
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 3970 3136 3976 3188
rect 4028 3176 4034 3188
rect 4617 3179 4675 3185
rect 4617 3176 4629 3179
rect 4028 3148 4629 3176
rect 4028 3136 4034 3148
rect 4617 3145 4629 3148
rect 4663 3145 4675 3179
rect 34238 3176 34244 3188
rect 34199 3148 34244 3176
rect 4617 3139 4675 3145
rect 34238 3136 34244 3148
rect 34296 3136 34302 3188
rect 37366 3176 37372 3188
rect 37327 3148 37372 3176
rect 37366 3136 37372 3148
rect 37424 3136 37430 3188
rect 38654 3176 38660 3188
rect 38615 3148 38660 3176
rect 38654 3136 38660 3148
rect 38712 3136 38718 3188
rect 43530 3136 43536 3188
rect 43588 3176 43594 3188
rect 46201 3179 46259 3185
rect 43588 3148 46152 3176
rect 43588 3136 43594 3148
rect 4062 3108 4068 3120
rect 2792 3080 4068 3108
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2792 3049 2820 3080
rect 4062 3068 4068 3080
rect 4120 3068 4126 3120
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 6273 3111 6331 3117
rect 6273 3108 6285 3111
rect 4764 3080 6285 3108
rect 4764 3068 4770 3080
rect 6273 3077 6285 3080
rect 6319 3077 6331 3111
rect 6273 3071 6331 3077
rect 29273 3111 29331 3117
rect 29273 3077 29285 3111
rect 29319 3108 29331 3111
rect 29319 3080 30144 3108
rect 29319 3077 29331 3080
rect 29273 3071 29331 3077
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2958 3040 2964 3052
rect 2919 3012 2964 3040
rect 2777 3003 2835 3009
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 30116 3049 30144 3080
rect 30484 3080 40724 3108
rect 28813 3043 28871 3049
rect 5460 3012 26234 3040
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 3752 2944 4813 2972
rect 3752 2932 3758 2944
rect 4801 2941 4813 2944
rect 4847 2972 4859 2975
rect 5350 2972 5356 2984
rect 4847 2944 5356 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 5350 2932 5356 2944
rect 5408 2932 5414 2984
rect 5460 2981 5488 3012
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 6273 2975 6331 2981
rect 6273 2941 6285 2975
rect 6319 2972 6331 2975
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6319 2944 6837 2972
rect 6319 2941 6331 2944
rect 6273 2935 6331 2941
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7064 2944 7481 2972
rect 7064 2932 7070 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 8846 2972 8852 2984
rect 8807 2944 8852 2972
rect 7469 2935 7527 2941
rect 8846 2932 8852 2944
rect 8904 2932 8910 2984
rect 26206 2972 26234 3012
rect 28813 3009 28825 3043
rect 28859 3040 28871 3043
rect 29917 3043 29975 3049
rect 29917 3040 29929 3043
rect 28859 3012 29929 3040
rect 28859 3009 28871 3012
rect 28813 3003 28871 3009
rect 29917 3009 29929 3012
rect 29963 3009 29975 3043
rect 29917 3003 29975 3009
rect 30101 3043 30159 3049
rect 30101 3009 30113 3043
rect 30147 3009 30159 3043
rect 30101 3003 30159 3009
rect 29457 2975 29515 2981
rect 29457 2972 29469 2975
rect 26206 2944 29469 2972
rect 29457 2941 29469 2944
rect 29503 2972 29515 2975
rect 30484 2972 30512 3080
rect 33689 3043 33747 3049
rect 33689 3009 33701 3043
rect 33735 3040 33747 3043
rect 33962 3040 33968 3052
rect 33735 3012 33968 3040
rect 33735 3009 33747 3012
rect 33689 3003 33747 3009
rect 33962 3000 33968 3012
rect 34020 3000 34026 3052
rect 35526 3040 35532 3052
rect 35487 3012 35532 3040
rect 35526 3000 35532 3012
rect 35584 3000 35590 3052
rect 38470 3040 38476 3052
rect 38431 3012 38476 3040
rect 38470 3000 38476 3012
rect 38528 3000 38534 3052
rect 40037 3043 40095 3049
rect 40037 3009 40049 3043
rect 40083 3040 40095 3043
rect 40494 3040 40500 3052
rect 40083 3012 40500 3040
rect 40083 3009 40095 3012
rect 40037 3003 40095 3009
rect 40494 3000 40500 3012
rect 40552 3000 40558 3052
rect 40696 3040 40724 3080
rect 41386 3080 44128 3108
rect 41386 3040 41414 3080
rect 40696 3012 41414 3040
rect 41966 3000 41972 3052
rect 42024 3040 42030 3052
rect 43717 3043 43775 3049
rect 43717 3040 43729 3043
rect 42024 3012 43729 3040
rect 42024 3000 42030 3012
rect 43717 3009 43729 3012
rect 43763 3009 43775 3043
rect 43717 3003 43775 3009
rect 31294 2972 31300 2984
rect 29503 2944 30512 2972
rect 31255 2944 31300 2972
rect 29503 2941 29515 2944
rect 29457 2935 29515 2941
rect 31294 2932 31300 2944
rect 31352 2932 31358 2984
rect 33229 2975 33287 2981
rect 33229 2941 33241 2975
rect 33275 2972 33287 2975
rect 33410 2972 33416 2984
rect 33275 2944 33416 2972
rect 33275 2941 33287 2944
rect 33229 2935 33287 2941
rect 33410 2932 33416 2944
rect 33468 2932 33474 2984
rect 33873 2975 33931 2981
rect 33873 2941 33885 2975
rect 33919 2941 33931 2975
rect 33873 2935 33931 2941
rect 35345 2975 35403 2981
rect 35345 2941 35357 2975
rect 35391 2972 35403 2975
rect 35894 2972 35900 2984
rect 35391 2944 35900 2972
rect 35391 2941 35403 2944
rect 35345 2935 35403 2941
rect 3970 2904 3976 2916
rect 3931 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4154 2904 4160 2916
rect 4115 2876 4160 2904
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 5626 2904 5632 2916
rect 4264 2876 5632 2904
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 4264 2836 4292 2876
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 31938 2904 31944 2916
rect 31899 2876 31944 2904
rect 31938 2864 31944 2876
rect 31996 2864 32002 2916
rect 32125 2907 32183 2913
rect 32125 2873 32137 2907
rect 32171 2904 32183 2907
rect 32306 2904 32312 2916
rect 32171 2876 32312 2904
rect 32171 2873 32183 2876
rect 32125 2867 32183 2873
rect 32306 2864 32312 2876
rect 32364 2864 32370 2916
rect 3292 2808 4292 2836
rect 3292 2796 3298 2808
rect 4338 2796 4344 2848
rect 4396 2836 4402 2848
rect 5074 2836 5080 2848
rect 4396 2808 5080 2836
rect 4396 2796 4402 2808
rect 5074 2796 5080 2808
rect 5132 2796 5138 2848
rect 5258 2836 5264 2848
rect 5219 2808 5264 2836
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 30558 2836 30564 2848
rect 30519 2808 30564 2836
rect 30558 2796 30564 2808
rect 30616 2796 30622 2848
rect 31113 2839 31171 2845
rect 31113 2805 31125 2839
rect 31159 2836 31171 2839
rect 32214 2836 32220 2848
rect 31159 2808 32220 2836
rect 31159 2805 31171 2808
rect 31113 2799 31171 2805
rect 32214 2796 32220 2808
rect 32272 2796 32278 2848
rect 33045 2839 33103 2845
rect 33045 2805 33057 2839
rect 33091 2836 33103 2839
rect 33888 2836 33916 2935
rect 35894 2932 35900 2944
rect 35952 2932 35958 2984
rect 37182 2972 37188 2984
rect 37143 2944 37188 2972
rect 37182 2932 37188 2944
rect 37240 2932 37246 2984
rect 38289 2975 38347 2981
rect 38289 2941 38301 2975
rect 38335 2972 38347 2975
rect 39114 2972 39120 2984
rect 38335 2944 39120 2972
rect 38335 2941 38347 2944
rect 38289 2935 38347 2941
rect 39114 2932 39120 2944
rect 39172 2932 39178 2984
rect 39577 2975 39635 2981
rect 39577 2941 39589 2975
rect 39623 2972 39635 2975
rect 39758 2972 39764 2984
rect 39623 2944 39764 2972
rect 39623 2941 39635 2944
rect 39577 2935 39635 2941
rect 35989 2907 36047 2913
rect 35989 2873 36001 2907
rect 36035 2904 36047 2907
rect 36541 2907 36599 2913
rect 36541 2904 36553 2907
rect 36035 2876 36553 2904
rect 36035 2873 36047 2876
rect 35989 2867 36047 2873
rect 36541 2873 36553 2876
rect 36587 2873 36599 2907
rect 36541 2867 36599 2873
rect 37366 2864 37372 2916
rect 37424 2904 37430 2916
rect 39592 2904 39620 2935
rect 39758 2932 39764 2944
rect 39816 2932 39822 2984
rect 40221 2975 40279 2981
rect 40221 2941 40233 2975
rect 40267 2941 40279 2975
rect 40221 2935 40279 2941
rect 37424 2876 39620 2904
rect 37424 2864 37430 2876
rect 33091 2808 33916 2836
rect 33091 2805 33103 2808
rect 33045 2799 33103 2805
rect 36078 2796 36084 2848
rect 36136 2836 36142 2848
rect 36633 2839 36691 2845
rect 36633 2836 36645 2839
rect 36136 2808 36645 2836
rect 36136 2796 36142 2808
rect 36633 2805 36645 2808
rect 36679 2805 36691 2839
rect 36633 2799 36691 2805
rect 39393 2839 39451 2845
rect 39393 2805 39405 2839
rect 39439 2836 39451 2839
rect 40236 2836 40264 2935
rect 42794 2932 42800 2984
rect 42852 2972 42858 2984
rect 43533 2975 43591 2981
rect 43533 2972 43545 2975
rect 42852 2944 43545 2972
rect 42852 2932 42858 2944
rect 43533 2941 43545 2944
rect 43579 2941 43591 2975
rect 44100 2972 44128 3080
rect 45462 3068 45468 3120
rect 45520 3108 45526 3120
rect 46124 3108 46152 3148
rect 46201 3145 46213 3179
rect 46247 3176 46259 3179
rect 47026 3176 47032 3188
rect 46247 3148 47032 3176
rect 46247 3145 46259 3148
rect 46201 3139 46259 3145
rect 47026 3136 47032 3148
rect 47084 3136 47090 3188
rect 47854 3176 47860 3188
rect 47815 3148 47860 3176
rect 47854 3136 47860 3148
rect 47912 3136 47918 3188
rect 49234 3136 49240 3188
rect 49292 3176 49298 3188
rect 51534 3176 51540 3188
rect 49292 3148 51540 3176
rect 49292 3136 49298 3148
rect 51534 3136 51540 3148
rect 51592 3136 51598 3188
rect 53006 3176 53012 3188
rect 52967 3148 53012 3176
rect 53006 3136 53012 3148
rect 53064 3136 53070 3188
rect 53098 3136 53104 3188
rect 53156 3176 53162 3188
rect 54846 3176 54852 3188
rect 53156 3148 54852 3176
rect 53156 3136 53162 3148
rect 54846 3136 54852 3148
rect 54904 3136 54910 3188
rect 55030 3136 55036 3188
rect 55088 3176 55094 3188
rect 55953 3179 56011 3185
rect 55953 3176 55965 3179
rect 55088 3148 55965 3176
rect 55088 3136 55094 3148
rect 55953 3145 55965 3148
rect 55999 3145 56011 3179
rect 55953 3139 56011 3145
rect 56226 3136 56232 3188
rect 56284 3176 56290 3188
rect 57977 3179 58035 3185
rect 56284 3148 57928 3176
rect 56284 3136 56290 3148
rect 57238 3108 57244 3120
rect 45520 3080 45784 3108
rect 46124 3080 56916 3108
rect 57199 3080 57244 3108
rect 45520 3068 45526 3080
rect 44177 3043 44235 3049
rect 44177 3009 44189 3043
rect 44223 3040 44235 3043
rect 45557 3043 45615 3049
rect 44223 3012 45508 3040
rect 44223 3009 44235 3012
rect 44177 3003 44235 3009
rect 45480 2972 45508 3012
rect 45557 3009 45569 3043
rect 45603 3040 45615 3043
rect 45646 3040 45652 3052
rect 45603 3012 45652 3040
rect 45603 3009 45615 3012
rect 45557 3003 45615 3009
rect 45646 3000 45652 3012
rect 45704 3000 45710 3052
rect 45756 3049 45784 3080
rect 45741 3043 45799 3049
rect 45741 3009 45753 3043
rect 45787 3009 45799 3043
rect 45741 3003 45799 3009
rect 47118 3000 47124 3052
rect 47176 3040 47182 3052
rect 47213 3043 47271 3049
rect 47213 3040 47225 3043
rect 47176 3012 47225 3040
rect 47176 3000 47182 3012
rect 47213 3009 47225 3012
rect 47259 3009 47271 3043
rect 47394 3040 47400 3052
rect 47355 3012 47400 3040
rect 47213 3003 47271 3009
rect 47394 3000 47400 3012
rect 47452 3000 47458 3052
rect 48590 3000 48596 3052
rect 48648 3040 48654 3052
rect 48777 3043 48835 3049
rect 48777 3040 48789 3043
rect 48648 3012 48789 3040
rect 48648 3000 48654 3012
rect 48777 3009 48789 3012
rect 48823 3009 48835 3043
rect 48958 3040 48964 3052
rect 48919 3012 48964 3040
rect 48777 3003 48835 3009
rect 48958 3000 48964 3012
rect 49016 3000 49022 3052
rect 52549 3043 52607 3049
rect 52549 3040 52561 3043
rect 51828 3012 52561 3040
rect 46750 2972 46756 2984
rect 44100 2944 45140 2972
rect 45480 2944 46756 2972
rect 43533 2935 43591 2941
rect 40681 2907 40739 2913
rect 40681 2873 40693 2907
rect 40727 2904 40739 2907
rect 41233 2907 41291 2913
rect 41233 2904 41245 2907
rect 40727 2876 41245 2904
rect 40727 2873 40739 2876
rect 40681 2867 40739 2873
rect 41233 2873 41245 2876
rect 41279 2873 41291 2907
rect 41966 2904 41972 2916
rect 41927 2876 41972 2904
rect 41233 2867 41291 2873
rect 41966 2864 41972 2876
rect 42024 2864 42030 2916
rect 44726 2904 44732 2916
rect 44687 2876 44732 2904
rect 44726 2864 44732 2876
rect 44784 2864 44790 2916
rect 39439 2808 40264 2836
rect 39439 2805 39451 2808
rect 39393 2799 39451 2805
rect 40770 2796 40776 2848
rect 40828 2836 40834 2848
rect 41325 2839 41383 2845
rect 41325 2836 41337 2839
rect 40828 2808 41337 2836
rect 40828 2796 40834 2808
rect 41325 2805 41337 2808
rect 41371 2805 41383 2839
rect 41325 2799 41383 2805
rect 41690 2796 41696 2848
rect 41748 2836 41754 2848
rect 42061 2839 42119 2845
rect 42061 2836 42073 2839
rect 41748 2808 42073 2836
rect 41748 2796 41754 2808
rect 42061 2805 42073 2808
rect 42107 2805 42119 2839
rect 42061 2799 42119 2805
rect 44450 2796 44456 2848
rect 44508 2836 44514 2848
rect 44821 2839 44879 2845
rect 44821 2836 44833 2839
rect 44508 2808 44833 2836
rect 44508 2796 44514 2808
rect 44821 2805 44833 2808
rect 44867 2805 44879 2839
rect 45112 2836 45140 2944
rect 46750 2932 46756 2944
rect 46808 2932 46814 2984
rect 49326 2932 49332 2984
rect 49384 2972 49390 2984
rect 51828 2972 51856 3012
rect 52549 3009 52561 3012
rect 52595 3009 52607 3043
rect 52549 3003 52607 3009
rect 55490 3000 55496 3052
rect 55548 3040 55554 3052
rect 56888 3049 56916 3080
rect 57238 3068 57244 3080
rect 57296 3068 57302 3120
rect 57900 3108 57928 3148
rect 57977 3145 57989 3179
rect 58023 3176 58035 3179
rect 58066 3176 58072 3188
rect 58023 3148 58072 3176
rect 58023 3145 58035 3148
rect 57977 3139 58035 3145
rect 58066 3136 58072 3148
rect 58124 3136 58130 3188
rect 58526 3108 58532 3120
rect 57900 3080 58532 3108
rect 58526 3068 58532 3080
rect 58584 3068 58590 3120
rect 55585 3043 55643 3049
rect 55585 3040 55597 3043
rect 55548 3012 55597 3040
rect 55548 3000 55554 3012
rect 55585 3009 55597 3012
rect 55631 3009 55643 3043
rect 55585 3003 55643 3009
rect 56873 3043 56931 3049
rect 56873 3009 56885 3043
rect 56919 3009 56931 3043
rect 57054 3040 57060 3052
rect 57015 3012 57060 3040
rect 56873 3003 56931 3009
rect 57054 3000 57060 3012
rect 57112 3000 57118 3052
rect 52362 2972 52368 2984
rect 49384 2944 51856 2972
rect 52323 2944 52368 2972
rect 49384 2932 49390 2944
rect 52362 2932 52368 2944
rect 52420 2932 52426 2984
rect 53392 2944 54340 2972
rect 45278 2864 45284 2916
rect 45336 2904 45342 2916
rect 49050 2904 49056 2916
rect 45336 2876 49056 2904
rect 45336 2864 45342 2876
rect 49050 2864 49056 2876
rect 49108 2864 49114 2916
rect 49421 2907 49479 2913
rect 49421 2873 49433 2907
rect 49467 2904 49479 2907
rect 49973 2907 50031 2913
rect 49973 2904 49985 2907
rect 49467 2876 49985 2904
rect 49467 2873 49479 2876
rect 49421 2867 49479 2873
rect 49973 2873 49985 2876
rect 50019 2873 50031 2907
rect 50706 2904 50712 2916
rect 50667 2876 50712 2904
rect 49973 2867 50031 2873
rect 50706 2864 50712 2876
rect 50764 2864 50770 2916
rect 51442 2904 51448 2916
rect 51403 2876 51448 2904
rect 51442 2864 51448 2876
rect 51500 2864 51506 2916
rect 51626 2864 51632 2916
rect 51684 2904 51690 2916
rect 53392 2904 53420 2944
rect 54110 2904 54116 2916
rect 51684 2876 53420 2904
rect 54071 2876 54116 2904
rect 51684 2864 51690 2876
rect 54110 2864 54116 2876
rect 54168 2864 54174 2916
rect 54312 2904 54340 2944
rect 54386 2932 54392 2984
rect 54444 2972 54450 2984
rect 54849 2975 54907 2981
rect 54849 2972 54861 2975
rect 54444 2944 54861 2972
rect 54444 2932 54450 2944
rect 54849 2941 54861 2944
rect 54895 2941 54907 2975
rect 54849 2935 54907 2941
rect 55769 2975 55827 2981
rect 55769 2941 55781 2975
rect 55815 2941 55827 2975
rect 55769 2935 55827 2941
rect 55784 2904 55812 2935
rect 55950 2932 55956 2984
rect 56008 2972 56014 2984
rect 58161 2975 58219 2981
rect 58161 2972 58173 2975
rect 56008 2944 58173 2972
rect 56008 2932 56014 2944
rect 58161 2941 58173 2944
rect 58207 2941 58219 2975
rect 58161 2935 58219 2941
rect 54312 2876 55812 2904
rect 55858 2864 55864 2916
rect 55916 2904 55922 2916
rect 59446 2904 59452 2916
rect 55916 2876 59452 2904
rect 55916 2864 55922 2876
rect 59446 2864 59452 2876
rect 59504 2864 59510 2916
rect 48406 2836 48412 2848
rect 45112 2808 48412 2836
rect 44821 2799 44879 2805
rect 48406 2796 48412 2808
rect 48464 2796 48470 2848
rect 49142 2796 49148 2848
rect 49200 2836 49206 2848
rect 50065 2839 50123 2845
rect 50065 2836 50077 2839
rect 49200 2808 50077 2836
rect 49200 2796 49206 2808
rect 50065 2805 50077 2808
rect 50111 2805 50123 2839
rect 50065 2799 50123 2805
rect 50154 2796 50160 2848
rect 50212 2836 50218 2848
rect 50801 2839 50859 2845
rect 50801 2836 50813 2839
rect 50212 2808 50813 2836
rect 50212 2796 50218 2808
rect 50801 2805 50813 2808
rect 50847 2805 50859 2839
rect 50801 2799 50859 2805
rect 51074 2796 51080 2848
rect 51132 2836 51138 2848
rect 51537 2839 51595 2845
rect 51537 2836 51549 2839
rect 51132 2808 51549 2836
rect 51132 2796 51138 2808
rect 51537 2805 51549 2808
rect 51583 2805 51595 2839
rect 51537 2799 51595 2805
rect 53834 2796 53840 2848
rect 53892 2836 53898 2848
rect 54205 2839 54263 2845
rect 54205 2836 54217 2839
rect 53892 2808 54217 2836
rect 53892 2796 53898 2808
rect 54205 2805 54217 2808
rect 54251 2805 54263 2839
rect 54205 2799 54263 2805
rect 54754 2796 54760 2848
rect 54812 2836 54818 2848
rect 54941 2839 54999 2845
rect 54941 2836 54953 2839
rect 54812 2808 54953 2836
rect 54812 2796 54818 2808
rect 54941 2805 54953 2808
rect 54987 2805 54999 2839
rect 54941 2799 54999 2805
rect 1104 2746 58880 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 50326 2746
rect 50378 2694 50390 2746
rect 50442 2694 50454 2746
rect 50506 2694 50518 2746
rect 50570 2694 58880 2746
rect 1104 2672 58880 2694
rect 2317 2635 2375 2641
rect 2317 2601 2329 2635
rect 2363 2632 2375 2635
rect 3970 2632 3976 2644
rect 2363 2604 3976 2632
rect 2363 2601 2375 2604
rect 2317 2595 2375 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 35345 2635 35403 2641
rect 35345 2601 35357 2635
rect 35391 2632 35403 2635
rect 35802 2632 35808 2644
rect 35391 2604 35808 2632
rect 35391 2601 35403 2604
rect 35345 2595 35403 2601
rect 35802 2592 35808 2604
rect 35860 2592 35866 2644
rect 36909 2635 36967 2641
rect 36909 2601 36921 2635
rect 36955 2632 36967 2635
rect 37090 2632 37096 2644
rect 36955 2604 37096 2632
rect 36955 2601 36967 2604
rect 36909 2595 36967 2601
rect 37090 2592 37096 2604
rect 37148 2592 37154 2644
rect 38930 2592 38936 2644
rect 38988 2632 38994 2644
rect 39577 2635 39635 2641
rect 39577 2632 39589 2635
rect 38988 2604 39589 2632
rect 38988 2592 38994 2604
rect 39577 2601 39589 2604
rect 39623 2601 39635 2635
rect 39577 2595 39635 2601
rect 44726 2592 44732 2644
rect 44784 2632 44790 2644
rect 44913 2635 44971 2641
rect 44913 2632 44925 2635
rect 44784 2604 44925 2632
rect 44784 2592 44790 2604
rect 44913 2601 44925 2604
rect 44959 2601 44971 2635
rect 44913 2595 44971 2601
rect 46017 2635 46075 2641
rect 46017 2601 46029 2635
rect 46063 2632 46075 2635
rect 46290 2632 46296 2644
rect 46063 2604 46296 2632
rect 46063 2601 46075 2604
rect 46017 2595 46075 2601
rect 46290 2592 46296 2604
rect 46348 2592 46354 2644
rect 47581 2635 47639 2641
rect 47581 2601 47593 2635
rect 47627 2632 47639 2635
rect 47762 2632 47768 2644
rect 47627 2604 47768 2632
rect 47627 2601 47639 2604
rect 47581 2595 47639 2601
rect 47762 2592 47768 2604
rect 47820 2592 47826 2644
rect 50249 2635 50307 2641
rect 50249 2601 50261 2635
rect 50295 2632 50307 2635
rect 50706 2632 50712 2644
rect 50295 2604 50712 2632
rect 50295 2601 50307 2604
rect 50249 2595 50307 2601
rect 50706 2592 50712 2604
rect 50764 2592 50770 2644
rect 51353 2635 51411 2641
rect 51353 2601 51365 2635
rect 51399 2632 51411 2635
rect 51442 2632 51448 2644
rect 51399 2604 51448 2632
rect 51399 2601 51411 2604
rect 51353 2595 51411 2601
rect 51442 2592 51448 2604
rect 51500 2592 51506 2644
rect 54021 2635 54079 2641
rect 54021 2601 54033 2635
rect 54067 2632 54079 2635
rect 54110 2632 54116 2644
rect 54067 2604 54116 2632
rect 54067 2601 54079 2604
rect 54021 2595 54079 2601
rect 54110 2592 54116 2604
rect 54168 2592 54174 2644
rect 55582 2632 55588 2644
rect 55543 2604 55588 2632
rect 55582 2592 55588 2604
rect 55640 2592 55646 2644
rect 56318 2592 56324 2644
rect 56376 2632 56382 2644
rect 56689 2635 56747 2641
rect 56689 2632 56701 2635
rect 56376 2604 56701 2632
rect 56376 2592 56382 2604
rect 56689 2601 56701 2604
rect 56735 2601 56747 2635
rect 56689 2595 56747 2601
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 4893 2567 4951 2573
rect 4893 2564 4905 2567
rect 2915 2536 4905 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 4893 2533 4905 2536
rect 4939 2533 4951 2567
rect 4893 2527 4951 2533
rect 5074 2524 5080 2576
rect 5132 2564 5138 2576
rect 29825 2567 29883 2573
rect 5132 2536 7604 2564
rect 5132 2524 5138 2536
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 4249 2499 4307 2505
rect 1719 2468 3372 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 3344 2428 3372 2468
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 4614 2496 4620 2508
rect 4295 2468 4620 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 7576 2505 7604 2536
rect 29825 2533 29837 2567
rect 29871 2564 29883 2567
rect 30558 2564 30564 2576
rect 29871 2536 30564 2564
rect 29871 2533 29883 2536
rect 29825 2527 29883 2533
rect 30558 2524 30564 2536
rect 30616 2524 30622 2576
rect 37829 2567 37887 2573
rect 37829 2533 37841 2567
rect 37875 2564 37887 2567
rect 40681 2567 40739 2573
rect 40681 2564 40693 2567
rect 37875 2536 40693 2564
rect 37875 2533 37887 2536
rect 37829 2527 37887 2533
rect 40681 2533 40693 2536
rect 40727 2533 40739 2567
rect 40681 2527 40739 2533
rect 46750 2524 46756 2576
rect 46808 2564 46814 2576
rect 48133 2567 48191 2573
rect 48133 2564 48145 2567
rect 46808 2536 48145 2564
rect 46808 2524 46814 2536
rect 48133 2533 48145 2536
rect 48179 2533 48191 2567
rect 48133 2527 48191 2533
rect 48866 2524 48872 2576
rect 48924 2564 48930 2576
rect 55214 2564 55220 2576
rect 48924 2536 50936 2564
rect 48924 2524 48930 2536
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 5684 2468 6929 2496
rect 5684 2456 5690 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8205 2499 8263 2505
rect 8205 2496 8217 2499
rect 7984 2468 8217 2496
rect 7984 2456 7990 2468
rect 8205 2465 8217 2468
rect 8251 2465 8263 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8205 2459 8263 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 10778 2496 10784 2508
rect 10739 2468 10784 2496
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11756 2468 12265 2496
rect 11756 2456 11762 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12676 2468 12909 2496
rect 12676 2456 12682 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 13538 2496 13544 2508
rect 13499 2468 13544 2496
rect 12897 2459 12955 2465
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 14458 2456 14464 2508
rect 14516 2496 14522 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14516 2468 14933 2496
rect 14516 2456 14522 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15470 2456 15476 2508
rect 15528 2496 15534 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15528 2468 15577 2496
rect 15528 2456 15534 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 16390 2496 16396 2508
rect 16351 2468 16396 2496
rect 15565 2459 15623 2465
rect 16390 2456 16396 2468
rect 16448 2456 16454 2508
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17368 2468 17601 2496
rect 17368 2456 17374 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 18230 2496 18236 2508
rect 18191 2468 18236 2496
rect 17589 2459 17647 2465
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 19150 2496 19156 2508
rect 19111 2468 19156 2496
rect 19150 2456 19156 2468
rect 19208 2456 19214 2508
rect 20070 2456 20076 2508
rect 20128 2496 20134 2508
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 20128 2468 20269 2496
rect 20128 2456 20134 2468
rect 20257 2465 20269 2468
rect 20303 2465 20315 2499
rect 21082 2496 21088 2508
rect 21043 2468 21088 2496
rect 20257 2459 20315 2465
rect 21082 2456 21088 2468
rect 21140 2456 21146 2508
rect 21821 2499 21879 2505
rect 21821 2465 21833 2499
rect 21867 2496 21879 2499
rect 22002 2496 22008 2508
rect 21867 2468 22008 2496
rect 21867 2465 21879 2468
rect 21821 2459 21879 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 22922 2496 22928 2508
rect 22883 2468 22928 2496
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 23842 2496 23848 2508
rect 23803 2468 23848 2496
rect 23842 2456 23848 2468
rect 23900 2456 23906 2508
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 24820 2468 25605 2496
rect 24820 2456 24826 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 25774 2456 25780 2508
rect 25832 2496 25838 2508
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25832 2468 26249 2496
rect 25832 2456 25838 2468
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 26694 2456 26700 2508
rect 26752 2496 26758 2508
rect 26881 2499 26939 2505
rect 26881 2496 26893 2499
rect 26752 2468 26893 2496
rect 26752 2456 26758 2468
rect 26881 2465 26893 2468
rect 26927 2465 26939 2499
rect 26881 2459 26939 2465
rect 27614 2456 27620 2508
rect 27672 2496 27678 2508
rect 28261 2499 28319 2505
rect 28261 2496 28273 2499
rect 27672 2468 28273 2496
rect 27672 2456 27678 2468
rect 28261 2465 28273 2468
rect 28307 2465 28319 2499
rect 28261 2459 28319 2465
rect 29089 2499 29147 2505
rect 29089 2465 29101 2499
rect 29135 2496 29147 2499
rect 30929 2499 30987 2505
rect 29135 2468 30604 2496
rect 29135 2465 29147 2468
rect 29089 2459 29147 2465
rect 4338 2428 4344 2440
rect 3344 2400 4344 2428
rect 1857 2391 1915 2397
rect 1872 2360 1900 2391
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 5258 2428 5264 2440
rect 4479 2400 5264 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5353 2363 5411 2369
rect 5353 2360 5365 2363
rect 1872 2332 5365 2360
rect 5353 2329 5365 2332
rect 5399 2329 5411 2363
rect 5353 2323 5411 2329
rect 30009 2363 30067 2369
rect 30009 2329 30021 2363
rect 30055 2360 30067 2363
rect 30466 2360 30472 2372
rect 30055 2332 30472 2360
rect 30055 2329 30067 2332
rect 30009 2323 30067 2329
rect 30466 2320 30472 2332
rect 30524 2320 30530 2372
rect 30576 2360 30604 2468
rect 30929 2465 30941 2499
rect 30975 2496 30987 2499
rect 31386 2496 31392 2508
rect 30975 2468 31392 2496
rect 30975 2465 30987 2468
rect 30929 2459 30987 2465
rect 31386 2456 31392 2468
rect 31444 2456 31450 2508
rect 32030 2496 32036 2508
rect 31991 2468 32036 2496
rect 32030 2456 32036 2468
rect 32088 2456 32094 2508
rect 32214 2496 32220 2508
rect 32175 2468 32220 2496
rect 32214 2456 32220 2468
rect 32272 2456 32278 2508
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 33597 2499 33655 2505
rect 33597 2496 33609 2499
rect 33192 2468 33609 2496
rect 33192 2456 33198 2468
rect 33597 2465 33609 2468
rect 33643 2465 33655 2499
rect 33778 2496 33784 2508
rect 33739 2468 33784 2496
rect 33597 2459 33655 2465
rect 33778 2456 33784 2468
rect 33836 2456 33842 2508
rect 34514 2456 34520 2508
rect 34572 2496 34578 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 34572 2468 34713 2496
rect 34572 2456 34578 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 34790 2456 34796 2508
rect 34848 2496 34854 2508
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 34848 2468 34897 2496
rect 34848 2456 34854 2468
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 34885 2459 34943 2465
rect 36170 2456 36176 2508
rect 36228 2496 36234 2508
rect 36449 2499 36507 2505
rect 36449 2496 36461 2499
rect 36228 2468 36461 2496
rect 36228 2456 36234 2468
rect 36449 2465 36461 2468
rect 36495 2465 36507 2499
rect 36449 2459 36507 2465
rect 38746 2456 38752 2508
rect 38804 2496 38810 2508
rect 38933 2499 38991 2505
rect 38933 2496 38945 2499
rect 38804 2468 38945 2496
rect 38804 2456 38810 2468
rect 38933 2465 38945 2468
rect 38979 2465 38991 2499
rect 38933 2459 38991 2465
rect 39022 2456 39028 2508
rect 39080 2496 39086 2508
rect 39117 2499 39175 2505
rect 39117 2496 39129 2499
rect 39080 2468 39129 2496
rect 39080 2456 39086 2468
rect 39117 2465 39129 2468
rect 39163 2465 39175 2499
rect 40034 2496 40040 2508
rect 39995 2468 40040 2496
rect 39117 2459 39175 2465
rect 40034 2456 40040 2468
rect 40092 2456 40098 2508
rect 40218 2496 40224 2508
rect 40179 2468 40224 2496
rect 40218 2456 40224 2468
rect 40276 2456 40282 2508
rect 41598 2496 41604 2508
rect 41559 2468 41604 2496
rect 41598 2456 41604 2468
rect 41656 2456 41662 2508
rect 41782 2496 41788 2508
rect 41743 2468 41788 2496
rect 41782 2456 41788 2468
rect 41840 2456 41846 2508
rect 42702 2496 42708 2508
rect 42663 2468 42708 2496
rect 42702 2456 42708 2468
rect 42760 2456 42766 2508
rect 42886 2496 42892 2508
rect 42847 2468 42892 2496
rect 42886 2456 42892 2468
rect 42944 2456 42950 2508
rect 44174 2456 44180 2508
rect 44232 2496 44238 2508
rect 44269 2499 44327 2505
rect 44269 2496 44281 2499
rect 44232 2468 44281 2496
rect 44232 2456 44238 2468
rect 44269 2465 44281 2468
rect 44315 2465 44327 2499
rect 44269 2459 44327 2465
rect 44358 2456 44364 2508
rect 44416 2496 44422 2508
rect 44453 2499 44511 2505
rect 44453 2496 44465 2499
rect 44416 2468 44465 2496
rect 44416 2456 44422 2468
rect 44453 2465 44465 2468
rect 44499 2465 44511 2499
rect 44453 2459 44511 2465
rect 45094 2456 45100 2508
rect 45152 2496 45158 2508
rect 45373 2499 45431 2505
rect 45373 2496 45385 2499
rect 45152 2468 45385 2496
rect 45152 2456 45158 2468
rect 45373 2465 45385 2468
rect 45419 2465 45431 2499
rect 45373 2459 45431 2465
rect 45554 2456 45560 2508
rect 45612 2496 45618 2508
rect 46934 2496 46940 2508
rect 45612 2468 45657 2496
rect 46895 2468 46940 2496
rect 45612 2456 45618 2468
rect 46934 2456 46940 2468
rect 46992 2456 46998 2508
rect 47121 2499 47179 2505
rect 47121 2465 47133 2499
rect 47167 2496 47179 2499
rect 47210 2496 47216 2508
rect 47167 2468 47216 2496
rect 47167 2465 47179 2468
rect 47121 2459 47179 2465
rect 47210 2456 47216 2468
rect 47268 2456 47274 2508
rect 48774 2456 48780 2508
rect 48832 2496 48838 2508
rect 49605 2499 49663 2505
rect 49605 2496 49617 2499
rect 48832 2468 49617 2496
rect 48832 2456 48838 2468
rect 49605 2465 49617 2468
rect 49651 2465 49663 2499
rect 49605 2459 49663 2465
rect 49694 2456 49700 2508
rect 49752 2496 49758 2508
rect 49789 2499 49847 2505
rect 49789 2496 49801 2499
rect 49752 2468 49801 2496
rect 49752 2456 49758 2468
rect 49789 2465 49801 2468
rect 49835 2465 49847 2499
rect 49789 2459 49847 2465
rect 31110 2428 31116 2440
rect 31071 2400 31116 2428
rect 31110 2388 31116 2400
rect 31168 2388 31174 2440
rect 36262 2428 36268 2440
rect 36223 2400 36268 2428
rect 36262 2388 36268 2400
rect 36320 2388 36326 2440
rect 43530 2388 43536 2440
rect 43588 2428 43594 2440
rect 50709 2431 50767 2437
rect 43588 2400 46888 2428
rect 43588 2388 43594 2400
rect 31297 2363 31355 2369
rect 31297 2360 31309 2363
rect 30576 2332 31309 2360
rect 31297 2329 31309 2332
rect 31343 2329 31355 2363
rect 31297 2323 31355 2329
rect 31938 2320 31944 2372
rect 31996 2360 32002 2372
rect 32401 2363 32459 2369
rect 32401 2360 32413 2363
rect 31996 2332 32413 2360
rect 31996 2320 32002 2332
rect 32401 2329 32413 2332
rect 32447 2329 32459 2363
rect 32401 2323 32459 2329
rect 33318 2320 33324 2372
rect 33376 2360 33382 2372
rect 33965 2363 34023 2369
rect 33965 2360 33977 2363
rect 33376 2332 33977 2360
rect 33376 2320 33382 2332
rect 33965 2329 33977 2332
rect 34011 2329 34023 2363
rect 33965 2323 34023 2329
rect 38013 2363 38071 2369
rect 38013 2329 38025 2363
rect 38059 2360 38071 2363
rect 39758 2360 39764 2372
rect 38059 2332 39764 2360
rect 38059 2329 38071 2332
rect 38013 2323 38071 2329
rect 39758 2320 39764 2332
rect 39816 2320 39822 2372
rect 41966 2360 41972 2372
rect 41927 2332 41972 2360
rect 41966 2320 41972 2332
rect 42024 2320 42030 2372
rect 43070 2360 43076 2372
rect 43031 2332 43076 2360
rect 43070 2320 43076 2332
rect 43128 2320 43134 2372
rect 45186 2320 45192 2372
rect 45244 2360 45250 2372
rect 46860 2360 46888 2400
rect 50709 2397 50721 2431
rect 50755 2428 50767 2431
rect 50798 2428 50804 2440
rect 50755 2400 50804 2428
rect 50755 2397 50767 2400
rect 50709 2391 50767 2397
rect 50798 2388 50804 2400
rect 50856 2388 50862 2440
rect 50908 2437 50936 2536
rect 51000 2536 53604 2564
rect 50893 2431 50951 2437
rect 50893 2397 50905 2431
rect 50939 2397 50951 2431
rect 50893 2391 50951 2397
rect 48317 2363 48375 2369
rect 48317 2360 48329 2363
rect 45244 2332 45554 2360
rect 46860 2332 48329 2360
rect 45244 2320 45250 2332
rect 2958 2292 2964 2304
rect 2919 2264 2964 2292
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 29181 2295 29239 2301
rect 29181 2261 29193 2295
rect 29227 2292 29239 2295
rect 31386 2292 31392 2304
rect 29227 2264 31392 2292
rect 29227 2261 29239 2264
rect 29181 2255 29239 2261
rect 31386 2252 31392 2264
rect 31444 2252 31450 2304
rect 45526 2292 45554 2332
rect 48317 2329 48329 2332
rect 48363 2329 48375 2363
rect 48317 2323 48375 2329
rect 49510 2320 49516 2372
rect 49568 2360 49574 2372
rect 51000 2360 51028 2536
rect 51350 2456 51356 2508
rect 51408 2496 51414 2508
rect 53576 2505 53604 2536
rect 54496 2536 55220 2564
rect 52273 2499 52331 2505
rect 52273 2496 52285 2499
rect 51408 2468 52285 2496
rect 51408 2456 51414 2468
rect 52273 2465 52285 2468
rect 52319 2465 52331 2499
rect 53377 2499 53435 2505
rect 53377 2496 53389 2499
rect 52273 2459 52331 2465
rect 52380 2468 53389 2496
rect 51810 2388 51816 2440
rect 51868 2428 51874 2440
rect 52380 2428 52408 2468
rect 53377 2465 53389 2468
rect 53423 2465 53435 2499
rect 53377 2459 53435 2465
rect 53561 2499 53619 2505
rect 53561 2465 53573 2499
rect 53607 2465 53619 2499
rect 53561 2459 53619 2465
rect 51868 2400 52408 2428
rect 52457 2431 52515 2437
rect 51868 2388 51874 2400
rect 52457 2397 52469 2431
rect 52503 2397 52515 2431
rect 52457 2391 52515 2397
rect 49568 2332 51028 2360
rect 49568 2320 49574 2332
rect 51166 2320 51172 2372
rect 51224 2360 51230 2372
rect 52472 2360 52500 2391
rect 52638 2360 52644 2372
rect 51224 2332 52500 2360
rect 52599 2332 52644 2360
rect 51224 2320 51230 2332
rect 52638 2320 52644 2332
rect 52696 2320 52702 2372
rect 54496 2292 54524 2536
rect 55214 2524 55220 2536
rect 55272 2524 55278 2576
rect 57974 2564 57980 2576
rect 57935 2536 57980 2564
rect 57974 2524 57980 2536
rect 58032 2524 58038 2576
rect 55306 2456 55312 2508
rect 55364 2496 55370 2508
rect 56045 2499 56103 2505
rect 56045 2496 56057 2499
rect 55364 2468 56057 2496
rect 55364 2456 55370 2468
rect 56045 2465 56057 2468
rect 56091 2465 56103 2499
rect 56045 2459 56103 2465
rect 54941 2431 54999 2437
rect 54941 2397 54953 2431
rect 54987 2397 54999 2431
rect 55122 2428 55128 2440
rect 55083 2400 55128 2428
rect 54941 2391 54999 2397
rect 45526 2264 54524 2292
rect 54662 2252 54668 2304
rect 54720 2292 54726 2304
rect 54757 2295 54815 2301
rect 54757 2292 54769 2295
rect 54720 2264 54769 2292
rect 54720 2252 54726 2264
rect 54757 2261 54769 2264
rect 54803 2292 54815 2295
rect 54956 2292 54984 2391
rect 55122 2388 55128 2400
rect 55180 2388 55186 2440
rect 56226 2428 56232 2440
rect 56187 2400 56232 2428
rect 56226 2388 56232 2400
rect 56284 2388 56290 2440
rect 54803 2264 54984 2292
rect 54803 2261 54815 2264
rect 54757 2255 54815 2261
rect 57882 2252 57888 2304
rect 57940 2292 57946 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 57940 2264 58081 2292
rect 57940 2252 57946 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 58880 2202
rect 1104 2128 58880 2150
rect 44910 2048 44916 2100
rect 44968 2088 44974 2100
rect 54662 2088 54668 2100
rect 44968 2060 54668 2088
rect 44968 2048 44974 2060
rect 54662 2048 54668 2060
rect 54720 2048 54726 2100
rect 47670 1980 47676 2032
rect 47728 2020 47734 2032
rect 51166 2020 51172 2032
rect 47728 1992 51172 2020
rect 47728 1980 47734 1992
rect 51166 1980 51172 1992
rect 51224 1980 51230 2032
rect 48130 1912 48136 1964
rect 48188 1952 48194 1964
rect 55122 1952 55128 1964
rect 48188 1924 55128 1952
rect 48188 1912 48194 1924
rect 55122 1912 55128 1924
rect 55180 1912 55186 1964
rect 49418 1844 49424 1896
rect 49476 1884 49482 1896
rect 56226 1884 56232 1896
rect 49476 1856 56232 1884
rect 49476 1844 49482 1856
rect 56226 1844 56232 1856
rect 56284 1844 56290 1896
rect 54478 1640 54484 1692
rect 54536 1680 54542 1692
rect 56686 1680 56692 1692
rect 54536 1652 56692 1680
rect 54536 1640 54542 1652
rect 56686 1640 56692 1652
rect 56744 1640 56750 1692
rect 44082 1300 44088 1352
rect 44140 1340 44146 1352
rect 55214 1340 55220 1352
rect 44140 1312 55220 1340
rect 44140 1300 44146 1312
rect 55214 1300 55220 1312
rect 55272 1300 55278 1352
<< via1 >>
rect 55220 58284 55272 58336
rect 56416 58284 56468 58336
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 59544 57536 59596 57588
rect 4620 57468 4672 57520
rect 24032 57468 24084 57520
rect 6644 57400 6696 57452
rect 1400 57375 1452 57384
rect 1400 57341 1409 57375
rect 1409 57341 1443 57375
rect 1443 57341 1452 57375
rect 1400 57332 1452 57341
rect 2044 57375 2096 57384
rect 2044 57341 2053 57375
rect 2053 57341 2087 57375
rect 2087 57341 2096 57375
rect 2044 57332 2096 57341
rect 2780 57332 2832 57384
rect 5080 57375 5132 57384
rect 5080 57341 5089 57375
rect 5089 57341 5123 57375
rect 5123 57341 5132 57375
rect 5080 57332 5132 57341
rect 5908 57332 5960 57384
rect 14556 57400 14608 57452
rect 7472 57332 7524 57384
rect 8208 57375 8260 57384
rect 8208 57341 8217 57375
rect 8217 57341 8251 57375
rect 8251 57341 8260 57375
rect 8208 57332 8260 57341
rect 9036 57332 9088 57384
rect 9772 57332 9824 57384
rect 10600 57332 10652 57384
rect 11428 57332 11480 57384
rect 12440 57332 12492 57384
rect 12992 57332 13044 57384
rect 13820 57332 13872 57384
rect 15384 57400 15436 57452
rect 20076 57400 20128 57452
rect 16948 57332 17000 57384
rect 17684 57332 17736 57384
rect 18512 57332 18564 57384
rect 19340 57332 19392 57384
rect 22468 57400 22520 57452
rect 20996 57332 21048 57384
rect 21640 57332 21692 57384
rect 23204 57400 23256 57452
rect 31944 57468 31996 57520
rect 25688 57400 25740 57452
rect 27988 57400 28040 57452
rect 4620 57264 4672 57316
rect 5080 57196 5132 57248
rect 24860 57196 24912 57248
rect 27160 57332 27212 57384
rect 30380 57400 30432 57452
rect 29000 57332 29052 57384
rect 29644 57332 29696 57384
rect 31116 57400 31168 57452
rect 55036 57468 55088 57520
rect 55496 57511 55548 57520
rect 55496 57477 55505 57511
rect 55505 57477 55539 57511
rect 55539 57477 55548 57511
rect 55496 57468 55548 57477
rect 33508 57400 33560 57452
rect 36636 57400 36688 57452
rect 32680 57264 32732 57316
rect 35256 57332 35308 57384
rect 39028 57400 39080 57452
rect 35900 57264 35952 57316
rect 37648 57332 37700 57384
rect 45376 57400 45428 57452
rect 42156 57375 42208 57384
rect 38200 57264 38252 57316
rect 42156 57341 42165 57375
rect 42165 57341 42199 57375
rect 42199 57341 42208 57375
rect 42156 57332 42208 57341
rect 42984 57375 43036 57384
rect 42984 57341 42993 57375
rect 42993 57341 43027 57375
rect 43027 57341 43036 57375
rect 42984 57332 43036 57341
rect 43720 57332 43772 57384
rect 44548 57332 44600 57384
rect 49240 57400 49292 57452
rect 46112 57332 46164 57384
rect 47032 57332 47084 57384
rect 47676 57332 47728 57384
rect 48504 57332 48556 57384
rect 50068 57400 50120 57452
rect 54944 57400 54996 57452
rect 55404 57332 55456 57384
rect 53104 57307 53156 57316
rect 53104 57273 53113 57307
rect 53113 57273 53147 57307
rect 53147 57273 53156 57307
rect 53104 57264 53156 57273
rect 53840 57307 53892 57316
rect 53840 57273 53849 57307
rect 53849 57273 53883 57307
rect 53883 57273 53892 57307
rect 53840 57264 53892 57273
rect 55772 57264 55824 57316
rect 57980 57307 58032 57316
rect 57980 57273 57989 57307
rect 57989 57273 58023 57307
rect 58023 57273 58032 57307
rect 57980 57264 58032 57273
rect 58164 57307 58216 57316
rect 58164 57273 58173 57307
rect 58173 57273 58207 57307
rect 58207 57273 58216 57307
rect 58164 57264 58216 57273
rect 58072 57196 58124 57248
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 50326 57094 50378 57146
rect 50390 57094 50442 57146
rect 50454 57094 50506 57146
rect 50518 57094 50570 57146
rect 53104 56992 53156 57044
rect 56600 56992 56652 57044
rect 57980 56992 58032 57044
rect 1400 56899 1452 56908
rect 1400 56865 1409 56899
rect 1409 56865 1443 56899
rect 1443 56865 1452 56899
rect 1400 56856 1452 56865
rect 2688 56856 2740 56908
rect 16120 56899 16172 56908
rect 16120 56865 16129 56899
rect 16129 56865 16163 56899
rect 16163 56865 16172 56899
rect 16120 56856 16172 56865
rect 26424 56899 26476 56908
rect 26424 56865 26433 56899
rect 26433 56865 26467 56899
rect 26467 56865 26476 56899
rect 26424 56856 26476 56865
rect 34244 56899 34296 56908
rect 34244 56865 34253 56899
rect 34253 56865 34287 56899
rect 34287 56865 34296 56899
rect 34244 56856 34296 56865
rect 39764 56899 39816 56908
rect 39764 56865 39773 56899
rect 39773 56865 39807 56899
rect 39807 56865 39816 56899
rect 39764 56856 39816 56865
rect 40592 56856 40644 56908
rect 41420 56856 41472 56908
rect 51080 56856 51132 56908
rect 51632 56856 51684 56908
rect 52460 56856 52512 56908
rect 55588 56856 55640 56908
rect 55772 56899 55824 56908
rect 55772 56865 55781 56899
rect 55781 56865 55815 56899
rect 55815 56865 55824 56899
rect 55772 56856 55824 56865
rect 57980 56856 58032 56908
rect 4712 56831 4764 56840
rect 4712 56797 4721 56831
rect 4721 56797 4755 56831
rect 4755 56797 4764 56831
rect 4712 56788 4764 56797
rect 53840 56788 53892 56840
rect 5448 56720 5500 56772
rect 56140 56720 56192 56772
rect 56324 56788 56376 56840
rect 57612 56788 57664 56840
rect 56876 56720 56928 56772
rect 57060 56763 57112 56772
rect 57060 56729 57069 56763
rect 57069 56729 57103 56763
rect 57103 56729 57112 56763
rect 57060 56720 57112 56729
rect 3332 56695 3384 56704
rect 3332 56661 3341 56695
rect 3341 56661 3375 56695
rect 3375 56661 3384 56695
rect 3332 56652 3384 56661
rect 57704 56652 57756 56704
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 388 56448 440 56500
rect 1308 56448 1360 56500
rect 4620 56448 4672 56500
rect 4712 56448 4764 56500
rect 5448 56491 5500 56500
rect 5448 56457 5457 56491
rect 5457 56457 5491 56491
rect 5491 56457 5500 56491
rect 5448 56448 5500 56457
rect 53932 56448 53984 56500
rect 54760 56448 54812 56500
rect 56324 56448 56376 56500
rect 56600 56491 56652 56500
rect 56600 56457 56609 56491
rect 56609 56457 56643 56491
rect 56643 56457 56652 56491
rect 56600 56448 56652 56457
rect 58072 56491 58124 56500
rect 58072 56457 58081 56491
rect 58081 56457 58115 56491
rect 58115 56457 58124 56491
rect 58072 56448 58124 56457
rect 3332 56312 3384 56364
rect 55404 56380 55456 56432
rect 1124 56244 1176 56296
rect 1952 56244 2004 56296
rect 55128 56312 55180 56364
rect 56232 56380 56284 56432
rect 58256 56380 58308 56432
rect 56876 56312 56928 56364
rect 57704 56355 57756 56364
rect 57704 56321 57713 56355
rect 57713 56321 57747 56355
rect 57747 56321 57756 56355
rect 57704 56312 57756 56321
rect 3700 56176 3752 56228
rect 53196 56244 53248 56296
rect 55772 56244 55824 56296
rect 56140 56287 56192 56296
rect 56140 56253 56149 56287
rect 56149 56253 56183 56287
rect 56183 56253 56192 56287
rect 56140 56244 56192 56253
rect 57152 56176 57204 56228
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 50326 56006 50378 56058
rect 50390 56006 50442 56058
rect 50454 56006 50506 56058
rect 50518 56006 50570 56058
rect 57612 55904 57664 55956
rect 1400 55811 1452 55820
rect 1400 55777 1409 55811
rect 1409 55777 1443 55811
rect 1443 55777 1452 55811
rect 1400 55768 1452 55777
rect 3516 55768 3568 55820
rect 54024 55768 54076 55820
rect 55680 55768 55732 55820
rect 55772 55811 55824 55820
rect 55772 55777 55781 55811
rect 55781 55777 55815 55811
rect 55815 55777 55824 55811
rect 55772 55768 55824 55777
rect 55312 55700 55364 55752
rect 58256 55836 58308 55888
rect 57336 55768 57388 55820
rect 56508 55700 56560 55752
rect 58716 55700 58768 55752
rect 58164 55675 58216 55684
rect 58164 55641 58173 55675
rect 58173 55641 58207 55675
rect 58207 55641 58216 55675
rect 58164 55632 58216 55641
rect 55496 55564 55548 55616
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 57244 55224 57296 55276
rect 53932 55156 53984 55208
rect 56324 55199 56376 55208
rect 56324 55165 56333 55199
rect 56333 55165 56367 55199
rect 56367 55165 56376 55199
rect 56324 55156 56376 55165
rect 56600 55156 56652 55208
rect 57980 55156 58032 55208
rect 56876 55131 56928 55140
rect 56876 55097 56885 55131
rect 56885 55097 56919 55131
rect 56919 55097 56928 55131
rect 56876 55088 56928 55097
rect 57060 55131 57112 55140
rect 57060 55097 57069 55131
rect 57069 55097 57103 55131
rect 57103 55097 57112 55131
rect 57060 55088 57112 55097
rect 56140 55063 56192 55072
rect 56140 55029 56149 55063
rect 56149 55029 56183 55063
rect 56183 55029 56192 55063
rect 56140 55020 56192 55029
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 50326 54918 50378 54970
rect 50390 54918 50442 54970
rect 50454 54918 50506 54970
rect 50518 54918 50570 54970
rect 55772 54859 55824 54868
rect 55772 54825 55781 54859
rect 55781 54825 55815 54859
rect 55815 54825 55824 54859
rect 55772 54816 55824 54825
rect 56324 54816 56376 54868
rect 57336 54859 57388 54868
rect 57336 54825 57345 54859
rect 57345 54825 57379 54859
rect 57379 54825 57388 54859
rect 57336 54816 57388 54825
rect 1400 54723 1452 54732
rect 1400 54689 1409 54723
rect 1409 54689 1443 54723
rect 1443 54689 1452 54723
rect 1400 54680 1452 54689
rect 56232 54748 56284 54800
rect 55312 54680 55364 54732
rect 56140 54680 56192 54732
rect 57980 54723 58032 54732
rect 57980 54689 57989 54723
rect 57989 54689 58023 54723
rect 58023 54689 58032 54723
rect 57980 54680 58032 54689
rect 55496 54612 55548 54664
rect 56324 54544 56376 54596
rect 58164 54587 58216 54596
rect 58164 54553 58173 54587
rect 58173 54553 58207 54587
rect 58207 54553 58216 54587
rect 58164 54544 58216 54553
rect 54944 54519 54996 54528
rect 54944 54485 54953 54519
rect 54953 54485 54987 54519
rect 54987 54485 54996 54519
rect 54944 54476 54996 54485
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 56600 54272 56652 54324
rect 56876 54272 56928 54324
rect 54944 54136 54996 54188
rect 55496 54111 55548 54120
rect 55496 54077 55505 54111
rect 55505 54077 55539 54111
rect 55539 54077 55548 54111
rect 55496 54068 55548 54077
rect 56324 54111 56376 54120
rect 56324 54077 56333 54111
rect 56333 54077 56367 54111
rect 56367 54077 56376 54111
rect 56324 54068 56376 54077
rect 57244 54136 57296 54188
rect 57428 54000 57480 54052
rect 56968 53975 57020 53984
rect 56968 53941 56977 53975
rect 56977 53941 57011 53975
rect 57011 53941 57020 53975
rect 56968 53932 57020 53941
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 50326 53830 50378 53882
rect 50390 53830 50442 53882
rect 50454 53830 50506 53882
rect 50518 53830 50570 53882
rect 1400 53635 1452 53644
rect 1400 53601 1409 53635
rect 1409 53601 1443 53635
rect 1443 53601 1452 53635
rect 1400 53592 1452 53601
rect 55588 53635 55640 53644
rect 55588 53601 55597 53635
rect 55597 53601 55631 53635
rect 55631 53601 55640 53635
rect 55588 53592 55640 53601
rect 56416 53524 56468 53576
rect 57244 53567 57296 53576
rect 57244 53533 57253 53567
rect 57253 53533 57287 53567
rect 57287 53533 57296 53567
rect 57244 53524 57296 53533
rect 57428 53499 57480 53508
rect 57428 53465 57437 53499
rect 57437 53465 57471 53499
rect 57471 53465 57480 53499
rect 57428 53456 57480 53465
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 56416 53227 56468 53236
rect 56416 53193 56425 53227
rect 56425 53193 56459 53227
rect 56459 53193 56468 53227
rect 56416 53184 56468 53193
rect 57244 53184 57296 53236
rect 57980 53227 58032 53236
rect 57980 53193 57989 53227
rect 57989 53193 58023 53227
rect 58023 53193 58032 53227
rect 57980 53184 58032 53193
rect 1400 53023 1452 53032
rect 1400 52989 1409 53023
rect 1409 52989 1443 53023
rect 1443 52989 1452 53023
rect 1400 52980 1452 52989
rect 56324 52980 56376 53032
rect 57244 52980 57296 53032
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 50326 52742 50378 52794
rect 50390 52742 50442 52794
rect 50454 52742 50506 52794
rect 50518 52742 50570 52794
rect 57244 52683 57296 52692
rect 57244 52649 57253 52683
rect 57253 52649 57287 52683
rect 57287 52649 57296 52683
rect 57244 52640 57296 52649
rect 57428 52547 57480 52556
rect 57428 52513 57437 52547
rect 57437 52513 57471 52547
rect 57471 52513 57480 52547
rect 57428 52504 57480 52513
rect 57980 52547 58032 52556
rect 57980 52513 57989 52547
rect 57989 52513 58023 52547
rect 58023 52513 58032 52547
rect 57980 52504 58032 52513
rect 57888 52436 57940 52488
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 57980 52139 58032 52148
rect 57980 52105 57989 52139
rect 57989 52105 58023 52139
rect 58023 52105 58032 52139
rect 57980 52096 58032 52105
rect 1400 51935 1452 51944
rect 1400 51901 1409 51935
rect 1409 51901 1443 51935
rect 1443 51901 1452 51935
rect 1400 51892 1452 51901
rect 55496 51935 55548 51944
rect 55496 51901 55505 51935
rect 55505 51901 55539 51935
rect 55539 51901 55548 51935
rect 55496 51892 55548 51901
rect 57520 51935 57572 51944
rect 56876 51867 56928 51876
rect 56876 51833 56885 51867
rect 56885 51833 56919 51867
rect 56919 51833 56928 51867
rect 56876 51824 56928 51833
rect 57060 51867 57112 51876
rect 57060 51833 57069 51867
rect 57069 51833 57103 51867
rect 57103 51833 57112 51867
rect 57060 51824 57112 51833
rect 57520 51901 57529 51935
rect 57529 51901 57563 51935
rect 57563 51901 57572 51935
rect 57520 51892 57572 51901
rect 57428 51824 57480 51876
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 50326 51654 50378 51706
rect 50390 51654 50442 51706
rect 50454 51654 50506 51706
rect 50518 51654 50570 51706
rect 56876 51552 56928 51604
rect 57520 51416 57572 51468
rect 57244 51391 57296 51400
rect 57244 51357 57253 51391
rect 57253 51357 57287 51391
rect 57287 51357 57296 51391
rect 57244 51348 57296 51357
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 57244 51008 57296 51060
rect 1400 50847 1452 50856
rect 1400 50813 1409 50847
rect 1409 50813 1443 50847
rect 1443 50813 1452 50847
rect 1400 50804 1452 50813
rect 56324 50804 56376 50856
rect 57428 50847 57480 50856
rect 57428 50813 57437 50847
rect 57437 50813 57471 50847
rect 57471 50813 57480 50847
rect 57428 50804 57480 50813
rect 57520 50736 57572 50788
rect 57980 50779 58032 50788
rect 57980 50745 57989 50779
rect 57989 50745 58023 50779
rect 58023 50745 58032 50779
rect 57980 50736 58032 50745
rect 58164 50779 58216 50788
rect 58164 50745 58173 50779
rect 58173 50745 58207 50779
rect 58207 50745 58216 50779
rect 58164 50736 58216 50745
rect 57704 50668 57756 50720
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 50326 50566 50378 50618
rect 50390 50566 50442 50618
rect 50454 50566 50506 50618
rect 50518 50566 50570 50618
rect 57980 50464 58032 50516
rect 1400 50371 1452 50380
rect 1400 50337 1409 50371
rect 1409 50337 1443 50371
rect 1443 50337 1452 50371
rect 1400 50328 1452 50337
rect 56876 50371 56928 50380
rect 56876 50337 56885 50371
rect 56885 50337 56919 50371
rect 56919 50337 56928 50371
rect 56876 50328 56928 50337
rect 57520 50371 57572 50380
rect 57520 50337 57529 50371
rect 57529 50337 57563 50371
rect 57563 50337 57572 50371
rect 57520 50328 57572 50337
rect 57704 50371 57756 50380
rect 57704 50337 57713 50371
rect 57713 50337 57747 50371
rect 57747 50337 57756 50371
rect 57704 50328 57756 50337
rect 57060 50235 57112 50244
rect 57060 50201 57069 50235
rect 57069 50201 57103 50235
rect 57103 50201 57112 50235
rect 57060 50192 57112 50201
rect 57152 50124 57204 50176
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 56324 49920 56376 49972
rect 56876 49920 56928 49972
rect 55956 49784 56008 49836
rect 57152 49827 57204 49836
rect 55220 49759 55272 49768
rect 55220 49725 55229 49759
rect 55229 49725 55263 49759
rect 55263 49725 55272 49759
rect 55220 49716 55272 49725
rect 56324 49716 56376 49768
rect 57152 49793 57161 49827
rect 57161 49793 57195 49827
rect 57195 49793 57204 49827
rect 57152 49784 57204 49793
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 50326 49478 50378 49530
rect 50390 49478 50442 49530
rect 50454 49478 50506 49530
rect 50518 49478 50570 49530
rect 1400 49283 1452 49292
rect 1400 49249 1409 49283
rect 1409 49249 1443 49283
rect 1443 49249 1452 49283
rect 1400 49240 1452 49249
rect 57428 49283 57480 49292
rect 57428 49249 57437 49283
rect 57437 49249 57471 49283
rect 57471 49249 57480 49283
rect 57428 49240 57480 49249
rect 57796 49240 57848 49292
rect 57980 49283 58032 49292
rect 57980 49249 57989 49283
rect 57989 49249 58023 49283
rect 58023 49249 58032 49283
rect 57980 49240 58032 49249
rect 58164 49283 58216 49292
rect 58164 49249 58173 49283
rect 58173 49249 58207 49283
rect 58207 49249 58216 49283
rect 58164 49240 58216 49249
rect 55772 49079 55824 49088
rect 55772 49045 55781 49079
rect 55781 49045 55815 49079
rect 55815 49045 55824 49079
rect 55772 49036 55824 49045
rect 57704 49036 57756 49088
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 57980 48875 58032 48884
rect 57980 48841 57989 48875
rect 57989 48841 58023 48875
rect 58023 48841 58032 48875
rect 57980 48832 58032 48841
rect 57060 48807 57112 48816
rect 57060 48773 57069 48807
rect 57069 48773 57103 48807
rect 57103 48773 57112 48807
rect 57060 48764 57112 48773
rect 55772 48696 55824 48748
rect 57704 48739 57756 48748
rect 57704 48705 57713 48739
rect 57713 48705 57747 48739
rect 57747 48705 57756 48739
rect 57704 48696 57756 48705
rect 55496 48671 55548 48680
rect 55496 48637 55505 48671
rect 55505 48637 55539 48671
rect 55539 48637 55548 48671
rect 55496 48628 55548 48637
rect 57060 48628 57112 48680
rect 57428 48560 57480 48612
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 50326 48390 50378 48442
rect 50390 48390 50442 48442
rect 50454 48390 50506 48442
rect 50518 48390 50570 48442
rect 1400 48195 1452 48204
rect 1400 48161 1409 48195
rect 1409 48161 1443 48195
rect 1443 48161 1452 48195
rect 1400 48152 1452 48161
rect 57060 48195 57112 48204
rect 57060 48161 57069 48195
rect 57069 48161 57103 48195
rect 57103 48161 57112 48195
rect 57060 48152 57112 48161
rect 55496 48084 55548 48136
rect 57428 48059 57480 48068
rect 57428 48025 57437 48059
rect 57437 48025 57471 48059
rect 57471 48025 57480 48059
rect 57428 48016 57480 48025
rect 57520 47948 57572 48000
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 55496 47787 55548 47796
rect 55496 47753 55505 47787
rect 55505 47753 55539 47787
rect 55539 47753 55548 47787
rect 55496 47744 55548 47753
rect 57060 47651 57112 47660
rect 57060 47617 57069 47651
rect 57069 47617 57103 47651
rect 57103 47617 57112 47651
rect 57060 47608 57112 47617
rect 57520 47651 57572 47660
rect 57520 47617 57529 47651
rect 57529 47617 57563 47651
rect 57563 47617 57572 47651
rect 57520 47608 57572 47617
rect 55680 47583 55732 47592
rect 55680 47549 55689 47583
rect 55689 47549 55723 47583
rect 55723 47549 55732 47583
rect 55680 47540 55732 47549
rect 57796 47540 57848 47592
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 50326 47302 50378 47354
rect 50390 47302 50442 47354
rect 50454 47302 50506 47354
rect 50518 47302 50570 47354
rect 1400 47107 1452 47116
rect 1400 47073 1409 47107
rect 1409 47073 1443 47107
rect 1443 47073 1452 47107
rect 1400 47064 1452 47073
rect 55220 47064 55272 47116
rect 55956 47064 56008 47116
rect 57244 47107 57296 47116
rect 57244 47073 57253 47107
rect 57253 47073 57287 47107
rect 57287 47073 57296 47107
rect 57244 47064 57296 47073
rect 57428 47107 57480 47116
rect 57428 47073 57437 47107
rect 57437 47073 57471 47107
rect 57471 47073 57480 47107
rect 57428 47064 57480 47073
rect 57980 47107 58032 47116
rect 57980 47073 57989 47107
rect 57989 47073 58023 47107
rect 58023 47073 58032 47107
rect 57980 47064 58032 47073
rect 57520 46928 57572 46980
rect 57888 46928 57940 46980
rect 55680 46860 55732 46912
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 57244 46656 57296 46708
rect 55036 46520 55088 46572
rect 58256 46520 58308 46572
rect 1400 46495 1452 46504
rect 1400 46461 1409 46495
rect 1409 46461 1443 46495
rect 1443 46461 1452 46495
rect 1400 46452 1452 46461
rect 54760 46452 54812 46504
rect 55680 46452 55732 46504
rect 57612 46427 57664 46436
rect 57612 46393 57621 46427
rect 57621 46393 57655 46427
rect 57655 46393 57664 46427
rect 57612 46384 57664 46393
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 50326 46214 50378 46266
rect 50390 46214 50442 46266
rect 50454 46214 50506 46266
rect 50518 46214 50570 46266
rect 55036 46155 55088 46164
rect 55036 46121 55045 46155
rect 55045 46121 55079 46155
rect 55079 46121 55088 46155
rect 55036 46112 55088 46121
rect 57612 46112 57664 46164
rect 57796 46112 57848 46164
rect 54944 46019 54996 46028
rect 54944 45985 54953 46019
rect 54953 45985 54987 46019
rect 54987 45985 54996 46019
rect 54944 45976 54996 45985
rect 55772 46019 55824 46028
rect 55036 45908 55088 45960
rect 51540 45840 51592 45892
rect 55772 45985 55781 46019
rect 55781 45985 55815 46019
rect 55815 45985 55824 46019
rect 55772 45976 55824 45985
rect 55956 45976 56008 46028
rect 58256 45976 58308 46028
rect 55772 45840 55824 45892
rect 56508 45772 56560 45824
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 57060 45543 57112 45552
rect 57060 45509 57069 45543
rect 57069 45509 57103 45543
rect 57103 45509 57112 45543
rect 57060 45500 57112 45509
rect 57980 45543 58032 45552
rect 57980 45509 57989 45543
rect 57989 45509 58023 45543
rect 58023 45509 58032 45543
rect 57980 45500 58032 45509
rect 57520 45475 57572 45484
rect 57520 45441 57529 45475
rect 57529 45441 57563 45475
rect 57563 45441 57572 45475
rect 57520 45432 57572 45441
rect 1400 45407 1452 45416
rect 1400 45373 1409 45407
rect 1409 45373 1443 45407
rect 1443 45373 1452 45407
rect 1400 45364 1452 45373
rect 53932 45364 53984 45416
rect 54208 45407 54260 45416
rect 54208 45373 54217 45407
rect 54217 45373 54251 45407
rect 54251 45373 54260 45407
rect 54208 45364 54260 45373
rect 52920 45296 52972 45348
rect 54944 45364 54996 45416
rect 55128 45364 55180 45416
rect 55680 45407 55732 45416
rect 55680 45373 55689 45407
rect 55689 45373 55723 45407
rect 55723 45373 55732 45407
rect 55680 45364 55732 45373
rect 57612 45364 57664 45416
rect 58072 45364 58124 45416
rect 57336 45296 57388 45348
rect 54116 45271 54168 45280
rect 54116 45237 54125 45271
rect 54125 45237 54159 45271
rect 54159 45237 54168 45271
rect 54116 45228 54168 45237
rect 55404 45228 55456 45280
rect 56048 45228 56100 45280
rect 57704 45228 57756 45280
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 50326 45126 50378 45178
rect 50390 45126 50442 45178
rect 50454 45126 50506 45178
rect 50518 45126 50570 45178
rect 52736 45024 52788 45076
rect 57336 45067 57388 45076
rect 57336 45033 57345 45067
rect 57345 45033 57379 45067
rect 57379 45033 57388 45067
rect 57336 45024 57388 45033
rect 52092 44888 52144 44940
rect 54208 44956 54260 45008
rect 51264 44820 51316 44872
rect 54116 44888 54168 44940
rect 54300 44888 54352 44940
rect 55588 44931 55640 44940
rect 55588 44897 55597 44931
rect 55597 44897 55631 44931
rect 55631 44897 55640 44931
rect 55588 44888 55640 44897
rect 56048 44888 56100 44940
rect 57980 44931 58032 44940
rect 57980 44897 57989 44931
rect 57989 44897 58023 44931
rect 58023 44897 58032 44931
rect 57980 44888 58032 44897
rect 53932 44820 53984 44872
rect 56692 44863 56744 44872
rect 56692 44829 56701 44863
rect 56701 44829 56735 44863
rect 56735 44829 56744 44863
rect 56692 44820 56744 44829
rect 54392 44752 54444 44804
rect 58164 44795 58216 44804
rect 58164 44761 58173 44795
rect 58173 44761 58207 44795
rect 58207 44761 58216 44795
rect 58164 44752 58216 44761
rect 54944 44727 54996 44736
rect 54944 44693 54953 44727
rect 54953 44693 54987 44727
rect 54987 44693 54996 44727
rect 54944 44684 54996 44693
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 51080 44480 51132 44532
rect 51264 44480 51316 44532
rect 52092 44480 52144 44532
rect 56692 44480 56744 44532
rect 57980 44523 58032 44532
rect 57980 44489 57989 44523
rect 57989 44489 58023 44523
rect 58023 44489 58032 44523
rect 57980 44480 58032 44489
rect 55588 44412 55640 44464
rect 1400 44319 1452 44328
rect 1400 44285 1409 44319
rect 1409 44285 1443 44319
rect 1443 44285 1452 44319
rect 1400 44276 1452 44285
rect 50712 44276 50764 44328
rect 52552 44344 52604 44396
rect 56508 44344 56560 44396
rect 57704 44387 57756 44396
rect 57704 44353 57713 44387
rect 57713 44353 57747 44387
rect 57747 44353 57756 44387
rect 57704 44344 57756 44353
rect 50620 44208 50672 44260
rect 52460 44276 52512 44328
rect 52920 44319 52972 44328
rect 52920 44285 52929 44319
rect 52929 44285 52963 44319
rect 52963 44285 52972 44319
rect 52920 44276 52972 44285
rect 54392 44276 54444 44328
rect 54484 44319 54536 44328
rect 54484 44285 54493 44319
rect 54493 44285 54527 44319
rect 54527 44285 54536 44319
rect 54484 44276 54536 44285
rect 55128 44208 55180 44260
rect 56876 44251 56928 44260
rect 56876 44217 56885 44251
rect 56885 44217 56919 44251
rect 56919 44217 56928 44251
rect 56876 44208 56928 44217
rect 57060 44251 57112 44260
rect 57060 44217 57069 44251
rect 57069 44217 57103 44251
rect 57103 44217 57112 44251
rect 57060 44208 57112 44217
rect 51448 44140 51500 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 50620 43936 50672 43988
rect 51540 43979 51592 43988
rect 51540 43945 51549 43979
rect 51549 43945 51583 43979
rect 51583 43945 51592 43979
rect 51540 43936 51592 43945
rect 52552 43979 52604 43988
rect 52552 43945 52561 43979
rect 52561 43945 52595 43979
rect 52595 43945 52604 43979
rect 52552 43936 52604 43945
rect 55128 43979 55180 43988
rect 55128 43945 55137 43979
rect 55137 43945 55171 43979
rect 55171 43945 55180 43979
rect 55128 43936 55180 43945
rect 56876 43936 56928 43988
rect 58072 43936 58124 43988
rect 50712 43868 50764 43920
rect 52644 43911 52696 43920
rect 51172 43800 51224 43852
rect 51448 43843 51500 43852
rect 51448 43809 51457 43843
rect 51457 43809 51491 43843
rect 51491 43809 51500 43843
rect 51448 43800 51500 43809
rect 52644 43877 52653 43911
rect 52653 43877 52687 43911
rect 52687 43877 52696 43911
rect 52644 43868 52696 43877
rect 54944 43868 54996 43920
rect 52736 43843 52788 43852
rect 52736 43809 52745 43843
rect 52745 43809 52779 43843
rect 52779 43809 52788 43843
rect 52736 43800 52788 43809
rect 53196 43800 53248 43852
rect 54116 43843 54168 43852
rect 54116 43809 54125 43843
rect 54125 43809 54159 43843
rect 54159 43809 54168 43843
rect 54116 43800 54168 43809
rect 54300 43843 54352 43852
rect 54300 43809 54309 43843
rect 54309 43809 54343 43843
rect 54343 43809 54352 43843
rect 54300 43800 54352 43809
rect 54392 43843 54444 43852
rect 54392 43809 54401 43843
rect 54401 43809 54435 43843
rect 54435 43809 54444 43843
rect 54392 43800 54444 43809
rect 53932 43639 53984 43648
rect 53932 43605 53941 43639
rect 53941 43605 53975 43639
rect 53975 43605 53984 43639
rect 53932 43596 53984 43605
rect 54208 43707 54260 43716
rect 54208 43673 54217 43707
rect 54217 43673 54251 43707
rect 54251 43673 54260 43707
rect 54852 43732 54904 43784
rect 55404 43800 55456 43852
rect 57612 43800 57664 43852
rect 54208 43664 54260 43673
rect 55680 43664 55732 43716
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 52644 43392 52696 43444
rect 52736 43324 52788 43376
rect 51172 43256 51224 43308
rect 1400 43231 1452 43240
rect 1400 43197 1409 43231
rect 1409 43197 1443 43231
rect 1443 43197 1452 43231
rect 1400 43188 1452 43197
rect 50620 43188 50672 43240
rect 52644 43256 52696 43308
rect 54208 43324 54260 43376
rect 55036 43324 55088 43376
rect 54116 43256 54168 43308
rect 54944 43256 54996 43308
rect 51632 43188 51684 43240
rect 52092 43231 52144 43240
rect 52092 43197 52101 43231
rect 52101 43197 52135 43231
rect 52135 43197 52144 43231
rect 52092 43188 52144 43197
rect 51540 43120 51592 43172
rect 53840 43188 53892 43240
rect 54208 43231 54260 43240
rect 54208 43197 54217 43231
rect 54217 43197 54251 43231
rect 54251 43197 54260 43231
rect 54208 43188 54260 43197
rect 52920 43120 52972 43172
rect 54024 43120 54076 43172
rect 54484 43120 54536 43172
rect 55128 43188 55180 43240
rect 55864 43120 55916 43172
rect 57980 43163 58032 43172
rect 57980 43129 57989 43163
rect 57989 43129 58023 43163
rect 58023 43129 58032 43163
rect 57980 43120 58032 43129
rect 58164 43163 58216 43172
rect 58164 43129 58173 43163
rect 58173 43129 58207 43163
rect 58207 43129 58216 43163
rect 58164 43120 58216 43129
rect 51172 43095 51224 43104
rect 51172 43061 51181 43095
rect 51181 43061 51215 43095
rect 51215 43061 51224 43095
rect 51172 43052 51224 43061
rect 51448 43052 51500 43104
rect 56416 43095 56468 43104
rect 56416 43061 56425 43095
rect 56425 43061 56459 43095
rect 56459 43061 56468 43095
rect 56416 43052 56468 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 50620 42848 50672 42900
rect 51632 42891 51684 42900
rect 51632 42857 51641 42891
rect 51641 42857 51675 42891
rect 51675 42857 51684 42891
rect 51632 42848 51684 42857
rect 52092 42848 52144 42900
rect 50528 42780 50580 42832
rect 51172 42780 51224 42832
rect 52828 42780 52880 42832
rect 1400 42755 1452 42764
rect 1400 42721 1409 42755
rect 1409 42721 1443 42755
rect 1443 42721 1452 42755
rect 1400 42712 1452 42721
rect 50988 42712 51040 42764
rect 51540 42712 51592 42764
rect 52920 42755 52972 42764
rect 52920 42721 52929 42755
rect 52929 42721 52963 42755
rect 52963 42721 52972 42755
rect 52920 42712 52972 42721
rect 54208 42780 54260 42832
rect 52736 42576 52788 42628
rect 53932 42712 53984 42764
rect 56416 42780 56468 42832
rect 53840 42687 53892 42696
rect 53840 42653 53849 42687
rect 53849 42653 53883 42687
rect 53883 42653 53892 42687
rect 53840 42644 53892 42653
rect 55036 42755 55088 42764
rect 55036 42721 55045 42755
rect 55045 42721 55079 42755
rect 55079 42721 55088 42755
rect 55036 42712 55088 42721
rect 55404 42644 55456 42696
rect 57152 42712 57204 42764
rect 57980 42848 58032 42900
rect 57704 42687 57756 42696
rect 57704 42653 57713 42687
rect 57713 42653 57747 42687
rect 57747 42653 57756 42687
rect 57704 42644 57756 42653
rect 55036 42576 55088 42628
rect 51080 42508 51132 42560
rect 51172 42508 51224 42560
rect 51632 42508 51684 42560
rect 54116 42508 54168 42560
rect 55128 42508 55180 42560
rect 56968 42551 57020 42560
rect 56968 42517 56977 42551
rect 56977 42517 57011 42551
rect 57011 42517 57020 42551
rect 56968 42508 57020 42517
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 50988 42347 51040 42356
rect 50988 42313 50997 42347
rect 50997 42313 51031 42347
rect 51031 42313 51040 42347
rect 50988 42304 51040 42313
rect 54208 42304 54260 42356
rect 55404 42347 55456 42356
rect 55404 42313 55413 42347
rect 55413 42313 55447 42347
rect 55447 42313 55456 42347
rect 55404 42304 55456 42313
rect 55864 42347 55916 42356
rect 55864 42313 55873 42347
rect 55873 42313 55907 42347
rect 55907 42313 55916 42347
rect 55864 42304 55916 42313
rect 57152 42347 57204 42356
rect 57152 42313 57161 42347
rect 57161 42313 57195 42347
rect 57195 42313 57204 42347
rect 57152 42304 57204 42313
rect 50436 42279 50488 42288
rect 50436 42245 50445 42279
rect 50445 42245 50479 42279
rect 50479 42245 50488 42279
rect 50436 42236 50488 42245
rect 52184 42279 52236 42288
rect 52184 42245 52193 42279
rect 52193 42245 52227 42279
rect 52227 42245 52236 42279
rect 52184 42236 52236 42245
rect 50528 42211 50580 42220
rect 50528 42177 50537 42211
rect 50537 42177 50571 42211
rect 50571 42177 50580 42211
rect 50528 42168 50580 42177
rect 55036 42168 55088 42220
rect 49424 42143 49476 42152
rect 49424 42109 49433 42143
rect 49433 42109 49467 42143
rect 49467 42109 49476 42143
rect 49424 42100 49476 42109
rect 50160 41964 50212 42016
rect 51172 42100 51224 42152
rect 51337 42143 51389 42152
rect 51337 42109 51362 42143
rect 51362 42109 51389 42143
rect 51337 42100 51389 42109
rect 52092 42143 52144 42152
rect 52092 42109 52101 42143
rect 52101 42109 52135 42143
rect 52135 42109 52144 42143
rect 52092 42100 52144 42109
rect 52736 42143 52788 42152
rect 52736 42109 52745 42143
rect 52745 42109 52779 42143
rect 52779 42109 52788 42143
rect 52736 42100 52788 42109
rect 52920 42143 52972 42152
rect 52920 42109 52929 42143
rect 52929 42109 52963 42143
rect 52963 42109 52972 42143
rect 52920 42100 52972 42109
rect 54024 42143 54076 42152
rect 54024 42109 54033 42143
rect 54033 42109 54067 42143
rect 54067 42109 54076 42143
rect 54024 42100 54076 42109
rect 54116 42100 54168 42152
rect 54852 42100 54904 42152
rect 56140 42100 56192 42152
rect 52828 42032 52880 42084
rect 55404 42032 55456 42084
rect 57980 42075 58032 42084
rect 57980 42041 57989 42075
rect 57989 42041 58023 42075
rect 58023 42041 58032 42075
rect 57980 42032 58032 42041
rect 58164 42075 58216 42084
rect 58164 42041 58173 42075
rect 58173 42041 58207 42075
rect 58207 42041 58216 42075
rect 58164 42032 58216 42041
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 52092 41760 52144 41812
rect 55404 41760 55456 41812
rect 57704 41760 57756 41812
rect 57980 41760 58032 41812
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 50068 41624 50120 41676
rect 51448 41667 51500 41676
rect 51448 41633 51457 41667
rect 51457 41633 51491 41667
rect 51491 41633 51500 41667
rect 51448 41624 51500 41633
rect 51632 41667 51684 41676
rect 51632 41633 51641 41667
rect 51641 41633 51675 41667
rect 51675 41633 51684 41667
rect 51632 41624 51684 41633
rect 53196 41624 53248 41676
rect 53380 41667 53432 41676
rect 53380 41633 53389 41667
rect 53389 41633 53423 41667
rect 53423 41633 53432 41667
rect 53380 41624 53432 41633
rect 53932 41624 53984 41676
rect 52460 41488 52512 41540
rect 53840 41556 53892 41608
rect 54852 41667 54904 41676
rect 54852 41633 54861 41667
rect 54861 41633 54895 41667
rect 54895 41633 54904 41667
rect 54852 41624 54904 41633
rect 54024 41488 54076 41540
rect 56140 41488 56192 41540
rect 54852 41463 54904 41472
rect 54852 41429 54861 41463
rect 54861 41429 54895 41463
rect 54895 41429 54904 41463
rect 54852 41420 54904 41429
rect 58256 41624 58308 41676
rect 57520 41599 57572 41608
rect 57520 41565 57529 41599
rect 57529 41565 57563 41599
rect 57563 41565 57572 41599
rect 57520 41556 57572 41565
rect 56416 41488 56468 41540
rect 57060 41463 57112 41472
rect 57060 41429 57069 41463
rect 57069 41429 57103 41463
rect 57103 41429 57112 41463
rect 57060 41420 57112 41429
rect 57612 41420 57664 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 51080 41012 51132 41064
rect 51448 41012 51500 41064
rect 50620 40944 50672 40996
rect 53380 41216 53432 41268
rect 53840 41216 53892 41268
rect 54116 41012 54168 41064
rect 54668 41012 54720 41064
rect 54852 41055 54904 41064
rect 54852 41021 54886 41055
rect 54886 41021 54904 41055
rect 54852 41012 54904 41021
rect 57520 41012 57572 41064
rect 57244 40987 57296 40996
rect 57244 40953 57253 40987
rect 57253 40953 57287 40987
rect 57287 40953 57296 40987
rect 57244 40944 57296 40953
rect 57428 40987 57480 40996
rect 57428 40953 57437 40987
rect 57437 40953 57471 40987
rect 57471 40953 57480 40987
rect 57428 40944 57480 40953
rect 57980 40987 58032 40996
rect 57980 40953 57989 40987
rect 57989 40953 58023 40987
rect 58023 40953 58032 40987
rect 57980 40944 58032 40953
rect 53840 40876 53892 40928
rect 54024 40876 54076 40928
rect 57888 40876 57940 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 1400 40579 1452 40588
rect 1400 40545 1409 40579
rect 1409 40545 1443 40579
rect 1443 40545 1452 40579
rect 1400 40536 1452 40545
rect 50620 40604 50672 40656
rect 51908 40647 51960 40656
rect 51908 40613 51917 40647
rect 51917 40613 51951 40647
rect 51951 40613 51960 40647
rect 51908 40604 51960 40613
rect 56416 40672 56468 40724
rect 57980 40672 58032 40724
rect 55220 40604 55272 40656
rect 50620 40468 50672 40520
rect 51816 40468 51868 40520
rect 52460 40536 52512 40588
rect 53472 40579 53524 40588
rect 53472 40545 53481 40579
rect 53481 40545 53515 40579
rect 53515 40545 53524 40579
rect 53472 40536 53524 40545
rect 53840 40579 53892 40588
rect 53840 40545 53849 40579
rect 53849 40545 53883 40579
rect 53883 40545 53892 40579
rect 53840 40536 53892 40545
rect 55128 40579 55180 40588
rect 53564 40511 53616 40520
rect 53564 40477 53573 40511
rect 53573 40477 53607 40511
rect 53607 40477 53616 40511
rect 53564 40468 53616 40477
rect 53932 40468 53984 40520
rect 54300 40468 54352 40520
rect 55128 40545 55137 40579
rect 55137 40545 55171 40579
rect 55171 40545 55180 40579
rect 55128 40536 55180 40545
rect 55496 40536 55548 40588
rect 56600 40536 56652 40588
rect 57060 40468 57112 40520
rect 57152 40468 57204 40520
rect 57612 40468 57664 40520
rect 54024 40400 54076 40452
rect 55036 40400 55088 40452
rect 55588 40400 55640 40452
rect 53104 40375 53156 40384
rect 53104 40341 53113 40375
rect 53113 40341 53147 40375
rect 53147 40341 53156 40375
rect 53104 40332 53156 40341
rect 55404 40332 55456 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 51908 40128 51960 40180
rect 54024 40103 54076 40112
rect 54024 40069 54033 40103
rect 54033 40069 54067 40103
rect 54067 40069 54076 40103
rect 54024 40060 54076 40069
rect 1400 39967 1452 39976
rect 1400 39933 1409 39967
rect 1409 39933 1443 39967
rect 1443 39933 1452 39967
rect 1400 39924 1452 39933
rect 50068 39924 50120 39976
rect 51172 39924 51224 39976
rect 51540 39967 51592 39976
rect 51540 39933 51549 39967
rect 51549 39933 51583 39967
rect 51583 39933 51592 39967
rect 51540 39924 51592 39933
rect 51816 39924 51868 39976
rect 52368 39967 52420 39976
rect 52368 39933 52377 39967
rect 52377 39933 52411 39967
rect 52411 39933 52420 39967
rect 52368 39924 52420 39933
rect 53748 39924 53800 39976
rect 53840 39924 53892 39976
rect 54300 39967 54352 39976
rect 54300 39933 54309 39967
rect 54309 39933 54343 39967
rect 54343 39933 54352 39967
rect 54484 39967 54536 39976
rect 54300 39924 54352 39933
rect 54484 39933 54493 39967
rect 54493 39933 54527 39967
rect 54527 39933 54536 39967
rect 54484 39924 54536 39933
rect 54852 39992 54904 40044
rect 57244 40128 57296 40180
rect 55036 39924 55088 39976
rect 55404 39924 55456 39976
rect 50712 39856 50764 39908
rect 53564 39788 53616 39840
rect 53748 39788 53800 39840
rect 54484 39788 54536 39840
rect 55496 39788 55548 39840
rect 56600 39788 56652 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 52368 39584 52420 39636
rect 53012 39584 53064 39636
rect 53840 39584 53892 39636
rect 54852 39584 54904 39636
rect 55496 39584 55548 39636
rect 51540 39516 51592 39568
rect 52552 39491 52604 39500
rect 52552 39457 52561 39491
rect 52561 39457 52595 39491
rect 52595 39457 52604 39491
rect 52552 39448 52604 39457
rect 52368 39380 52420 39432
rect 52736 39491 52788 39500
rect 52736 39457 52745 39491
rect 52745 39457 52779 39491
rect 52779 39457 52788 39491
rect 52736 39448 52788 39457
rect 53012 39448 53064 39500
rect 55864 39516 55916 39568
rect 51908 39312 51960 39364
rect 53748 39423 53800 39432
rect 53748 39389 53757 39423
rect 53757 39389 53791 39423
rect 53791 39389 53800 39423
rect 53748 39380 53800 39389
rect 55036 39312 55088 39364
rect 56692 39380 56744 39432
rect 57520 39380 57572 39432
rect 56968 39355 57020 39364
rect 56968 39321 56977 39355
rect 56977 39321 57011 39355
rect 57011 39321 57020 39355
rect 56968 39312 57020 39321
rect 57152 39244 57204 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 51172 39040 51224 39092
rect 52368 39040 52420 39092
rect 52644 39040 52696 39092
rect 55588 39040 55640 39092
rect 1400 38879 1452 38888
rect 1400 38845 1409 38879
rect 1409 38845 1443 38879
rect 1443 38845 1452 38879
rect 1400 38836 1452 38845
rect 55220 38972 55272 39024
rect 50712 38904 50764 38956
rect 52552 38904 52604 38956
rect 52644 38904 52696 38956
rect 53196 38904 53248 38956
rect 53288 38904 53340 38956
rect 51172 38836 51224 38888
rect 51908 38879 51960 38888
rect 51908 38845 51917 38879
rect 51917 38845 51951 38879
rect 51951 38845 51960 38879
rect 51908 38836 51960 38845
rect 52460 38836 52512 38888
rect 53012 38879 53064 38888
rect 53012 38845 53021 38879
rect 53021 38845 53055 38879
rect 53055 38845 53064 38879
rect 53012 38836 53064 38845
rect 53564 38836 53616 38888
rect 55036 38879 55088 38888
rect 55036 38845 55045 38879
rect 55045 38845 55079 38879
rect 55079 38845 55088 38879
rect 55036 38836 55088 38845
rect 55496 38836 55548 38888
rect 56232 38836 56284 38888
rect 52000 38700 52052 38752
rect 53196 38700 53248 38752
rect 54116 38743 54168 38752
rect 54116 38709 54125 38743
rect 54125 38709 54159 38743
rect 54159 38709 54168 38743
rect 54116 38700 54168 38709
rect 56600 38768 56652 38820
rect 57704 38768 57756 38820
rect 57520 38700 57572 38752
rect 57888 38700 57940 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 50712 38496 50764 38548
rect 52828 38496 52880 38548
rect 49700 38360 49752 38412
rect 52552 38428 52604 38480
rect 52000 38403 52052 38412
rect 52000 38369 52009 38403
rect 52009 38369 52043 38403
rect 52043 38369 52052 38403
rect 52000 38360 52052 38369
rect 52644 38360 52696 38412
rect 54116 38496 54168 38548
rect 54208 38496 54260 38548
rect 56692 38496 56744 38548
rect 57612 38496 57664 38548
rect 53196 38428 53248 38480
rect 54024 38360 54076 38412
rect 54760 38360 54812 38412
rect 53104 38292 53156 38344
rect 53380 38335 53432 38344
rect 53380 38301 53389 38335
rect 53389 38301 53423 38335
rect 53423 38301 53432 38335
rect 53380 38292 53432 38301
rect 57060 38360 57112 38412
rect 57980 38403 58032 38412
rect 57980 38369 57989 38403
rect 57989 38369 58023 38403
rect 58023 38369 58032 38403
rect 57980 38360 58032 38369
rect 58164 38403 58216 38412
rect 58164 38369 58173 38403
rect 58173 38369 58207 38403
rect 58207 38369 58216 38403
rect 58164 38360 58216 38369
rect 55588 38292 55640 38344
rect 50068 38156 50120 38208
rect 56968 38224 57020 38276
rect 55588 38156 55640 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 53012 37995 53064 38004
rect 53012 37961 53021 37995
rect 53021 37961 53055 37995
rect 53055 37961 53064 37995
rect 53012 37952 53064 37961
rect 53472 37952 53524 38004
rect 57980 37995 58032 38004
rect 56968 37927 57020 37936
rect 56968 37893 56977 37927
rect 56977 37893 57011 37927
rect 57011 37893 57020 37927
rect 56968 37884 57020 37893
rect 54024 37859 54076 37868
rect 54024 37825 54033 37859
rect 54033 37825 54067 37859
rect 54067 37825 54076 37859
rect 54024 37816 54076 37825
rect 1400 37791 1452 37800
rect 1400 37757 1409 37791
rect 1409 37757 1443 37791
rect 1443 37757 1452 37791
rect 1400 37748 1452 37757
rect 50068 37791 50120 37800
rect 50068 37757 50077 37791
rect 50077 37757 50111 37791
rect 50111 37757 50120 37791
rect 50068 37748 50120 37757
rect 50620 37748 50672 37800
rect 51356 37748 51408 37800
rect 53472 37748 53524 37800
rect 54760 37816 54812 37868
rect 57980 37961 57989 37995
rect 57989 37961 58023 37995
rect 58023 37961 58032 37995
rect 57980 37952 58032 37961
rect 54668 37748 54720 37800
rect 54852 37748 54904 37800
rect 49056 37612 49108 37664
rect 54944 37680 54996 37732
rect 55496 37680 55548 37732
rect 55220 37612 55272 37664
rect 57612 37748 57664 37800
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 54944 37451 54996 37460
rect 49056 37315 49108 37324
rect 49056 37281 49065 37315
rect 49065 37281 49099 37315
rect 49099 37281 49108 37315
rect 49056 37272 49108 37281
rect 49700 37315 49752 37324
rect 49700 37281 49709 37315
rect 49709 37281 49743 37315
rect 49743 37281 49752 37315
rect 49700 37272 49752 37281
rect 49792 37247 49844 37256
rect 49792 37213 49801 37247
rect 49801 37213 49835 37247
rect 49835 37213 49844 37247
rect 49792 37204 49844 37213
rect 51172 37272 51224 37324
rect 51908 37315 51960 37324
rect 51908 37281 51917 37315
rect 51917 37281 51951 37315
rect 51951 37281 51960 37315
rect 51908 37272 51960 37281
rect 52092 37315 52144 37324
rect 52092 37281 52101 37315
rect 52101 37281 52135 37315
rect 52135 37281 52144 37315
rect 52092 37272 52144 37281
rect 52460 37272 52512 37324
rect 54668 37383 54720 37392
rect 54668 37349 54677 37383
rect 54677 37349 54711 37383
rect 54711 37349 54720 37383
rect 54668 37340 54720 37349
rect 54944 37417 54953 37451
rect 54953 37417 54987 37451
rect 54987 37417 54996 37451
rect 54944 37408 54996 37417
rect 55496 37451 55548 37460
rect 55496 37417 55505 37451
rect 55505 37417 55539 37451
rect 55539 37417 55548 37451
rect 55496 37408 55548 37417
rect 57704 37451 57756 37460
rect 57704 37417 57713 37451
rect 57713 37417 57747 37451
rect 57747 37417 57756 37451
rect 57704 37408 57756 37417
rect 54576 37315 54628 37324
rect 52368 37204 52420 37256
rect 52000 37179 52052 37188
rect 52000 37145 52009 37179
rect 52009 37145 52043 37179
rect 52043 37145 52052 37179
rect 52000 37136 52052 37145
rect 51356 37068 51408 37120
rect 53840 37204 53892 37256
rect 54576 37281 54585 37315
rect 54585 37281 54619 37315
rect 54619 37281 54628 37315
rect 54576 37272 54628 37281
rect 54760 37315 54812 37324
rect 54760 37281 54769 37315
rect 54769 37281 54803 37315
rect 54803 37281 54812 37315
rect 54760 37272 54812 37281
rect 55128 37272 55180 37324
rect 55588 37315 55640 37324
rect 55588 37281 55597 37315
rect 55597 37281 55631 37315
rect 55631 37281 55640 37315
rect 55588 37272 55640 37281
rect 57060 37247 57112 37256
rect 57060 37213 57069 37247
rect 57069 37213 57103 37247
rect 57103 37213 57112 37247
rect 57060 37204 57112 37213
rect 54024 37068 54076 37120
rect 54576 37068 54628 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 52460 36864 52512 36916
rect 53840 36864 53892 36916
rect 52092 36796 52144 36848
rect 53748 36796 53800 36848
rect 1400 36703 1452 36712
rect 1400 36669 1409 36703
rect 1409 36669 1443 36703
rect 1443 36669 1452 36703
rect 1400 36660 1452 36669
rect 50160 36660 50212 36712
rect 51356 36592 51408 36644
rect 52736 36703 52788 36712
rect 52736 36669 52750 36703
rect 52750 36669 52784 36703
rect 52784 36669 52788 36703
rect 52736 36660 52788 36669
rect 53012 36660 53064 36712
rect 54024 36703 54076 36712
rect 54024 36669 54033 36703
rect 54033 36669 54067 36703
rect 54067 36669 54076 36703
rect 54024 36660 54076 36669
rect 54300 36660 54352 36712
rect 54852 36660 54904 36712
rect 57612 36864 57664 36916
rect 58164 36771 58216 36780
rect 58164 36737 58173 36771
rect 58173 36737 58207 36771
rect 58207 36737 58216 36771
rect 58164 36728 58216 36737
rect 57428 36703 57480 36712
rect 57428 36669 57437 36703
rect 57437 36669 57471 36703
rect 57471 36669 57480 36703
rect 57428 36660 57480 36669
rect 54668 36592 54720 36644
rect 57980 36635 58032 36644
rect 57980 36601 57989 36635
rect 57989 36601 58023 36635
rect 58023 36601 58032 36635
rect 57980 36592 58032 36601
rect 51080 36524 51132 36576
rect 52644 36524 52696 36576
rect 54116 36567 54168 36576
rect 54116 36533 54125 36567
rect 54125 36533 54159 36567
rect 54159 36533 54168 36567
rect 54116 36524 54168 36533
rect 54852 36524 54904 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 52552 36320 52604 36372
rect 52644 36320 52696 36372
rect 54668 36363 54720 36372
rect 54668 36329 54677 36363
rect 54677 36329 54711 36363
rect 54711 36329 54720 36363
rect 54668 36320 54720 36329
rect 56968 36363 57020 36372
rect 56968 36329 56977 36363
rect 56977 36329 57011 36363
rect 57011 36329 57020 36363
rect 56968 36320 57020 36329
rect 57980 36320 58032 36372
rect 52000 36252 52052 36304
rect 1400 36227 1452 36236
rect 1400 36193 1409 36227
rect 1409 36193 1443 36227
rect 1443 36193 1452 36227
rect 1400 36184 1452 36193
rect 51264 36184 51316 36236
rect 53012 36252 53064 36304
rect 54024 36252 54076 36304
rect 53840 36227 53892 36236
rect 53840 36193 53849 36227
rect 53849 36193 53883 36227
rect 53883 36193 53892 36227
rect 54116 36227 54168 36236
rect 53840 36184 53892 36193
rect 54116 36193 54125 36227
rect 54125 36193 54159 36227
rect 54159 36193 54168 36227
rect 54116 36184 54168 36193
rect 55404 36252 55456 36304
rect 55588 36227 55640 36236
rect 52368 36116 52420 36168
rect 52828 36159 52880 36168
rect 52828 36125 52837 36159
rect 52837 36125 52871 36159
rect 52871 36125 52880 36159
rect 52828 36116 52880 36125
rect 55588 36193 55597 36227
rect 55597 36193 55631 36227
rect 55631 36193 55640 36227
rect 55588 36184 55640 36193
rect 56876 36227 56928 36236
rect 56876 36193 56885 36227
rect 56885 36193 56919 36227
rect 56919 36193 56928 36227
rect 56876 36184 56928 36193
rect 56968 36184 57020 36236
rect 52736 35980 52788 36032
rect 52828 35980 52880 36032
rect 54852 35980 54904 36032
rect 54944 35980 54996 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 55220 35776 55272 35828
rect 56876 35776 56928 35828
rect 51172 35640 51224 35692
rect 50896 35572 50948 35624
rect 51724 35615 51776 35624
rect 51724 35581 51733 35615
rect 51733 35581 51767 35615
rect 51767 35581 51776 35615
rect 51724 35572 51776 35581
rect 50620 35504 50672 35556
rect 52092 35572 52144 35624
rect 56968 35640 57020 35692
rect 51264 35436 51316 35488
rect 51816 35479 51868 35488
rect 51816 35445 51825 35479
rect 51825 35445 51859 35479
rect 51859 35445 51868 35479
rect 51816 35436 51868 35445
rect 53104 35615 53156 35624
rect 53104 35581 53113 35615
rect 53113 35581 53147 35615
rect 53147 35581 53156 35615
rect 53104 35572 53156 35581
rect 53932 35572 53984 35624
rect 58072 35572 58124 35624
rect 58348 35572 58400 35624
rect 53012 35504 53064 35556
rect 55404 35547 55456 35556
rect 55404 35513 55413 35547
rect 55413 35513 55447 35547
rect 55447 35513 55456 35547
rect 55404 35504 55456 35513
rect 56232 35547 56284 35556
rect 56232 35513 56241 35547
rect 56241 35513 56275 35547
rect 56275 35513 56284 35547
rect 56232 35504 56284 35513
rect 56692 35504 56744 35556
rect 53104 35436 53156 35488
rect 54392 35436 54444 35488
rect 55128 35436 55180 35488
rect 56324 35479 56376 35488
rect 56324 35445 56333 35479
rect 56333 35445 56367 35479
rect 56367 35445 56376 35479
rect 56324 35436 56376 35445
rect 56600 35436 56652 35488
rect 57428 35436 57480 35488
rect 57888 35436 57940 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 53932 35232 53984 35284
rect 56968 35275 57020 35284
rect 56968 35241 56977 35275
rect 56977 35241 57011 35275
rect 57011 35241 57020 35275
rect 56968 35232 57020 35241
rect 51816 35164 51868 35216
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 49700 35139 49752 35148
rect 49700 35105 49709 35139
rect 49709 35105 49743 35139
rect 49743 35105 49752 35139
rect 49700 35096 49752 35105
rect 49884 35139 49936 35148
rect 49884 35105 49893 35139
rect 49893 35105 49927 35139
rect 49927 35105 49936 35139
rect 49884 35096 49936 35105
rect 51172 35096 51224 35148
rect 56324 35164 56376 35216
rect 50068 35028 50120 35080
rect 50344 35003 50396 35012
rect 50344 34969 50353 35003
rect 50353 34969 50387 35003
rect 50387 34969 50396 35003
rect 50344 34960 50396 34969
rect 51448 34960 51500 35012
rect 53196 35003 53248 35012
rect 53196 34969 53205 35003
rect 53205 34969 53239 35003
rect 53239 34969 53248 35003
rect 54392 35096 54444 35148
rect 55036 35096 55088 35148
rect 53840 35028 53892 35080
rect 54300 35071 54352 35080
rect 54300 35037 54309 35071
rect 54309 35037 54343 35071
rect 54343 35037 54352 35071
rect 54300 35028 54352 35037
rect 58256 35028 58308 35080
rect 53196 34960 53248 34969
rect 50160 34892 50212 34944
rect 53012 34892 53064 34944
rect 54208 34892 54260 34944
rect 54300 34892 54352 34944
rect 55588 34892 55640 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 50160 34688 50212 34740
rect 50896 34688 50948 34740
rect 51724 34688 51776 34740
rect 52092 34688 52144 34740
rect 54300 34688 54352 34740
rect 55036 34731 55088 34740
rect 55036 34697 55045 34731
rect 55045 34697 55079 34731
rect 55079 34697 55088 34731
rect 55036 34688 55088 34697
rect 55128 34688 55180 34740
rect 50988 34484 51040 34536
rect 51908 34527 51960 34536
rect 51908 34493 51917 34527
rect 51917 34493 51951 34527
rect 51951 34493 51960 34527
rect 51908 34484 51960 34493
rect 53564 34484 53616 34536
rect 54208 34527 54260 34536
rect 54208 34493 54217 34527
rect 54217 34493 54251 34527
rect 54251 34493 54260 34527
rect 54208 34484 54260 34493
rect 54944 34620 54996 34672
rect 56416 34663 56468 34672
rect 56416 34629 56425 34663
rect 56425 34629 56459 34663
rect 56459 34629 56468 34663
rect 56416 34620 56468 34629
rect 54668 34552 54720 34604
rect 54852 34552 54904 34604
rect 57060 34595 57112 34604
rect 54576 34527 54628 34536
rect 54576 34493 54585 34527
rect 54585 34493 54619 34527
rect 54619 34493 54628 34527
rect 54576 34484 54628 34493
rect 57060 34561 57069 34595
rect 57069 34561 57103 34595
rect 57103 34561 57112 34595
rect 57060 34552 57112 34561
rect 56876 34527 56928 34536
rect 50804 34416 50856 34468
rect 51080 34459 51132 34468
rect 51080 34425 51089 34459
rect 51089 34425 51123 34459
rect 51123 34425 51132 34459
rect 51080 34416 51132 34425
rect 52368 34416 52420 34468
rect 54852 34416 54904 34468
rect 56876 34493 56885 34527
rect 56885 34493 56919 34527
rect 56919 34493 56928 34527
rect 56876 34484 56928 34493
rect 55404 34416 55456 34468
rect 55956 34416 56008 34468
rect 57980 34527 58032 34536
rect 57980 34493 57989 34527
rect 57989 34493 58023 34527
rect 58023 34493 58032 34527
rect 57980 34484 58032 34493
rect 50712 34348 50764 34400
rect 52736 34348 52788 34400
rect 52920 34348 52972 34400
rect 57152 34348 57204 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 50620 34144 50672 34196
rect 51908 34187 51960 34196
rect 51908 34153 51917 34187
rect 51917 34153 51951 34187
rect 51951 34153 51960 34187
rect 51908 34144 51960 34153
rect 52736 34144 52788 34196
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 55220 34076 55272 34128
rect 50068 34008 50120 34060
rect 52184 34008 52236 34060
rect 52460 33940 52512 33992
rect 53380 34051 53432 34060
rect 53380 34017 53389 34051
rect 53389 34017 53423 34051
rect 53423 34017 53432 34051
rect 53380 34008 53432 34017
rect 56048 34008 56100 34060
rect 56692 34144 56744 34196
rect 56784 34119 56836 34128
rect 56784 34085 56793 34119
rect 56793 34085 56827 34119
rect 56827 34085 56836 34119
rect 56784 34076 56836 34085
rect 53012 33872 53064 33924
rect 53288 33847 53340 33856
rect 53288 33813 53297 33847
rect 53297 33813 53331 33847
rect 53331 33813 53340 33847
rect 53288 33804 53340 33813
rect 53840 33940 53892 33992
rect 57612 33940 57664 33992
rect 57980 33940 58032 33992
rect 55404 33872 55456 33924
rect 55128 33804 55180 33856
rect 57980 33847 58032 33856
rect 57980 33813 57989 33847
rect 57989 33813 58023 33847
rect 58023 33813 58032 33847
rect 57980 33804 58032 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 50712 33600 50764 33652
rect 52460 33600 52512 33652
rect 52920 33532 52972 33584
rect 54392 33532 54444 33584
rect 55588 33600 55640 33652
rect 56048 33643 56100 33652
rect 56048 33609 56057 33643
rect 56057 33609 56091 33643
rect 56091 33609 56100 33643
rect 56048 33600 56100 33609
rect 58164 33575 58216 33584
rect 50896 33464 50948 33516
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 50068 33396 50120 33448
rect 50712 33396 50764 33448
rect 53380 33464 53432 33516
rect 52552 33439 52604 33448
rect 52552 33405 52561 33439
rect 52561 33405 52595 33439
rect 52595 33405 52604 33439
rect 52552 33396 52604 33405
rect 52828 33439 52880 33448
rect 52828 33405 52837 33439
rect 52837 33405 52871 33439
rect 52871 33405 52880 33439
rect 52828 33396 52880 33405
rect 53288 33396 53340 33448
rect 53472 33396 53524 33448
rect 54392 33396 54444 33448
rect 54760 33464 54812 33516
rect 54668 33396 54720 33448
rect 55496 33396 55548 33448
rect 56048 33439 56100 33448
rect 56048 33405 56057 33439
rect 56057 33405 56091 33439
rect 56091 33405 56100 33439
rect 56048 33396 56100 33405
rect 58164 33541 58173 33575
rect 58173 33541 58207 33575
rect 58207 33541 58216 33575
rect 58164 33532 58216 33541
rect 57980 33439 58032 33448
rect 57980 33405 57989 33439
rect 57989 33405 58023 33439
rect 58023 33405 58032 33439
rect 57980 33396 58032 33405
rect 51356 33260 51408 33312
rect 52276 33260 52328 33312
rect 57520 33328 57572 33380
rect 53196 33260 53248 33312
rect 55036 33303 55088 33312
rect 55036 33269 55045 33303
rect 55045 33269 55079 33303
rect 55079 33269 55088 33303
rect 55036 33260 55088 33269
rect 57336 33303 57388 33312
rect 57336 33269 57345 33303
rect 57345 33269 57379 33303
rect 57379 33269 57388 33303
rect 57336 33260 57388 33269
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 49700 32963 49752 32972
rect 49700 32929 49709 32963
rect 49709 32929 49743 32963
rect 49743 32929 49752 32963
rect 49700 32920 49752 32929
rect 52644 33056 52696 33108
rect 52828 33099 52880 33108
rect 52828 33065 52837 33099
rect 52837 33065 52871 33099
rect 52871 33065 52880 33099
rect 52828 33056 52880 33065
rect 53564 33099 53616 33108
rect 53564 33065 53573 33099
rect 53573 33065 53607 33099
rect 53607 33065 53616 33099
rect 53564 33056 53616 33065
rect 54300 33056 54352 33108
rect 55128 33056 55180 33108
rect 52368 32988 52420 33040
rect 54116 32988 54168 33040
rect 51540 32920 51592 32972
rect 53656 32963 53708 32972
rect 53656 32929 53665 32963
rect 53665 32929 53699 32963
rect 53699 32929 53708 32963
rect 53656 32920 53708 32929
rect 54300 32963 54352 32972
rect 54300 32929 54309 32963
rect 54309 32929 54343 32963
rect 54343 32929 54352 32963
rect 54300 32920 54352 32929
rect 57152 32963 57204 32972
rect 49516 32784 49568 32836
rect 57152 32929 57161 32963
rect 57161 32929 57195 32963
rect 57195 32929 57204 32963
rect 57152 32920 57204 32929
rect 57336 32895 57388 32904
rect 52552 32784 52604 32836
rect 54024 32784 54076 32836
rect 54484 32784 54536 32836
rect 54760 32784 54812 32836
rect 57336 32861 57345 32895
rect 57345 32861 57379 32895
rect 57379 32861 57388 32895
rect 57336 32852 57388 32861
rect 55496 32784 55548 32836
rect 57520 32827 57572 32836
rect 57520 32793 57529 32827
rect 57529 32793 57563 32827
rect 57563 32793 57572 32827
rect 57520 32784 57572 32793
rect 52736 32716 52788 32768
rect 54300 32716 54352 32768
rect 54852 32716 54904 32768
rect 56600 32716 56652 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 51540 32555 51592 32564
rect 51540 32521 51549 32555
rect 51549 32521 51583 32555
rect 51583 32521 51592 32555
rect 51540 32512 51592 32521
rect 52736 32512 52788 32564
rect 52184 32444 52236 32496
rect 54944 32444 54996 32496
rect 56600 32444 56652 32496
rect 1400 32351 1452 32360
rect 1400 32317 1409 32351
rect 1409 32317 1443 32351
rect 1443 32317 1452 32351
rect 1400 32308 1452 32317
rect 53012 32376 53064 32428
rect 53656 32376 53708 32428
rect 53748 32376 53800 32428
rect 54300 32419 54352 32428
rect 54300 32385 54309 32419
rect 54309 32385 54343 32419
rect 54343 32385 54352 32419
rect 54300 32376 54352 32385
rect 55036 32376 55088 32428
rect 51724 32240 51776 32292
rect 52000 32351 52052 32360
rect 52000 32317 52009 32351
rect 52009 32317 52043 32351
rect 52043 32317 52052 32351
rect 52184 32351 52236 32360
rect 52000 32308 52052 32317
rect 52184 32317 52193 32351
rect 52193 32317 52227 32351
rect 52227 32317 52236 32351
rect 52184 32308 52236 32317
rect 53288 32308 53340 32360
rect 52276 32240 52328 32292
rect 55956 32308 56008 32360
rect 55404 32240 55456 32292
rect 50712 32172 50764 32224
rect 54116 32172 54168 32224
rect 54300 32172 54352 32224
rect 57980 32172 58032 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 51724 32011 51776 32020
rect 51724 31977 51733 32011
rect 51733 31977 51767 32011
rect 51767 31977 51776 32011
rect 51724 31968 51776 31977
rect 54484 31968 54536 32020
rect 48320 31832 48372 31884
rect 54300 31900 54352 31952
rect 55128 31943 55180 31952
rect 55128 31909 55137 31943
rect 55137 31909 55171 31943
rect 55171 31909 55180 31943
rect 57980 31943 58032 31952
rect 55128 31900 55180 31909
rect 57980 31909 57989 31943
rect 57989 31909 58023 31943
rect 58023 31909 58032 31943
rect 57980 31900 58032 31909
rect 58164 31943 58216 31952
rect 58164 31909 58173 31943
rect 58173 31909 58207 31943
rect 58207 31909 58216 31943
rect 58164 31900 58216 31909
rect 51816 31832 51868 31884
rect 52368 31832 52420 31884
rect 52460 31832 52512 31884
rect 54576 31832 54628 31884
rect 54944 31832 54996 31884
rect 58072 31832 58124 31884
rect 51908 31807 51960 31816
rect 51908 31773 51917 31807
rect 51917 31773 51951 31807
rect 51951 31773 51960 31807
rect 51908 31764 51960 31773
rect 52552 31696 52604 31748
rect 52184 31628 52236 31680
rect 52460 31628 52512 31680
rect 52736 31807 52788 31816
rect 52736 31773 52745 31807
rect 52745 31773 52779 31807
rect 52779 31773 52788 31807
rect 57428 31807 57480 31816
rect 52736 31764 52788 31773
rect 57428 31773 57437 31807
rect 57437 31773 57471 31807
rect 57471 31773 57480 31807
rect 57428 31764 57480 31773
rect 54576 31696 54628 31748
rect 56416 31696 56468 31748
rect 54392 31628 54444 31680
rect 54668 31628 54720 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 51264 31424 51316 31476
rect 51448 31424 51500 31476
rect 52736 31424 52788 31476
rect 54392 31467 54444 31476
rect 54392 31433 54401 31467
rect 54401 31433 54435 31467
rect 54435 31433 54444 31467
rect 54392 31424 54444 31433
rect 54760 31467 54812 31476
rect 54760 31433 54769 31467
rect 54769 31433 54803 31467
rect 54803 31433 54812 31467
rect 54760 31424 54812 31433
rect 51540 31356 51592 31408
rect 52000 31356 52052 31408
rect 57336 31424 57388 31476
rect 58072 31467 58124 31476
rect 58072 31433 58081 31467
rect 58081 31433 58115 31467
rect 58115 31433 58124 31467
rect 58072 31424 58124 31433
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 48872 31220 48924 31272
rect 52000 31220 52052 31272
rect 52368 31220 52420 31272
rect 51172 31152 51224 31204
rect 51540 31084 51592 31136
rect 51724 31152 51776 31204
rect 54668 31220 54720 31272
rect 54852 31263 54904 31272
rect 54852 31229 54861 31263
rect 54861 31229 54895 31263
rect 54895 31229 54904 31263
rect 54852 31220 54904 31229
rect 54944 31220 54996 31272
rect 55956 31220 56008 31272
rect 57428 31263 57480 31272
rect 57428 31229 57437 31263
rect 57437 31229 57471 31263
rect 57471 31229 57480 31263
rect 57428 31220 57480 31229
rect 55220 31152 55272 31204
rect 55680 31152 55732 31204
rect 52092 31084 52144 31136
rect 52828 31084 52880 31136
rect 52920 31084 52972 31136
rect 56416 31084 56468 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 50712 30880 50764 30932
rect 52184 30923 52236 30932
rect 52184 30889 52193 30923
rect 52193 30889 52227 30923
rect 52227 30889 52236 30923
rect 52184 30880 52236 30889
rect 52368 30880 52420 30932
rect 55404 30923 55456 30932
rect 55404 30889 55413 30923
rect 55413 30889 55447 30923
rect 55447 30889 55456 30923
rect 55404 30880 55456 30889
rect 49056 30812 49108 30864
rect 1400 30787 1452 30796
rect 1400 30753 1409 30787
rect 1409 30753 1443 30787
rect 1443 30753 1452 30787
rect 1400 30744 1452 30753
rect 52000 30812 52052 30864
rect 50528 30787 50580 30796
rect 50528 30753 50537 30787
rect 50537 30753 50571 30787
rect 50571 30753 50580 30787
rect 50528 30744 50580 30753
rect 50620 30744 50672 30796
rect 51724 30787 51776 30796
rect 51724 30753 51733 30787
rect 51733 30753 51767 30787
rect 51767 30753 51776 30787
rect 51724 30744 51776 30753
rect 52368 30744 52420 30796
rect 52644 30787 52696 30796
rect 52644 30753 52653 30787
rect 52653 30753 52687 30787
rect 52687 30753 52696 30787
rect 52828 30787 52880 30796
rect 52644 30744 52696 30753
rect 52828 30753 52837 30787
rect 52837 30753 52871 30787
rect 52871 30753 52880 30787
rect 52828 30744 52880 30753
rect 53656 30744 53708 30796
rect 53840 30787 53892 30796
rect 53840 30753 53849 30787
rect 53849 30753 53883 30787
rect 53883 30753 53892 30787
rect 54484 30787 54536 30796
rect 53840 30744 53892 30753
rect 54484 30753 54493 30787
rect 54493 30753 54527 30787
rect 54527 30753 54536 30787
rect 54484 30744 54536 30753
rect 54576 30787 54628 30796
rect 54576 30753 54585 30787
rect 54585 30753 54619 30787
rect 54619 30753 54628 30787
rect 54576 30744 54628 30753
rect 54760 30744 54812 30796
rect 55312 30787 55364 30796
rect 55312 30753 55321 30787
rect 55321 30753 55355 30787
rect 55355 30753 55364 30787
rect 55312 30744 55364 30753
rect 55496 30787 55548 30796
rect 55496 30753 55505 30787
rect 55505 30753 55539 30787
rect 55539 30753 55548 30787
rect 55496 30744 55548 30753
rect 57244 30787 57296 30796
rect 57244 30753 57253 30787
rect 57253 30753 57287 30787
rect 57287 30753 57296 30787
rect 57244 30744 57296 30753
rect 57980 30787 58032 30796
rect 57980 30753 57989 30787
rect 57989 30753 58023 30787
rect 58023 30753 58032 30787
rect 57980 30744 58032 30753
rect 51448 30608 51500 30660
rect 52920 30608 52972 30660
rect 54208 30608 54260 30660
rect 56048 30676 56100 30728
rect 56508 30608 56560 30660
rect 57428 30651 57480 30660
rect 57428 30617 57437 30651
rect 57437 30617 57471 30651
rect 57471 30617 57480 30651
rect 57428 30608 57480 30617
rect 58164 30651 58216 30660
rect 58164 30617 58173 30651
rect 58173 30617 58207 30651
rect 58207 30617 58216 30651
rect 58164 30608 58216 30617
rect 51264 30540 51316 30592
rect 57520 30540 57572 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 49056 30336 49108 30388
rect 48780 30200 48832 30252
rect 49516 30243 49568 30252
rect 49516 30209 49525 30243
rect 49525 30209 49559 30243
rect 49559 30209 49568 30243
rect 49516 30200 49568 30209
rect 51540 30336 51592 30388
rect 52644 30336 52696 30388
rect 52276 30268 52328 30320
rect 52368 30268 52420 30320
rect 53472 30336 53524 30388
rect 54760 30336 54812 30388
rect 55128 30379 55180 30388
rect 55128 30345 55137 30379
rect 55137 30345 55171 30379
rect 55171 30345 55180 30379
rect 55128 30336 55180 30345
rect 55680 30379 55732 30388
rect 55680 30345 55689 30379
rect 55689 30345 55723 30379
rect 55723 30345 55732 30379
rect 55680 30336 55732 30345
rect 57980 30379 58032 30388
rect 57980 30345 57989 30379
rect 57989 30345 58023 30379
rect 58023 30345 58032 30379
rect 57980 30336 58032 30345
rect 54024 30243 54076 30252
rect 54024 30209 54033 30243
rect 54033 30209 54067 30243
rect 54067 30209 54076 30243
rect 54024 30200 54076 30209
rect 55128 30200 55180 30252
rect 57520 30243 57572 30252
rect 47860 30132 47912 30184
rect 52368 30132 52420 30184
rect 52460 30132 52512 30184
rect 54208 30175 54260 30184
rect 1860 30107 1912 30116
rect 1860 30073 1869 30107
rect 1869 30073 1903 30107
rect 1903 30073 1912 30107
rect 1860 30064 1912 30073
rect 49424 30064 49476 30116
rect 49884 30064 49936 30116
rect 54208 30141 54217 30175
rect 54217 30141 54251 30175
rect 54251 30141 54260 30175
rect 54208 30132 54260 30141
rect 54668 30132 54720 30184
rect 55312 30132 55364 30184
rect 57520 30209 57529 30243
rect 57529 30209 57563 30243
rect 57563 30209 57572 30243
rect 57520 30200 57572 30209
rect 1952 30039 2004 30048
rect 1952 30005 1961 30039
rect 1961 30005 1995 30039
rect 1995 30005 2004 30039
rect 1952 29996 2004 30005
rect 48872 30039 48924 30048
rect 48872 30005 48881 30039
rect 48881 30005 48915 30039
rect 48915 30005 48924 30039
rect 48872 29996 48924 30005
rect 48964 29996 49016 30048
rect 50160 29996 50212 30048
rect 50620 29996 50672 30048
rect 50896 30039 50948 30048
rect 50896 30005 50905 30039
rect 50905 30005 50939 30039
rect 50939 30005 50948 30039
rect 50896 29996 50948 30005
rect 54116 29996 54168 30048
rect 56784 30064 56836 30116
rect 56876 30064 56928 30116
rect 57520 29996 57572 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 49424 29835 49476 29844
rect 49424 29801 49433 29835
rect 49433 29801 49467 29835
rect 49467 29801 49476 29835
rect 49424 29792 49476 29801
rect 2136 29656 2188 29708
rect 48964 29656 49016 29708
rect 51264 29724 51316 29776
rect 52000 29724 52052 29776
rect 52828 29724 52880 29776
rect 53288 29767 53340 29776
rect 53288 29733 53297 29767
rect 53297 29733 53331 29767
rect 53331 29733 53340 29767
rect 53288 29724 53340 29733
rect 54944 29724 54996 29776
rect 49976 29631 50028 29640
rect 49976 29597 49985 29631
rect 49985 29597 50019 29631
rect 50019 29597 50028 29631
rect 49976 29588 50028 29597
rect 50896 29656 50948 29708
rect 52368 29699 52420 29708
rect 52368 29665 52377 29699
rect 52377 29665 52411 29699
rect 52411 29665 52420 29699
rect 52368 29656 52420 29665
rect 52460 29656 52512 29708
rect 50436 29588 50488 29640
rect 52276 29631 52328 29640
rect 52276 29597 52285 29631
rect 52285 29597 52319 29631
rect 52319 29597 52328 29631
rect 54024 29656 54076 29708
rect 54852 29656 54904 29708
rect 58256 29792 58308 29844
rect 54208 29631 54260 29640
rect 52276 29588 52328 29597
rect 54208 29597 54217 29631
rect 54217 29597 54251 29631
rect 54251 29597 54260 29631
rect 54208 29588 54260 29597
rect 53748 29520 53800 29572
rect 57888 29656 57940 29708
rect 55956 29588 56008 29640
rect 57244 29563 57296 29572
rect 57244 29529 57253 29563
rect 57253 29529 57287 29563
rect 57287 29529 57296 29563
rect 57244 29520 57296 29529
rect 1400 29452 1452 29504
rect 2688 29495 2740 29504
rect 2688 29461 2697 29495
rect 2697 29461 2731 29495
rect 2731 29461 2740 29495
rect 2688 29452 2740 29461
rect 51540 29495 51592 29504
rect 51540 29461 51549 29495
rect 51549 29461 51583 29495
rect 51583 29461 51592 29495
rect 51540 29452 51592 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1860 29248 1912 29300
rect 48320 29248 48372 29300
rect 49884 29248 49936 29300
rect 49976 29248 50028 29300
rect 50436 29248 50488 29300
rect 50620 29180 50672 29232
rect 2688 29112 2740 29164
rect 49516 29155 49568 29164
rect 49516 29121 49525 29155
rect 49525 29121 49559 29155
rect 49559 29121 49568 29155
rect 49516 29112 49568 29121
rect 1768 29087 1820 29096
rect 1768 29053 1777 29087
rect 1777 29053 1811 29087
rect 1811 29053 1820 29087
rect 1768 29044 1820 29053
rect 47860 29087 47912 29096
rect 47860 29053 47869 29087
rect 47869 29053 47903 29087
rect 47903 29053 47912 29087
rect 47860 29044 47912 29053
rect 49056 29044 49108 29096
rect 50712 29112 50764 29164
rect 51540 29248 51592 29300
rect 54024 29291 54076 29300
rect 54024 29257 54033 29291
rect 54033 29257 54067 29291
rect 54067 29257 54076 29291
rect 54024 29248 54076 29257
rect 56876 29248 56928 29300
rect 57612 29248 57664 29300
rect 51448 29180 51500 29232
rect 55496 29180 55548 29232
rect 56508 29223 56560 29232
rect 56508 29189 56517 29223
rect 56517 29189 56551 29223
rect 56551 29189 56560 29223
rect 56508 29180 56560 29189
rect 50896 29044 50948 29096
rect 51448 29087 51500 29096
rect 51448 29053 51457 29087
rect 51457 29053 51491 29087
rect 51491 29053 51500 29087
rect 51448 29044 51500 29053
rect 52368 29112 52420 29164
rect 51724 29087 51776 29096
rect 51724 29053 51733 29087
rect 51733 29053 51767 29087
rect 51767 29053 51776 29087
rect 51724 29044 51776 29053
rect 51172 28976 51224 29028
rect 52000 29044 52052 29096
rect 52644 29044 52696 29096
rect 51908 28976 51960 29028
rect 53748 29112 53800 29164
rect 53472 29044 53524 29096
rect 54116 29044 54168 29096
rect 54944 29087 54996 29096
rect 54944 29053 54953 29087
rect 54953 29053 54987 29087
rect 54987 29053 54996 29087
rect 54944 29044 54996 29053
rect 55128 29087 55180 29096
rect 55128 29053 55137 29087
rect 55137 29053 55171 29087
rect 55171 29053 55180 29087
rect 55128 29044 55180 29053
rect 56232 29044 56284 29096
rect 56416 29087 56468 29096
rect 56416 29053 56425 29087
rect 56425 29053 56459 29087
rect 56459 29053 56468 29087
rect 56416 29044 56468 29053
rect 57888 29044 57940 29096
rect 55220 28976 55272 29028
rect 57980 29019 58032 29028
rect 57980 28985 57989 29019
rect 57989 28985 58023 29019
rect 58023 28985 58032 29019
rect 57980 28976 58032 28985
rect 58164 29019 58216 29028
rect 58164 28985 58173 29019
rect 58173 28985 58207 29019
rect 58207 28985 58216 29019
rect 58164 28976 58216 28985
rect 49240 28908 49292 28960
rect 50988 28908 51040 28960
rect 51724 28908 51776 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 50326 28806 50378 28858
rect 50390 28806 50442 28858
rect 50454 28806 50506 28858
rect 50518 28806 50570 28858
rect 47860 28704 47912 28756
rect 3976 28568 4028 28620
rect 49424 28704 49476 28756
rect 51448 28704 51500 28756
rect 52460 28747 52512 28756
rect 51632 28636 51684 28688
rect 52460 28713 52469 28747
rect 52469 28713 52503 28747
rect 52503 28713 52512 28747
rect 52460 28704 52512 28713
rect 55128 28704 55180 28756
rect 57980 28704 58032 28756
rect 49056 28611 49108 28620
rect 3148 28500 3200 28552
rect 49056 28577 49065 28611
rect 49065 28577 49099 28611
rect 49099 28577 49108 28611
rect 49056 28568 49108 28577
rect 49240 28611 49292 28620
rect 49240 28577 49249 28611
rect 49249 28577 49283 28611
rect 49283 28577 49292 28611
rect 49240 28568 49292 28577
rect 49700 28611 49752 28620
rect 49700 28577 49709 28611
rect 49709 28577 49743 28611
rect 49743 28577 49752 28611
rect 49700 28568 49752 28577
rect 49976 28568 50028 28620
rect 50620 28568 50672 28620
rect 51724 28611 51776 28620
rect 51724 28577 51733 28611
rect 51733 28577 51767 28611
rect 51767 28577 51776 28611
rect 51724 28568 51776 28577
rect 51908 28611 51960 28620
rect 51908 28577 51917 28611
rect 51917 28577 51951 28611
rect 51951 28577 51960 28611
rect 51908 28568 51960 28577
rect 55312 28636 55364 28688
rect 52184 28568 52236 28620
rect 52460 28568 52512 28620
rect 48872 28500 48924 28552
rect 53196 28500 53248 28552
rect 2136 28475 2188 28484
rect 2136 28441 2145 28475
rect 2145 28441 2179 28475
rect 2179 28441 2188 28475
rect 2136 28432 2188 28441
rect 52184 28432 52236 28484
rect 52920 28432 52972 28484
rect 48780 28364 48832 28416
rect 54208 28364 54260 28416
rect 54300 28364 54352 28416
rect 56876 28611 56928 28620
rect 56876 28577 56885 28611
rect 56885 28577 56919 28611
rect 56919 28577 56928 28611
rect 56876 28568 56928 28577
rect 57060 28611 57112 28620
rect 57060 28577 57069 28611
rect 57069 28577 57103 28611
rect 57103 28577 57112 28611
rect 57060 28568 57112 28577
rect 57520 28611 57572 28620
rect 57520 28577 57529 28611
rect 57529 28577 57563 28611
rect 57563 28577 57572 28611
rect 57520 28568 57572 28577
rect 56600 28500 56652 28552
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1768 28160 1820 28212
rect 3148 28203 3200 28212
rect 3148 28169 3157 28203
rect 3157 28169 3191 28203
rect 3191 28169 3200 28203
rect 3148 28160 3200 28169
rect 3976 28203 4028 28212
rect 3976 28169 3985 28203
rect 3985 28169 4019 28203
rect 4019 28169 4028 28203
rect 3976 28160 4028 28169
rect 50620 28160 50672 28212
rect 52460 28203 52512 28212
rect 52460 28169 52469 28203
rect 52469 28169 52503 28203
rect 52503 28169 52512 28203
rect 52460 28160 52512 28169
rect 52828 28092 52880 28144
rect 2688 27999 2740 28008
rect 2688 27965 2697 27999
rect 2697 27965 2731 27999
rect 2731 27965 2740 27999
rect 2688 27956 2740 27965
rect 48780 27999 48832 28008
rect 48780 27965 48789 27999
rect 48789 27965 48823 27999
rect 48823 27965 48832 27999
rect 48780 27956 48832 27965
rect 2044 27888 2096 27940
rect 1952 27863 2004 27872
rect 1952 27829 1961 27863
rect 1961 27829 1995 27863
rect 1995 27829 2004 27863
rect 1952 27820 2004 27829
rect 50712 27956 50764 28008
rect 51080 27956 51132 28008
rect 51540 27956 51592 28008
rect 52276 27956 52328 28008
rect 52736 27999 52788 28008
rect 52736 27965 52745 27999
rect 52745 27965 52779 27999
rect 52779 27965 52788 27999
rect 52736 27956 52788 27965
rect 53012 27956 53064 28008
rect 56876 28160 56928 28212
rect 54208 28092 54260 28144
rect 55128 28092 55180 28144
rect 54668 28024 54720 28076
rect 55036 27956 55088 28008
rect 55220 27956 55272 28008
rect 57244 27999 57296 28008
rect 49240 27820 49292 27872
rect 52184 27888 52236 27940
rect 57244 27965 57253 27999
rect 57253 27965 57287 27999
rect 57287 27965 57296 27999
rect 57244 27956 57296 27965
rect 53472 27820 53524 27872
rect 54024 27863 54076 27872
rect 54024 27829 54033 27863
rect 54033 27829 54067 27863
rect 54067 27829 54076 27863
rect 54024 27820 54076 27829
rect 56508 27863 56560 27872
rect 56508 27829 56517 27863
rect 56517 27829 56551 27863
rect 56551 27829 56560 27863
rect 56508 27820 56560 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 50326 27718 50378 27770
rect 50390 27718 50442 27770
rect 50454 27718 50506 27770
rect 50518 27718 50570 27770
rect 49700 27616 49752 27668
rect 49884 27616 49936 27668
rect 3332 27480 3384 27532
rect 48320 27480 48372 27532
rect 49056 27523 49108 27532
rect 49056 27489 49065 27523
rect 49065 27489 49099 27523
rect 49099 27489 49108 27523
rect 49056 27480 49108 27489
rect 50252 27548 50304 27600
rect 49976 27480 50028 27532
rect 50160 27480 50212 27532
rect 51264 27616 51316 27668
rect 53472 27659 53524 27668
rect 53472 27625 53481 27659
rect 53481 27625 53515 27659
rect 53515 27625 53524 27659
rect 53472 27616 53524 27625
rect 2504 27412 2556 27464
rect 51724 27480 51776 27532
rect 51816 27480 51868 27532
rect 52736 27548 52788 27600
rect 52828 27548 52880 27600
rect 54300 27523 54352 27532
rect 54300 27489 54309 27523
rect 54309 27489 54343 27523
rect 54343 27489 54352 27523
rect 54300 27480 54352 27489
rect 55220 27548 55272 27600
rect 57060 27591 57112 27600
rect 57060 27557 57069 27591
rect 57069 27557 57103 27591
rect 57103 27557 57112 27591
rect 57060 27548 57112 27557
rect 54668 27523 54720 27532
rect 54668 27489 54677 27523
rect 54677 27489 54711 27523
rect 54711 27489 54720 27523
rect 54668 27480 54720 27489
rect 55312 27523 55364 27532
rect 55312 27489 55321 27523
rect 55321 27489 55355 27523
rect 55355 27489 55364 27523
rect 55312 27480 55364 27489
rect 55496 27523 55548 27532
rect 55496 27489 55505 27523
rect 55505 27489 55539 27523
rect 55539 27489 55548 27523
rect 55496 27480 55548 27489
rect 55680 27523 55732 27532
rect 55680 27489 55689 27523
rect 55689 27489 55723 27523
rect 55723 27489 55732 27523
rect 55680 27480 55732 27489
rect 51172 27412 51224 27464
rect 52736 27455 52788 27464
rect 52736 27421 52745 27455
rect 52745 27421 52779 27455
rect 52779 27421 52788 27455
rect 52736 27412 52788 27421
rect 54116 27412 54168 27464
rect 54208 27412 54260 27464
rect 54576 27455 54628 27464
rect 54576 27421 54585 27455
rect 54585 27421 54619 27455
rect 54619 27421 54628 27455
rect 54576 27412 54628 27421
rect 57704 27455 57756 27464
rect 2044 27387 2096 27396
rect 2044 27353 2053 27387
rect 2053 27353 2087 27387
rect 2087 27353 2096 27387
rect 2044 27344 2096 27353
rect 53012 27344 53064 27396
rect 53196 27344 53248 27396
rect 48412 27319 48464 27328
rect 48412 27285 48421 27319
rect 48421 27285 48455 27319
rect 48455 27285 48464 27319
rect 48412 27276 48464 27285
rect 49608 27276 49660 27328
rect 51632 27276 51684 27328
rect 52000 27276 52052 27328
rect 52368 27319 52420 27328
rect 52368 27285 52377 27319
rect 52377 27285 52411 27319
rect 52411 27285 52420 27319
rect 52368 27276 52420 27285
rect 52644 27276 52696 27328
rect 52828 27276 52880 27328
rect 57704 27421 57713 27455
rect 57713 27421 57747 27455
rect 57747 27421 57756 27455
rect 57704 27412 57756 27421
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 2504 27115 2556 27124
rect 2504 27081 2513 27115
rect 2513 27081 2547 27115
rect 2547 27081 2556 27115
rect 2504 27072 2556 27081
rect 3332 27115 3384 27124
rect 3332 27081 3341 27115
rect 3341 27081 3375 27115
rect 3375 27081 3384 27115
rect 3332 27072 3384 27081
rect 49884 27072 49936 27124
rect 51632 27072 51684 27124
rect 54116 27115 54168 27124
rect 52736 27004 52788 27056
rect 54116 27081 54125 27115
rect 54125 27081 54159 27115
rect 54159 27081 54168 27115
rect 54116 27072 54168 27081
rect 55680 27072 55732 27124
rect 57244 27004 57296 27056
rect 51172 26936 51224 26988
rect 2688 26911 2740 26920
rect 2688 26877 2697 26911
rect 2697 26877 2731 26911
rect 2731 26877 2740 26911
rect 2688 26868 2740 26877
rect 2872 26868 2924 26920
rect 49240 26911 49292 26920
rect 49240 26877 49249 26911
rect 49249 26877 49283 26911
rect 49283 26877 49292 26911
rect 49240 26868 49292 26877
rect 50988 26868 51040 26920
rect 52368 26936 52420 26988
rect 54208 26936 54260 26988
rect 51724 26911 51776 26920
rect 2320 26800 2372 26852
rect 51724 26877 51733 26911
rect 51733 26877 51767 26911
rect 51767 26877 51776 26911
rect 51724 26868 51776 26877
rect 53012 26868 53064 26920
rect 53196 26868 53248 26920
rect 55220 26936 55272 26988
rect 55312 26868 55364 26920
rect 56508 26868 56560 26920
rect 57152 26911 57204 26920
rect 57152 26877 57161 26911
rect 57161 26877 57195 26911
rect 57195 26877 57204 26911
rect 57152 26868 57204 26877
rect 52644 26800 52696 26852
rect 1952 26775 2004 26784
rect 1952 26741 1961 26775
rect 1961 26741 1995 26775
rect 1995 26741 2004 26775
rect 1952 26732 2004 26741
rect 50620 26775 50672 26784
rect 50620 26741 50629 26775
rect 50629 26741 50663 26775
rect 50663 26741 50672 26775
rect 50620 26732 50672 26741
rect 53932 26800 53984 26852
rect 54300 26800 54352 26852
rect 55036 26843 55088 26852
rect 55036 26809 55045 26843
rect 55045 26809 55079 26843
rect 55079 26809 55088 26843
rect 55036 26800 55088 26809
rect 55220 26800 55272 26852
rect 53012 26775 53064 26784
rect 53012 26741 53021 26775
rect 53021 26741 53055 26775
rect 53055 26741 53064 26775
rect 53012 26732 53064 26741
rect 54024 26732 54076 26784
rect 54576 26732 54628 26784
rect 57244 26732 57296 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 50326 26630 50378 26682
rect 50390 26630 50442 26682
rect 50454 26630 50506 26682
rect 50518 26630 50570 26682
rect 2320 26571 2372 26580
rect 2320 26537 2329 26571
rect 2329 26537 2363 26571
rect 2363 26537 2372 26571
rect 2320 26528 2372 26537
rect 50988 26528 51040 26580
rect 54300 26571 54352 26580
rect 54300 26537 54309 26571
rect 54309 26537 54343 26571
rect 54343 26537 54352 26571
rect 54300 26528 54352 26537
rect 55036 26528 55088 26580
rect 55496 26528 55548 26580
rect 57336 26571 57388 26580
rect 57336 26537 57345 26571
rect 57345 26537 57379 26571
rect 57379 26537 57388 26571
rect 57336 26528 57388 26537
rect 55220 26460 55272 26512
rect 49976 26392 50028 26444
rect 50620 26392 50672 26444
rect 51724 26435 51776 26444
rect 51724 26401 51733 26435
rect 51733 26401 51767 26435
rect 51767 26401 51776 26435
rect 51724 26392 51776 26401
rect 51908 26392 51960 26444
rect 52920 26435 52972 26444
rect 52920 26401 52929 26435
rect 52929 26401 52963 26435
rect 52963 26401 52972 26435
rect 52920 26392 52972 26401
rect 54116 26392 54168 26444
rect 54392 26392 54444 26444
rect 57244 26503 57296 26512
rect 57244 26469 57253 26503
rect 57253 26469 57287 26503
rect 57287 26469 57296 26503
rect 57244 26460 57296 26469
rect 57980 26435 58032 26444
rect 1860 26367 1912 26376
rect 1860 26333 1869 26367
rect 1869 26333 1903 26367
rect 1903 26333 1912 26367
rect 1860 26324 1912 26333
rect 50160 26324 50212 26376
rect 54208 26324 54260 26376
rect 54852 26324 54904 26376
rect 57980 26401 57989 26435
rect 57989 26401 58023 26435
rect 58023 26401 58032 26435
rect 57980 26392 58032 26401
rect 52828 26256 52880 26308
rect 49424 26188 49476 26240
rect 51816 26188 51868 26240
rect 52000 26188 52052 26240
rect 52460 26188 52512 26240
rect 55496 26256 55548 26308
rect 57888 26256 57940 26308
rect 55312 26188 55364 26240
rect 56324 26188 56376 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 1860 25984 1912 26036
rect 1308 25916 1360 25968
rect 46204 25984 46256 26036
rect 49240 25984 49292 26036
rect 50620 25984 50672 26036
rect 51724 25984 51776 26036
rect 1860 25755 1912 25764
rect 1860 25721 1869 25755
rect 1869 25721 1903 25755
rect 1903 25721 1912 25755
rect 1860 25712 1912 25721
rect 2044 25755 2096 25764
rect 2044 25721 2053 25755
rect 2053 25721 2087 25755
rect 2087 25721 2096 25755
rect 2044 25712 2096 25721
rect 2780 25780 2832 25832
rect 50160 25823 50212 25832
rect 3148 25712 3200 25764
rect 50160 25789 50169 25823
rect 50169 25789 50203 25823
rect 50203 25789 50212 25823
rect 50160 25780 50212 25789
rect 50620 25823 50672 25832
rect 50620 25789 50629 25823
rect 50629 25789 50663 25823
rect 50663 25789 50672 25823
rect 50620 25780 50672 25789
rect 52092 25984 52144 26036
rect 52092 25848 52144 25900
rect 57152 25984 57204 26036
rect 57980 26027 58032 26036
rect 57980 25993 57989 26027
rect 57989 25993 58023 26027
rect 58023 25993 58032 26027
rect 57980 25984 58032 25993
rect 56324 25959 56376 25968
rect 56324 25925 56333 25959
rect 56333 25925 56367 25959
rect 56367 25925 56376 25959
rect 56324 25916 56376 25925
rect 52736 25848 52788 25900
rect 54300 25823 54352 25832
rect 54300 25789 54309 25823
rect 54309 25789 54343 25823
rect 54343 25789 54352 25823
rect 54300 25780 54352 25789
rect 54760 25780 54812 25832
rect 56600 25848 56652 25900
rect 57704 25823 57756 25832
rect 51080 25712 51132 25764
rect 51632 25712 51684 25764
rect 54852 25712 54904 25764
rect 55036 25712 55088 25764
rect 55128 25712 55180 25764
rect 55312 25712 55364 25764
rect 57704 25789 57713 25823
rect 57713 25789 57747 25823
rect 57747 25789 57756 25823
rect 57704 25780 57756 25789
rect 52460 25644 52512 25696
rect 54392 25687 54444 25696
rect 54392 25653 54401 25687
rect 54401 25653 54435 25687
rect 54435 25653 54444 25687
rect 54392 25644 54444 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 50326 25542 50378 25594
rect 50390 25542 50442 25594
rect 50454 25542 50506 25594
rect 50518 25542 50570 25594
rect 1860 25440 1912 25492
rect 51816 25440 51868 25492
rect 55128 25483 55180 25492
rect 55128 25449 55137 25483
rect 55137 25449 55171 25483
rect 55171 25449 55180 25483
rect 55128 25440 55180 25449
rect 46204 25372 46256 25424
rect 54392 25372 54444 25424
rect 58164 25415 58216 25424
rect 2780 25304 2832 25356
rect 3148 25347 3200 25356
rect 3148 25313 3157 25347
rect 3157 25313 3191 25347
rect 3191 25313 3200 25347
rect 3148 25304 3200 25313
rect 49056 25304 49108 25356
rect 51632 25304 51684 25356
rect 52000 25304 52052 25356
rect 54944 25304 54996 25356
rect 58164 25381 58173 25415
rect 58173 25381 58207 25415
rect 58207 25381 58216 25415
rect 58164 25372 58216 25381
rect 56692 25304 56744 25356
rect 55312 25236 55364 25288
rect 52092 25100 52144 25152
rect 52736 25100 52788 25152
rect 53656 25168 53708 25220
rect 57704 25100 57756 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 50804 24896 50856 24948
rect 53656 24896 53708 24948
rect 2780 24803 2832 24812
rect 2780 24769 2789 24803
rect 2789 24769 2823 24803
rect 2823 24769 2832 24803
rect 2780 24760 2832 24769
rect 3148 24692 3200 24744
rect 50160 24735 50212 24744
rect 50160 24701 50169 24735
rect 50169 24701 50203 24735
rect 50203 24701 50212 24735
rect 50160 24692 50212 24701
rect 50620 24692 50672 24744
rect 55220 24896 55272 24948
rect 53840 24760 53892 24812
rect 54116 24803 54168 24812
rect 54116 24769 54125 24803
rect 54125 24769 54159 24803
rect 54159 24769 54168 24803
rect 54116 24760 54168 24769
rect 53932 24692 53984 24744
rect 54760 24760 54812 24812
rect 57336 24692 57388 24744
rect 58348 24692 58400 24744
rect 2044 24624 2096 24676
rect 2596 24667 2648 24676
rect 2596 24633 2605 24667
rect 2605 24633 2639 24667
rect 2639 24633 2648 24667
rect 2596 24624 2648 24633
rect 50068 24624 50120 24676
rect 50988 24624 51040 24676
rect 51080 24667 51132 24676
rect 51080 24633 51089 24667
rect 51089 24633 51123 24667
rect 51123 24633 51132 24667
rect 51080 24624 51132 24633
rect 52368 24624 52420 24676
rect 1952 24599 2004 24608
rect 1952 24565 1961 24599
rect 1961 24565 1995 24599
rect 1995 24565 2004 24599
rect 1952 24556 2004 24565
rect 3240 24599 3292 24608
rect 3240 24565 3249 24599
rect 3249 24565 3283 24599
rect 3283 24565 3292 24599
rect 3240 24556 3292 24565
rect 49976 24556 50028 24608
rect 54852 24624 54904 24676
rect 55036 24624 55088 24676
rect 56232 24624 56284 24676
rect 57980 24667 58032 24676
rect 53748 24556 53800 24608
rect 54208 24556 54260 24608
rect 55956 24556 56008 24608
rect 57980 24633 57989 24667
rect 57989 24633 58023 24667
rect 58023 24633 58032 24667
rect 57980 24624 58032 24633
rect 58164 24667 58216 24676
rect 58164 24633 58173 24667
rect 58173 24633 58207 24667
rect 58207 24633 58216 24667
rect 58164 24624 58216 24633
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 50326 24454 50378 24506
rect 50390 24454 50442 24506
rect 50454 24454 50506 24506
rect 50518 24454 50570 24506
rect 2596 24352 2648 24404
rect 51908 24395 51960 24404
rect 51908 24361 51917 24395
rect 51917 24361 51951 24395
rect 51951 24361 51960 24395
rect 51908 24352 51960 24361
rect 53012 24327 53064 24336
rect 52092 24259 52144 24268
rect 52092 24225 52101 24259
rect 52101 24225 52135 24259
rect 52135 24225 52144 24259
rect 52092 24216 52144 24225
rect 53012 24293 53021 24327
rect 53021 24293 53055 24327
rect 53055 24293 53064 24327
rect 53012 24284 53064 24293
rect 3240 24148 3292 24200
rect 52828 24148 52880 24200
rect 54576 24352 54628 24404
rect 54668 24284 54720 24336
rect 53748 24259 53800 24268
rect 53748 24225 53757 24259
rect 53757 24225 53791 24259
rect 53791 24225 53800 24259
rect 53748 24216 53800 24225
rect 54576 24216 54628 24268
rect 57980 24352 58032 24404
rect 56876 24259 56928 24268
rect 56876 24225 56885 24259
rect 56885 24225 56919 24259
rect 56919 24225 56928 24259
rect 56876 24216 56928 24225
rect 54208 24191 54260 24200
rect 54208 24157 54217 24191
rect 54217 24157 54251 24191
rect 54251 24157 54260 24191
rect 54208 24148 54260 24157
rect 57704 24191 57756 24200
rect 57704 24157 57713 24191
rect 57713 24157 57747 24191
rect 57747 24157 57756 24191
rect 57704 24148 57756 24157
rect 52460 24012 52512 24064
rect 55128 24012 55180 24064
rect 56968 24055 57020 24064
rect 56968 24021 56977 24055
rect 56977 24021 57011 24055
rect 57011 24021 57020 24055
rect 56968 24012 57020 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 2044 23851 2096 23860
rect 2044 23817 2053 23851
rect 2053 23817 2087 23851
rect 2087 23817 2096 23851
rect 2044 23808 2096 23817
rect 50804 23808 50856 23860
rect 52368 23808 52420 23860
rect 53012 23808 53064 23860
rect 55036 23808 55088 23860
rect 57704 23740 57756 23792
rect 50160 23672 50212 23724
rect 50804 23672 50856 23724
rect 1860 23647 1912 23656
rect 1860 23613 1869 23647
rect 1869 23613 1903 23647
rect 1903 23613 1912 23647
rect 1860 23604 1912 23613
rect 50712 23647 50764 23656
rect 50712 23613 50721 23647
rect 50721 23613 50755 23647
rect 50755 23613 50764 23647
rect 50712 23604 50764 23613
rect 52092 23672 52144 23724
rect 56232 23672 56284 23724
rect 52460 23647 52512 23656
rect 52460 23613 52469 23647
rect 52469 23613 52503 23647
rect 52503 23613 52512 23647
rect 52460 23604 52512 23613
rect 52552 23604 52604 23656
rect 52736 23604 52788 23656
rect 54392 23647 54444 23656
rect 54392 23613 54401 23647
rect 54401 23613 54435 23647
rect 54435 23613 54444 23647
rect 54392 23604 54444 23613
rect 54484 23647 54536 23656
rect 54484 23613 54493 23647
rect 54493 23613 54527 23647
rect 54527 23613 54536 23647
rect 54944 23647 54996 23656
rect 54484 23604 54536 23613
rect 54944 23613 54953 23647
rect 54953 23613 54987 23647
rect 54987 23613 54996 23647
rect 54944 23604 54996 23613
rect 55128 23647 55180 23656
rect 55128 23613 55137 23647
rect 55137 23613 55171 23647
rect 55171 23613 55180 23647
rect 55128 23604 55180 23613
rect 55956 23647 56008 23656
rect 55956 23613 55965 23647
rect 55965 23613 55999 23647
rect 55999 23613 56008 23647
rect 55956 23604 56008 23613
rect 55220 23536 55272 23588
rect 57244 23579 57296 23588
rect 57244 23545 57253 23579
rect 57253 23545 57287 23579
rect 57287 23545 57296 23579
rect 57244 23536 57296 23545
rect 57428 23579 57480 23588
rect 57428 23545 57437 23579
rect 57437 23545 57471 23579
rect 57471 23545 57480 23579
rect 57428 23536 57480 23545
rect 57980 23579 58032 23588
rect 57980 23545 57989 23579
rect 57989 23545 58023 23579
rect 58023 23545 58032 23579
rect 57980 23536 58032 23545
rect 49884 23511 49936 23520
rect 49884 23477 49893 23511
rect 49893 23477 49927 23511
rect 49927 23477 49936 23511
rect 49884 23468 49936 23477
rect 50712 23468 50764 23520
rect 52552 23468 52604 23520
rect 53656 23468 53708 23520
rect 56048 23511 56100 23520
rect 56048 23477 56057 23511
rect 56057 23477 56091 23511
rect 56091 23477 56100 23511
rect 56048 23468 56100 23477
rect 57888 23468 57940 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 50326 23366 50378 23418
rect 50390 23366 50442 23418
rect 50454 23366 50506 23418
rect 50518 23366 50570 23418
rect 1860 23264 1912 23316
rect 49884 23264 49936 23316
rect 50436 23239 50488 23248
rect 50436 23205 50445 23239
rect 50445 23205 50479 23239
rect 50479 23205 50488 23239
rect 50436 23196 50488 23205
rect 1860 23171 1912 23180
rect 1860 23137 1869 23171
rect 1869 23137 1903 23171
rect 1903 23137 1912 23171
rect 1860 23128 1912 23137
rect 3148 23128 3200 23180
rect 49884 23128 49936 23180
rect 52092 23128 52144 23180
rect 54208 23128 54260 23180
rect 54484 23171 54536 23180
rect 54484 23137 54493 23171
rect 54493 23137 54527 23171
rect 54527 23137 54536 23171
rect 54484 23128 54536 23137
rect 56048 23196 56100 23248
rect 55128 23128 55180 23180
rect 55588 23171 55640 23180
rect 55588 23137 55597 23171
rect 55597 23137 55631 23171
rect 55631 23137 55640 23171
rect 55588 23128 55640 23137
rect 57152 23171 57204 23180
rect 57152 23137 57161 23171
rect 57161 23137 57195 23171
rect 57195 23137 57204 23171
rect 57152 23128 57204 23137
rect 49976 23060 50028 23112
rect 54668 23103 54720 23112
rect 54668 23069 54677 23103
rect 54677 23069 54711 23103
rect 54711 23069 54720 23103
rect 54668 23060 54720 23069
rect 1584 22992 1636 23044
rect 53840 22992 53892 23044
rect 54392 22992 54444 23044
rect 56876 22992 56928 23044
rect 1952 22967 2004 22976
rect 1952 22933 1961 22967
rect 1961 22933 1995 22967
rect 1995 22933 2004 22967
rect 1952 22924 2004 22933
rect 49792 22924 49844 22976
rect 52000 22924 52052 22976
rect 54116 22924 54168 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 1860 22720 1912 22772
rect 3148 22720 3200 22772
rect 51724 22720 51776 22772
rect 52092 22763 52144 22772
rect 52092 22729 52101 22763
rect 52101 22729 52135 22763
rect 52135 22729 52144 22763
rect 52092 22720 52144 22729
rect 53748 22720 53800 22772
rect 1584 22627 1636 22636
rect 1584 22593 1593 22627
rect 1593 22593 1627 22627
rect 1627 22593 1636 22627
rect 1584 22584 1636 22593
rect 53748 22584 53800 22636
rect 2964 22516 3016 22568
rect 3148 22516 3200 22568
rect 49884 22516 49936 22568
rect 50620 22516 50672 22568
rect 50712 22516 50764 22568
rect 52368 22559 52420 22568
rect 52368 22525 52377 22559
rect 52377 22525 52411 22559
rect 52411 22525 52420 22559
rect 52368 22516 52420 22525
rect 52736 22559 52788 22568
rect 52276 22448 52328 22500
rect 52736 22525 52745 22559
rect 52745 22525 52779 22559
rect 52779 22525 52788 22559
rect 52736 22516 52788 22525
rect 52644 22448 52696 22500
rect 55588 22720 55640 22772
rect 56232 22763 56284 22772
rect 56232 22729 56241 22763
rect 56241 22729 56275 22763
rect 56275 22729 56284 22763
rect 56232 22720 56284 22729
rect 57244 22720 57296 22772
rect 54116 22559 54168 22568
rect 54116 22525 54125 22559
rect 54125 22525 54159 22559
rect 54159 22525 54168 22559
rect 54116 22516 54168 22525
rect 54852 22559 54904 22568
rect 54852 22525 54861 22559
rect 54861 22525 54895 22559
rect 54895 22525 54904 22559
rect 54852 22516 54904 22525
rect 52000 22380 52052 22432
rect 53380 22380 53432 22432
rect 54208 22423 54260 22432
rect 54208 22389 54217 22423
rect 54217 22389 54251 22423
rect 54251 22389 54260 22423
rect 54208 22380 54260 22389
rect 54944 22448 54996 22500
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 50326 22278 50378 22330
rect 50390 22278 50442 22330
rect 50454 22278 50506 22330
rect 50518 22278 50570 22330
rect 50620 22176 50672 22228
rect 54300 22176 54352 22228
rect 54944 22219 54996 22228
rect 54944 22185 54953 22219
rect 54953 22185 54987 22219
rect 54987 22185 54996 22219
rect 54944 22176 54996 22185
rect 2964 22108 3016 22160
rect 51356 22108 51408 22160
rect 52368 22108 52420 22160
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 49332 22040 49384 22092
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 2044 21947 2096 21956
rect 2044 21913 2053 21947
rect 2053 21913 2087 21947
rect 2087 21913 2096 21947
rect 2044 21904 2096 21913
rect 52552 22040 52604 22092
rect 52828 22083 52880 22092
rect 52828 22049 52837 22083
rect 52837 22049 52871 22083
rect 52871 22049 52880 22083
rect 52828 22040 52880 22049
rect 54208 22108 54260 22160
rect 54024 22083 54076 22092
rect 54024 22049 54033 22083
rect 54033 22049 54067 22083
rect 54067 22049 54076 22083
rect 54024 22040 54076 22049
rect 54760 22040 54812 22092
rect 54944 22040 54996 22092
rect 58072 22108 58124 22160
rect 55128 22040 55180 22092
rect 55680 22083 55732 22092
rect 55680 22049 55689 22083
rect 55689 22049 55723 22083
rect 55723 22049 55732 22083
rect 55680 22040 55732 22049
rect 56232 21972 56284 22024
rect 57704 22015 57756 22024
rect 31300 21836 31352 21888
rect 49056 21879 49108 21888
rect 49056 21845 49065 21879
rect 49065 21845 49099 21879
rect 49099 21845 49108 21879
rect 49056 21836 49108 21845
rect 52644 21836 52696 21888
rect 54116 21904 54168 21956
rect 54300 21947 54352 21956
rect 54300 21913 54309 21947
rect 54309 21913 54343 21947
rect 54343 21913 54352 21947
rect 54300 21904 54352 21913
rect 54392 21904 54444 21956
rect 57704 21981 57713 22015
rect 57713 21981 57747 22015
rect 57747 21981 57756 22015
rect 57704 21972 57756 21981
rect 57980 21947 58032 21956
rect 57980 21913 57989 21947
rect 57989 21913 58023 21947
rect 58023 21913 58032 21947
rect 57980 21904 58032 21913
rect 55220 21836 55272 21888
rect 55496 21879 55548 21888
rect 55496 21845 55505 21879
rect 55505 21845 55539 21879
rect 55539 21845 55548 21879
rect 55496 21836 55548 21845
rect 56508 21836 56560 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 1860 21632 1912 21684
rect 51816 21632 51868 21684
rect 3148 21564 3200 21616
rect 51724 21564 51776 21616
rect 52736 21564 52788 21616
rect 53196 21632 53248 21684
rect 53380 21632 53432 21684
rect 57704 21632 57756 21684
rect 58072 21675 58124 21684
rect 58072 21641 58081 21675
rect 58081 21641 58115 21675
rect 58115 21641 58124 21675
rect 58072 21632 58124 21641
rect 52920 21564 52972 21616
rect 3056 21428 3108 21480
rect 49884 21471 49936 21480
rect 49884 21437 49893 21471
rect 49893 21437 49927 21471
rect 49927 21437 49936 21471
rect 49884 21428 49936 21437
rect 3240 21360 3292 21412
rect 2872 21292 2924 21344
rect 49976 21335 50028 21344
rect 49976 21301 49985 21335
rect 49985 21301 50019 21335
rect 50019 21301 50028 21335
rect 49976 21292 50028 21301
rect 50160 21428 50212 21480
rect 50620 21360 50672 21412
rect 51632 21292 51684 21344
rect 52736 21471 52788 21480
rect 52736 21437 52745 21471
rect 52745 21437 52779 21471
rect 52779 21437 52788 21471
rect 52736 21428 52788 21437
rect 54116 21428 54168 21480
rect 54484 21539 54536 21548
rect 54484 21505 54493 21539
rect 54493 21505 54527 21539
rect 54527 21505 54536 21539
rect 54484 21496 54536 21505
rect 54576 21360 54628 21412
rect 53288 21292 53340 21344
rect 54024 21292 54076 21344
rect 55036 21428 55088 21480
rect 56600 21428 56652 21480
rect 55496 21360 55548 21412
rect 56048 21292 56100 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 50326 21190 50378 21242
rect 50390 21190 50442 21242
rect 50454 21190 50506 21242
rect 50518 21190 50570 21242
rect 1860 20995 1912 21004
rect 1860 20961 1869 20995
rect 1869 20961 1903 20995
rect 1903 20961 1912 20995
rect 1860 20952 1912 20961
rect 2596 20995 2648 21004
rect 2596 20961 2605 20995
rect 2605 20961 2639 20995
rect 2639 20961 2648 20995
rect 2596 20952 2648 20961
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 47860 20952 47912 21004
rect 49976 21088 50028 21140
rect 50620 21020 50672 21072
rect 49056 20952 49108 21004
rect 49792 20952 49844 21004
rect 52552 21020 52604 21072
rect 53288 21063 53340 21072
rect 53288 21029 53297 21063
rect 53297 21029 53331 21063
rect 53331 21029 53340 21063
rect 54116 21088 54168 21140
rect 53288 21020 53340 21029
rect 52644 20995 52696 21004
rect 51264 20884 51316 20936
rect 51724 20816 51776 20868
rect 52644 20961 52653 20995
rect 52653 20961 52687 20995
rect 52687 20961 52696 20995
rect 52644 20952 52696 20961
rect 52552 20884 52604 20936
rect 52736 20884 52788 20936
rect 52920 20995 52972 21004
rect 52920 20961 52929 20995
rect 52929 20961 52963 20995
rect 52963 20961 52972 20995
rect 53748 20995 53800 21004
rect 52920 20952 52972 20961
rect 53748 20961 53757 20995
rect 53757 20961 53791 20995
rect 53791 20961 53800 20995
rect 53748 20952 53800 20961
rect 54300 20995 54352 21004
rect 54300 20961 54309 20995
rect 54309 20961 54343 20995
rect 54343 20961 54352 20995
rect 54300 20952 54352 20961
rect 54576 20952 54628 21004
rect 53104 20884 53156 20936
rect 53656 20884 53708 20936
rect 53840 20816 53892 20868
rect 54116 20927 54168 20936
rect 54116 20893 54125 20927
rect 54125 20893 54159 20927
rect 54159 20893 54168 20927
rect 55680 20952 55732 21004
rect 54116 20884 54168 20893
rect 56048 20884 56100 20936
rect 57244 20927 57296 20936
rect 57244 20893 57253 20927
rect 57253 20893 57287 20927
rect 57287 20893 57296 20927
rect 57244 20884 57296 20893
rect 1952 20791 2004 20800
rect 1952 20757 1961 20791
rect 1961 20757 1995 20791
rect 1995 20757 2004 20791
rect 1952 20748 2004 20757
rect 48412 20791 48464 20800
rect 48412 20757 48421 20791
rect 48421 20757 48455 20791
rect 48455 20757 48464 20791
rect 48412 20748 48464 20757
rect 52000 20791 52052 20800
rect 52000 20757 52009 20791
rect 52009 20757 52043 20791
rect 52043 20757 52052 20791
rect 52000 20748 52052 20757
rect 52920 20748 52972 20800
rect 54300 20816 54352 20868
rect 56600 20816 56652 20868
rect 54024 20748 54076 20800
rect 55496 20791 55548 20800
rect 55496 20757 55505 20791
rect 55505 20757 55539 20791
rect 55539 20757 55548 20791
rect 55496 20748 55548 20757
rect 57428 20791 57480 20800
rect 57428 20757 57437 20791
rect 57437 20757 57471 20791
rect 57471 20757 57480 20791
rect 57428 20748 57480 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 2596 20544 2648 20596
rect 3240 20587 3292 20596
rect 3240 20553 3249 20587
rect 3249 20553 3283 20587
rect 3283 20553 3292 20587
rect 3240 20544 3292 20553
rect 51264 20587 51316 20596
rect 51264 20553 51273 20587
rect 51273 20553 51307 20587
rect 51307 20553 51316 20587
rect 51264 20544 51316 20553
rect 54300 20544 54352 20596
rect 54484 20544 54536 20596
rect 55680 20544 55732 20596
rect 2872 20408 2924 20460
rect 57244 20476 57296 20528
rect 57520 20476 57572 20528
rect 52828 20451 52880 20460
rect 52828 20417 52837 20451
rect 52837 20417 52871 20451
rect 52871 20417 52880 20451
rect 52828 20408 52880 20417
rect 53288 20408 53340 20460
rect 3056 20340 3108 20392
rect 3240 20340 3292 20392
rect 50068 20340 50120 20392
rect 50712 20340 50764 20392
rect 51448 20340 51500 20392
rect 53104 20340 53156 20392
rect 54300 20383 54352 20392
rect 54300 20349 54309 20383
rect 54309 20349 54343 20383
rect 54343 20349 54352 20383
rect 54300 20340 54352 20349
rect 54576 20383 54628 20392
rect 54576 20349 54585 20383
rect 54585 20349 54619 20383
rect 54619 20349 54628 20383
rect 54576 20340 54628 20349
rect 55496 20408 55548 20460
rect 56048 20383 56100 20392
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 50620 20204 50672 20256
rect 50988 20204 51040 20256
rect 51448 20247 51500 20256
rect 51448 20213 51457 20247
rect 51457 20213 51491 20247
rect 51491 20213 51500 20247
rect 51448 20204 51500 20213
rect 52276 20204 52328 20256
rect 52828 20272 52880 20324
rect 54484 20315 54536 20324
rect 54484 20281 54493 20315
rect 54493 20281 54527 20315
rect 54527 20281 54536 20315
rect 54484 20272 54536 20281
rect 56048 20349 56057 20383
rect 56057 20349 56091 20383
rect 56091 20349 56100 20383
rect 56048 20340 56100 20349
rect 57428 20340 57480 20392
rect 57980 20315 58032 20324
rect 57980 20281 57989 20315
rect 57989 20281 58023 20315
rect 58023 20281 58032 20315
rect 57980 20272 58032 20281
rect 58164 20315 58216 20324
rect 58164 20281 58173 20315
rect 58173 20281 58207 20315
rect 58207 20281 58216 20315
rect 58164 20272 58216 20281
rect 54300 20204 54352 20256
rect 55128 20204 55180 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 50326 20102 50378 20154
rect 50390 20102 50442 20154
rect 50454 20102 50506 20154
rect 50518 20102 50570 20154
rect 1860 20000 1912 20052
rect 51448 20000 51500 20052
rect 52276 20000 52328 20052
rect 55312 20000 55364 20052
rect 57980 20000 58032 20052
rect 3884 19932 3936 19984
rect 2964 19864 3016 19916
rect 49056 19864 49108 19916
rect 50712 19864 50764 19916
rect 50896 19864 50948 19916
rect 52368 19907 52420 19916
rect 52368 19873 52377 19907
rect 52377 19873 52411 19907
rect 52411 19873 52420 19907
rect 52368 19864 52420 19873
rect 50068 19796 50120 19848
rect 52276 19796 52328 19848
rect 50620 19728 50672 19780
rect 50896 19728 50948 19780
rect 51448 19728 51500 19780
rect 53012 19864 53064 19916
rect 53104 19907 53156 19916
rect 53104 19873 53113 19907
rect 53113 19873 53147 19907
rect 53147 19873 53156 19907
rect 53104 19864 53156 19873
rect 53380 19907 53432 19916
rect 53380 19873 53414 19907
rect 53414 19873 53432 19907
rect 53380 19864 53432 19873
rect 54760 19864 54812 19916
rect 55128 19907 55180 19916
rect 55128 19873 55137 19907
rect 55137 19873 55171 19907
rect 55171 19873 55180 19907
rect 55128 19864 55180 19873
rect 55220 19864 55272 19916
rect 56876 19907 56928 19916
rect 56876 19873 56885 19907
rect 56885 19873 56919 19907
rect 56919 19873 56928 19907
rect 56876 19864 56928 19873
rect 3240 19660 3292 19712
rect 49056 19703 49108 19712
rect 49056 19669 49065 19703
rect 49065 19669 49099 19703
rect 49099 19669 49108 19703
rect 49056 19660 49108 19669
rect 50068 19660 50120 19712
rect 50712 19660 50764 19712
rect 51540 19660 51592 19712
rect 54392 19796 54444 19848
rect 54208 19660 54260 19712
rect 55128 19728 55180 19780
rect 57060 19771 57112 19780
rect 57060 19737 57069 19771
rect 57069 19737 57103 19771
rect 57103 19737 57112 19771
rect 57060 19728 57112 19737
rect 54484 19703 54536 19712
rect 54484 19669 54493 19703
rect 54493 19669 54527 19703
rect 54527 19669 54536 19703
rect 54484 19660 54536 19669
rect 55220 19660 55272 19712
rect 55312 19660 55364 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 52368 19456 52420 19508
rect 53104 19456 53156 19508
rect 54300 19456 54352 19508
rect 56876 19456 56928 19508
rect 54392 19388 54444 19440
rect 2872 19252 2924 19304
rect 47860 19295 47912 19304
rect 47860 19261 47869 19295
rect 47869 19261 47903 19295
rect 47903 19261 47912 19295
rect 47860 19252 47912 19261
rect 49056 19252 49108 19304
rect 49792 19295 49844 19304
rect 49792 19261 49801 19295
rect 49801 19261 49835 19295
rect 49835 19261 49844 19295
rect 49792 19252 49844 19261
rect 1860 19227 1912 19236
rect 1860 19193 1869 19227
rect 1869 19193 1903 19227
rect 1903 19193 1912 19227
rect 1860 19184 1912 19193
rect 2596 19227 2648 19236
rect 2596 19193 2605 19227
rect 2605 19193 2639 19227
rect 2639 19193 2648 19227
rect 2596 19184 2648 19193
rect 2780 19227 2832 19236
rect 2780 19193 2789 19227
rect 2789 19193 2823 19227
rect 2823 19193 2832 19227
rect 2780 19184 2832 19193
rect 49976 19252 50028 19304
rect 52092 19252 52144 19304
rect 53288 19320 53340 19372
rect 54576 19320 54628 19372
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 49700 19116 49752 19168
rect 50160 19116 50212 19168
rect 51908 19184 51960 19236
rect 52552 19184 52604 19236
rect 53104 19295 53156 19304
rect 53104 19261 53113 19295
rect 53113 19261 53147 19295
rect 53147 19261 53156 19295
rect 53104 19252 53156 19261
rect 54116 19252 54168 19304
rect 54484 19252 54536 19304
rect 54668 19252 54720 19304
rect 55036 19252 55088 19304
rect 55220 19295 55272 19304
rect 55220 19261 55254 19295
rect 55254 19261 55272 19295
rect 55220 19252 55272 19261
rect 56968 19295 57020 19304
rect 56968 19261 56977 19295
rect 56977 19261 57011 19295
rect 57011 19261 57020 19295
rect 56968 19252 57020 19261
rect 57152 19295 57204 19304
rect 57152 19261 57161 19295
rect 57161 19261 57195 19295
rect 57195 19261 57204 19295
rect 57152 19252 57204 19261
rect 53840 19184 53892 19236
rect 54208 19184 54260 19236
rect 54392 19227 54444 19236
rect 54392 19193 54401 19227
rect 54401 19193 54435 19227
rect 54435 19193 54444 19227
rect 54392 19184 54444 19193
rect 54576 19184 54628 19236
rect 55312 19184 55364 19236
rect 50896 19116 50948 19168
rect 51632 19159 51684 19168
rect 51632 19125 51641 19159
rect 51641 19125 51675 19159
rect 51675 19125 51684 19159
rect 51632 19116 51684 19125
rect 52736 19116 52788 19168
rect 53932 19116 53984 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 50326 19014 50378 19066
rect 50390 19014 50442 19066
rect 50454 19014 50506 19066
rect 50518 19014 50570 19066
rect 2596 18955 2648 18964
rect 2596 18921 2605 18955
rect 2605 18921 2639 18955
rect 2639 18921 2648 18955
rect 2596 18912 2648 18921
rect 49976 18912 50028 18964
rect 50712 18912 50764 18964
rect 57152 18912 57204 18964
rect 2872 18776 2924 18828
rect 3240 18819 3292 18828
rect 3240 18785 3249 18819
rect 3249 18785 3283 18819
rect 3283 18785 3292 18819
rect 3240 18776 3292 18785
rect 49056 18776 49108 18828
rect 55220 18844 55272 18896
rect 49884 18776 49936 18828
rect 51448 18776 51500 18828
rect 51632 18819 51684 18828
rect 51632 18785 51641 18819
rect 51641 18785 51675 18819
rect 51675 18785 51684 18819
rect 51632 18776 51684 18785
rect 52644 18776 52696 18828
rect 52920 18819 52972 18828
rect 52920 18785 52929 18819
rect 52929 18785 52963 18819
rect 52963 18785 52972 18819
rect 52920 18776 52972 18785
rect 53380 18776 53432 18828
rect 54116 18819 54168 18828
rect 54116 18785 54125 18819
rect 54125 18785 54159 18819
rect 54159 18785 54168 18819
rect 54116 18776 54168 18785
rect 54300 18776 54352 18828
rect 54392 18776 54444 18828
rect 56692 18844 56744 18896
rect 57336 18844 57388 18896
rect 56140 18776 56192 18828
rect 56784 18819 56836 18828
rect 56784 18785 56793 18819
rect 56793 18785 56827 18819
rect 56827 18785 56836 18819
rect 56784 18776 56836 18785
rect 57980 18819 58032 18828
rect 57980 18785 57989 18819
rect 57989 18785 58023 18819
rect 58023 18785 58032 18819
rect 57980 18776 58032 18785
rect 50620 18708 50672 18760
rect 52276 18708 52328 18760
rect 51080 18640 51132 18692
rect 51264 18640 51316 18692
rect 51448 18572 51500 18624
rect 51816 18572 51868 18624
rect 52828 18615 52880 18624
rect 52828 18581 52837 18615
rect 52837 18581 52871 18615
rect 52871 18581 52880 18615
rect 52828 18572 52880 18581
rect 53288 18572 53340 18624
rect 53932 18615 53984 18624
rect 53932 18581 53941 18615
rect 53941 18581 53975 18615
rect 53975 18581 53984 18615
rect 53932 18572 53984 18581
rect 54208 18572 54260 18624
rect 54392 18615 54444 18624
rect 54392 18581 54401 18615
rect 54401 18581 54435 18615
rect 54435 18581 54444 18615
rect 54392 18572 54444 18581
rect 58164 18683 58216 18692
rect 58164 18649 58173 18683
rect 58173 18649 58207 18683
rect 58207 18649 58216 18683
rect 58164 18640 58216 18649
rect 55588 18572 55640 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 1860 18368 1912 18420
rect 56140 18411 56192 18420
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 51448 18300 51500 18352
rect 51908 18343 51960 18352
rect 51908 18309 51917 18343
rect 51917 18309 51951 18343
rect 51951 18309 51960 18343
rect 51908 18300 51960 18309
rect 53104 18300 53156 18352
rect 56140 18377 56149 18411
rect 56149 18377 56183 18411
rect 56183 18377 56192 18411
rect 56140 18368 56192 18377
rect 57980 18411 58032 18420
rect 57980 18377 57989 18411
rect 57989 18377 58023 18411
rect 58023 18377 58032 18411
rect 57980 18368 58032 18377
rect 52000 18232 52052 18284
rect 50160 18207 50212 18216
rect 50160 18173 50169 18207
rect 50169 18173 50203 18207
rect 50203 18173 50212 18207
rect 50160 18164 50212 18173
rect 50712 18164 50764 18216
rect 51172 18164 51224 18216
rect 51540 18164 51592 18216
rect 52460 18164 52512 18216
rect 54668 18232 54720 18284
rect 53012 18207 53064 18216
rect 52368 18096 52420 18148
rect 49792 18028 49844 18080
rect 50712 18028 50764 18080
rect 51448 18028 51500 18080
rect 53012 18173 53021 18207
rect 53021 18173 53055 18207
rect 53055 18173 53064 18207
rect 53012 18164 53064 18173
rect 53288 18164 53340 18216
rect 54208 18207 54260 18216
rect 54208 18173 54217 18207
rect 54217 18173 54251 18207
rect 54251 18173 54260 18207
rect 54208 18164 54260 18173
rect 52920 18096 52972 18148
rect 53196 18096 53248 18148
rect 55588 18164 55640 18216
rect 57520 18207 57572 18216
rect 57520 18173 57529 18207
rect 57529 18173 57563 18207
rect 57563 18173 57572 18207
rect 57520 18164 57572 18173
rect 54852 18096 54904 18148
rect 56876 18139 56928 18148
rect 56876 18105 56885 18139
rect 56885 18105 56919 18139
rect 56919 18105 56928 18139
rect 56876 18096 56928 18105
rect 57060 18139 57112 18148
rect 57060 18105 57069 18139
rect 57069 18105 57103 18139
rect 57103 18105 57112 18139
rect 57060 18096 57112 18105
rect 52828 18028 52880 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 50326 17926 50378 17978
rect 50390 17926 50442 17978
rect 50454 17926 50506 17978
rect 50518 17926 50570 17978
rect 1768 17824 1820 17876
rect 54852 17867 54904 17876
rect 1860 17731 1912 17740
rect 1860 17697 1869 17731
rect 1869 17697 1903 17731
rect 1903 17697 1912 17731
rect 1860 17688 1912 17697
rect 3240 17688 3292 17740
rect 54852 17833 54861 17867
rect 54861 17833 54895 17867
rect 54895 17833 54904 17867
rect 54852 17824 54904 17833
rect 49792 17688 49844 17740
rect 52736 17756 52788 17808
rect 50528 17731 50580 17740
rect 50528 17697 50537 17731
rect 50537 17697 50571 17731
rect 50571 17697 50580 17731
rect 50528 17688 50580 17697
rect 51172 17688 51224 17740
rect 51724 17731 51776 17740
rect 51724 17697 51733 17731
rect 51733 17697 51767 17731
rect 51767 17697 51776 17731
rect 52000 17731 52052 17740
rect 51724 17688 51776 17697
rect 52000 17697 52009 17731
rect 52009 17697 52043 17731
rect 52043 17697 52052 17731
rect 52000 17688 52052 17697
rect 52460 17731 52512 17740
rect 52460 17697 52469 17731
rect 52469 17697 52503 17731
rect 52503 17697 52512 17731
rect 52460 17688 52512 17697
rect 52552 17688 52604 17740
rect 52828 17731 52880 17740
rect 52828 17697 52837 17731
rect 52837 17697 52871 17731
rect 52871 17697 52880 17731
rect 52828 17688 52880 17697
rect 52920 17688 52972 17740
rect 53380 17688 53432 17740
rect 53932 17731 53984 17740
rect 53932 17697 53941 17731
rect 53941 17697 53975 17731
rect 53975 17697 53984 17731
rect 53932 17688 53984 17697
rect 54760 17731 54812 17740
rect 51356 17620 51408 17672
rect 51448 17620 51500 17672
rect 53472 17620 53524 17672
rect 53840 17620 53892 17672
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 52828 17552 52880 17604
rect 54760 17697 54769 17731
rect 54769 17697 54803 17731
rect 54803 17697 54812 17731
rect 54760 17688 54812 17697
rect 54944 17731 54996 17740
rect 54944 17697 54953 17731
rect 54953 17697 54987 17731
rect 54987 17697 54996 17731
rect 54944 17688 54996 17697
rect 55496 17731 55548 17740
rect 55496 17697 55505 17731
rect 55505 17697 55539 17731
rect 55539 17697 55548 17731
rect 55496 17688 55548 17697
rect 56508 17620 56560 17672
rect 56968 17663 57020 17672
rect 56968 17629 56977 17663
rect 56977 17629 57011 17663
rect 57011 17629 57020 17663
rect 56968 17620 57020 17629
rect 57152 17663 57204 17672
rect 57152 17629 57161 17663
rect 57161 17629 57195 17663
rect 57195 17629 57204 17663
rect 57152 17620 57204 17629
rect 56876 17552 56928 17604
rect 51356 17484 51408 17536
rect 51632 17484 51684 17536
rect 54208 17484 54260 17536
rect 54300 17484 54352 17536
rect 57520 17484 57572 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 1860 17280 1912 17332
rect 2504 17076 2556 17128
rect 55220 17280 55272 17332
rect 55496 17323 55548 17332
rect 55496 17289 55505 17323
rect 55505 17289 55539 17323
rect 55539 17289 55548 17323
rect 55496 17280 55548 17289
rect 55680 17280 55732 17332
rect 51172 17255 51224 17264
rect 51172 17221 51181 17255
rect 51181 17221 51215 17255
rect 51215 17221 51224 17255
rect 51172 17212 51224 17221
rect 51356 17212 51408 17264
rect 49700 17144 49752 17196
rect 51632 17187 51684 17196
rect 51632 17153 51641 17187
rect 51641 17153 51675 17187
rect 51675 17153 51684 17187
rect 51632 17144 51684 17153
rect 54116 17212 54168 17264
rect 53104 17187 53156 17196
rect 52828 17119 52880 17128
rect 50160 17008 50212 17060
rect 52828 17085 52837 17119
rect 52837 17085 52871 17119
rect 52871 17085 52880 17119
rect 52828 17076 52880 17085
rect 53104 17153 53113 17187
rect 53113 17153 53147 17187
rect 53147 17153 53156 17187
rect 53104 17144 53156 17153
rect 53012 17119 53064 17128
rect 53012 17085 53021 17119
rect 53021 17085 53055 17119
rect 53055 17085 53064 17119
rect 53012 17076 53064 17085
rect 53932 17076 53984 17128
rect 54208 17076 54260 17128
rect 55588 17212 55640 17264
rect 56232 17119 56284 17128
rect 56232 17085 56241 17119
rect 56241 17085 56275 17119
rect 56275 17085 56284 17119
rect 56508 17119 56560 17128
rect 56232 17076 56284 17085
rect 56508 17085 56517 17119
rect 56517 17085 56551 17119
rect 56551 17085 56560 17119
rect 56508 17076 56560 17085
rect 53472 17008 53524 17060
rect 54576 17008 54628 17060
rect 55220 17008 55272 17060
rect 57244 17051 57296 17060
rect 57244 17017 57253 17051
rect 57253 17017 57287 17051
rect 57287 17017 57296 17051
rect 57244 17008 57296 17017
rect 57428 17051 57480 17060
rect 57428 17017 57437 17051
rect 57437 17017 57471 17051
rect 57471 17017 57480 17051
rect 57428 17008 57480 17017
rect 57980 17051 58032 17060
rect 57980 17017 57989 17051
rect 57989 17017 58023 17051
rect 58023 17017 58032 17051
rect 57980 17008 58032 17017
rect 58164 17051 58216 17060
rect 58164 17017 58173 17051
rect 58173 17017 58207 17051
rect 58207 17017 58216 17051
rect 58164 17008 58216 17017
rect 50712 16940 50764 16992
rect 52368 16940 52420 16992
rect 56968 16940 57020 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 50326 16838 50378 16890
rect 50390 16838 50442 16890
rect 50454 16838 50506 16890
rect 50518 16838 50570 16890
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 49884 16736 49936 16788
rect 50160 16736 50212 16788
rect 52552 16736 52604 16788
rect 52736 16736 52788 16788
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 3056 16600 3108 16652
rect 49976 16600 50028 16652
rect 50712 16668 50764 16720
rect 53012 16668 53064 16720
rect 54760 16736 54812 16788
rect 51356 16600 51408 16652
rect 51448 16643 51500 16652
rect 51448 16609 51457 16643
rect 51457 16609 51491 16643
rect 51491 16609 51500 16643
rect 51632 16643 51684 16652
rect 51448 16600 51500 16609
rect 51632 16609 51641 16643
rect 51641 16609 51675 16643
rect 51675 16609 51684 16643
rect 51632 16600 51684 16609
rect 52276 16643 52328 16652
rect 52276 16609 52285 16643
rect 52285 16609 52319 16643
rect 52319 16609 52328 16643
rect 52276 16600 52328 16609
rect 52828 16600 52880 16652
rect 53104 16643 53156 16652
rect 53104 16609 53113 16643
rect 53113 16609 53147 16643
rect 53147 16609 53156 16643
rect 53104 16600 53156 16609
rect 51172 16532 51224 16584
rect 52920 16532 52972 16584
rect 53196 16575 53248 16584
rect 53196 16541 53205 16575
rect 53205 16541 53239 16575
rect 53239 16541 53248 16575
rect 53196 16532 53248 16541
rect 53288 16575 53340 16584
rect 53288 16541 53297 16575
rect 53297 16541 53331 16575
rect 53331 16541 53340 16575
rect 54208 16600 54260 16652
rect 54484 16600 54536 16652
rect 55220 16643 55272 16652
rect 55220 16609 55229 16643
rect 55229 16609 55263 16643
rect 55263 16609 55272 16643
rect 55220 16600 55272 16609
rect 56600 16600 56652 16652
rect 57980 16736 58032 16788
rect 53288 16532 53340 16541
rect 1952 16439 2004 16448
rect 1952 16405 1961 16439
rect 1961 16405 1995 16439
rect 1995 16405 2004 16439
rect 1952 16396 2004 16405
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 52460 16439 52512 16448
rect 52460 16405 52469 16439
rect 52469 16405 52503 16439
rect 52503 16405 52512 16439
rect 52460 16396 52512 16405
rect 53012 16396 53064 16448
rect 56692 16396 56744 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 1860 16192 1912 16244
rect 3148 16056 3200 16108
rect 52552 16099 52604 16108
rect 52552 16065 52561 16099
rect 52561 16065 52595 16099
rect 52595 16065 52604 16099
rect 52552 16056 52604 16065
rect 53012 16056 53064 16108
rect 53932 16056 53984 16108
rect 57244 16192 57296 16244
rect 3056 15988 3108 16040
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 50804 15988 50856 16040
rect 51264 15988 51316 16040
rect 51632 15988 51684 16040
rect 52000 15988 52052 16040
rect 53288 15988 53340 16040
rect 54852 15988 54904 16040
rect 55680 15988 55732 16040
rect 51356 15920 51408 15972
rect 53012 15920 53064 15972
rect 3240 15895 3292 15904
rect 3240 15861 3249 15895
rect 3249 15861 3283 15895
rect 3283 15861 3292 15895
rect 3240 15852 3292 15861
rect 49976 15852 50028 15904
rect 52552 15852 52604 15904
rect 52644 15852 52696 15904
rect 54484 15852 54536 15904
rect 55496 15852 55548 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 50326 15750 50378 15802
rect 50390 15750 50442 15802
rect 50454 15750 50506 15802
rect 50518 15750 50570 15802
rect 1860 15555 1912 15564
rect 1860 15521 1869 15555
rect 1869 15521 1903 15555
rect 1903 15521 1912 15555
rect 1860 15512 1912 15521
rect 2596 15555 2648 15564
rect 2596 15521 2605 15555
rect 2605 15521 2639 15555
rect 2639 15521 2648 15555
rect 2596 15512 2648 15521
rect 49700 15555 49752 15564
rect 49700 15521 49709 15555
rect 49709 15521 49743 15555
rect 49743 15521 49752 15555
rect 49700 15512 49752 15521
rect 51172 15648 51224 15700
rect 52644 15648 52696 15700
rect 53012 15648 53064 15700
rect 53288 15648 53340 15700
rect 55128 15648 55180 15700
rect 55956 15648 56008 15700
rect 56324 15648 56376 15700
rect 51908 15623 51960 15632
rect 50712 15512 50764 15564
rect 51908 15589 51917 15623
rect 51917 15589 51951 15623
rect 51951 15589 51960 15623
rect 51908 15580 51960 15589
rect 53840 15580 53892 15632
rect 52000 15555 52052 15564
rect 52000 15521 52009 15555
rect 52009 15521 52043 15555
rect 52043 15521 52052 15555
rect 52000 15512 52052 15521
rect 53012 15512 53064 15564
rect 2780 15419 2832 15428
rect 2780 15385 2789 15419
rect 2789 15385 2823 15419
rect 2823 15385 2832 15419
rect 2780 15376 2832 15385
rect 53288 15555 53340 15564
rect 53288 15521 53297 15555
rect 53297 15521 53331 15555
rect 53331 15521 53340 15555
rect 53288 15512 53340 15521
rect 53472 15555 53524 15564
rect 53472 15521 53481 15555
rect 53481 15521 53515 15555
rect 53515 15521 53524 15555
rect 53472 15512 53524 15521
rect 54484 15512 54536 15564
rect 55220 15512 55272 15564
rect 55680 15512 55732 15564
rect 56600 15512 56652 15564
rect 57980 15555 58032 15564
rect 57980 15521 57989 15555
rect 57989 15521 58023 15555
rect 58023 15521 58032 15555
rect 57980 15512 58032 15521
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 51264 15308 51316 15360
rect 53196 15308 53248 15360
rect 54024 15351 54076 15360
rect 54024 15317 54033 15351
rect 54033 15317 54067 15351
rect 54067 15317 54076 15351
rect 54024 15308 54076 15317
rect 54668 15308 54720 15360
rect 55772 15308 55824 15360
rect 57888 15308 57940 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 2596 15104 2648 15156
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 4068 15036 4120 15088
rect 3240 14968 3292 15020
rect 49792 14968 49844 15020
rect 51908 15104 51960 15156
rect 52460 15104 52512 15156
rect 53472 15104 53524 15156
rect 54576 15147 54628 15156
rect 54576 15113 54585 15147
rect 54585 15113 54619 15147
rect 54619 15113 54628 15147
rect 54576 15104 54628 15113
rect 57980 15147 58032 15156
rect 52000 15036 52052 15088
rect 57980 15113 57989 15147
rect 57989 15113 58023 15147
rect 58023 15113 58032 15147
rect 57980 15104 58032 15113
rect 2964 14900 3016 14952
rect 52460 14943 52512 14952
rect 52460 14909 52469 14943
rect 52469 14909 52503 14943
rect 52503 14909 52512 14943
rect 52460 14900 52512 14909
rect 52552 14900 52604 14952
rect 52736 14943 52788 14952
rect 52736 14909 52745 14943
rect 52745 14909 52779 14943
rect 52779 14909 52788 14943
rect 52736 14900 52788 14909
rect 54024 14900 54076 14952
rect 54300 14943 54352 14952
rect 54300 14909 54309 14943
rect 54309 14909 54343 14943
rect 54343 14909 54352 14943
rect 54300 14900 54352 14909
rect 51448 14832 51500 14884
rect 54116 14764 54168 14816
rect 54944 14900 54996 14952
rect 54760 14832 54812 14884
rect 55312 14832 55364 14884
rect 55220 14764 55272 14816
rect 55588 14764 55640 14816
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 50326 14662 50378 14714
rect 50390 14662 50442 14714
rect 50454 14662 50506 14714
rect 50518 14662 50570 14714
rect 1860 14560 1912 14612
rect 54024 14560 54076 14612
rect 54208 14603 54260 14612
rect 54208 14569 54217 14603
rect 54217 14569 54251 14603
rect 54251 14569 54260 14603
rect 54208 14560 54260 14569
rect 54300 14560 54352 14612
rect 54576 14560 54628 14612
rect 55588 14560 55640 14612
rect 2504 14356 2556 14408
rect 49976 14424 50028 14476
rect 51264 14424 51316 14476
rect 52368 14467 52420 14476
rect 50252 14356 50304 14408
rect 51356 14356 51408 14408
rect 52368 14433 52377 14467
rect 52377 14433 52411 14467
rect 52411 14433 52420 14467
rect 52368 14424 52420 14433
rect 52644 14467 52696 14476
rect 52644 14433 52678 14467
rect 52678 14433 52696 14467
rect 54392 14467 54444 14476
rect 52644 14424 52696 14433
rect 54392 14433 54401 14467
rect 54401 14433 54435 14467
rect 54435 14433 54444 14467
rect 54392 14424 54444 14433
rect 54484 14467 54536 14476
rect 54484 14433 54493 14467
rect 54493 14433 54527 14467
rect 54527 14433 54536 14467
rect 54484 14424 54536 14433
rect 54668 14424 54720 14476
rect 55220 14424 55272 14476
rect 55588 14424 55640 14476
rect 55772 14467 55824 14476
rect 55772 14433 55781 14467
rect 55781 14433 55815 14467
rect 55815 14433 55824 14467
rect 55772 14424 55824 14433
rect 55956 14424 56008 14476
rect 3976 14288 4028 14340
rect 51448 14331 51500 14340
rect 51448 14297 51457 14331
rect 51457 14297 51491 14331
rect 51491 14297 51500 14331
rect 51448 14288 51500 14297
rect 54484 14288 54536 14340
rect 54024 14220 54076 14272
rect 54668 14263 54720 14272
rect 54668 14229 54677 14263
rect 54677 14229 54711 14263
rect 54711 14229 54720 14263
rect 54668 14220 54720 14229
rect 55128 14220 55180 14272
rect 55772 14220 55824 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 2504 14059 2556 14068
rect 2504 14025 2513 14059
rect 2513 14025 2547 14059
rect 2547 14025 2556 14059
rect 2504 14016 2556 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 49700 14016 49752 14068
rect 50988 14016 51040 14068
rect 52000 14016 52052 14068
rect 52644 14016 52696 14068
rect 53932 14016 53984 14068
rect 54668 14016 54720 14068
rect 54760 13991 54812 14000
rect 54760 13957 54769 13991
rect 54769 13957 54803 13991
rect 54803 13957 54812 13991
rect 55496 13991 55548 14000
rect 54760 13948 54812 13957
rect 55496 13957 55505 13991
rect 55505 13957 55539 13991
rect 55539 13957 55548 13991
rect 55496 13948 55548 13957
rect 3056 13812 3108 13864
rect 49148 13855 49200 13864
rect 49148 13821 49157 13855
rect 49157 13821 49191 13855
rect 49191 13821 49200 13855
rect 49148 13812 49200 13821
rect 50436 13855 50488 13864
rect 50436 13821 50445 13855
rect 50445 13821 50479 13855
rect 50479 13821 50488 13855
rect 50436 13812 50488 13821
rect 2044 13744 2096 13796
rect 49424 13744 49476 13796
rect 50252 13744 50304 13796
rect 50712 13812 50764 13864
rect 52920 13880 52972 13932
rect 55680 13880 55732 13932
rect 51264 13812 51316 13864
rect 51540 13812 51592 13864
rect 52092 13855 52144 13864
rect 51632 13744 51684 13796
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 3148 13719 3200 13728
rect 3148 13685 3157 13719
rect 3157 13685 3191 13719
rect 3191 13685 3200 13719
rect 3148 13676 3200 13685
rect 51080 13676 51132 13728
rect 52092 13821 52101 13855
rect 52101 13821 52135 13855
rect 52135 13821 52144 13855
rect 52092 13812 52144 13821
rect 52552 13855 52604 13864
rect 52552 13821 52561 13855
rect 52561 13821 52595 13855
rect 52595 13821 52604 13855
rect 52736 13855 52788 13864
rect 52552 13812 52604 13821
rect 52736 13821 52745 13855
rect 52745 13821 52779 13855
rect 52779 13821 52788 13855
rect 52736 13812 52788 13821
rect 54300 13812 54352 13864
rect 54392 13855 54444 13864
rect 54392 13821 54401 13855
rect 54401 13821 54435 13855
rect 54435 13821 54444 13855
rect 54392 13812 54444 13821
rect 54116 13744 54168 13796
rect 55772 13812 55824 13864
rect 56048 13855 56100 13864
rect 56048 13821 56057 13855
rect 56057 13821 56091 13855
rect 56091 13821 56100 13855
rect 56048 13812 56100 13821
rect 57060 13855 57112 13864
rect 57060 13821 57069 13855
rect 57069 13821 57103 13855
rect 57103 13821 57112 13855
rect 57060 13812 57112 13821
rect 57520 13855 57572 13864
rect 57520 13821 57529 13855
rect 57529 13821 57563 13855
rect 57563 13821 57572 13855
rect 57520 13812 57572 13821
rect 57704 13855 57756 13864
rect 57704 13821 57713 13855
rect 57713 13821 57747 13855
rect 57747 13821 57756 13855
rect 57704 13812 57756 13821
rect 52552 13676 52604 13728
rect 54576 13676 54628 13728
rect 56140 13719 56192 13728
rect 56140 13685 56149 13719
rect 56149 13685 56183 13719
rect 56183 13685 56192 13719
rect 56140 13676 56192 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 50326 13574 50378 13626
rect 50390 13574 50442 13626
rect 50454 13574 50506 13626
rect 50518 13574 50570 13626
rect 55312 13515 55364 13524
rect 51080 13404 51132 13456
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 3148 13268 3200 13320
rect 2044 13243 2096 13252
rect 2044 13209 2053 13243
rect 2053 13209 2087 13243
rect 2087 13209 2096 13243
rect 2044 13200 2096 13209
rect 5080 13175 5132 13184
rect 5080 13141 5089 13175
rect 5089 13141 5123 13175
rect 5123 13141 5132 13175
rect 47492 13336 47544 13388
rect 49884 13379 49936 13388
rect 49884 13345 49893 13379
rect 49893 13345 49927 13379
rect 49927 13345 49936 13379
rect 49884 13336 49936 13345
rect 51356 13336 51408 13388
rect 50436 13311 50488 13320
rect 50436 13277 50445 13311
rect 50445 13277 50479 13311
rect 50479 13277 50488 13311
rect 51448 13311 51500 13320
rect 50436 13268 50488 13277
rect 51448 13277 51457 13311
rect 51457 13277 51491 13311
rect 51491 13277 51500 13311
rect 51448 13268 51500 13277
rect 53932 13447 53984 13456
rect 53932 13413 53941 13447
rect 53941 13413 53975 13447
rect 53975 13413 53984 13447
rect 53932 13404 53984 13413
rect 54024 13404 54076 13456
rect 55312 13481 55321 13515
rect 55321 13481 55355 13515
rect 55355 13481 55364 13515
rect 55312 13472 55364 13481
rect 53196 13336 53248 13388
rect 54392 13336 54444 13388
rect 54576 13379 54628 13388
rect 54576 13345 54585 13379
rect 54585 13345 54619 13379
rect 54619 13345 54628 13379
rect 54576 13336 54628 13345
rect 55220 13379 55272 13388
rect 55220 13345 55229 13379
rect 55229 13345 55263 13379
rect 55263 13345 55272 13379
rect 55220 13336 55272 13345
rect 55956 13336 56008 13388
rect 52000 13311 52052 13320
rect 52000 13277 52009 13311
rect 52009 13277 52043 13311
rect 52043 13277 52052 13311
rect 52000 13268 52052 13277
rect 54300 13268 54352 13320
rect 55772 13268 55824 13320
rect 5080 13132 5132 13141
rect 47584 13132 47636 13184
rect 52920 13132 52972 13184
rect 53104 13132 53156 13184
rect 57244 13132 57296 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 50988 12928 51040 12980
rect 51448 12928 51500 12980
rect 52000 12928 52052 12980
rect 54208 12928 54260 12980
rect 55220 12928 55272 12980
rect 57336 12971 57388 12980
rect 57336 12937 57345 12971
rect 57345 12937 57379 12971
rect 57379 12937 57388 12971
rect 57336 12928 57388 12937
rect 51264 12792 51316 12844
rect 5080 12724 5132 12776
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 50436 12724 50488 12776
rect 51724 12724 51776 12776
rect 51816 12724 51868 12776
rect 52828 12767 52880 12776
rect 52828 12733 52837 12767
rect 52837 12733 52871 12767
rect 52871 12733 52880 12767
rect 54300 12792 54352 12844
rect 54944 12792 54996 12844
rect 52828 12724 52880 12733
rect 53104 12767 53156 12776
rect 53104 12733 53113 12767
rect 53113 12733 53147 12767
rect 53147 12733 53156 12767
rect 53104 12724 53156 12733
rect 53932 12724 53984 12776
rect 54208 12767 54260 12776
rect 54208 12733 54217 12767
rect 54217 12733 54251 12767
rect 54251 12733 54260 12767
rect 54208 12724 54260 12733
rect 57520 12792 57572 12844
rect 57244 12767 57296 12776
rect 57244 12733 57253 12767
rect 57253 12733 57287 12767
rect 57287 12733 57296 12767
rect 57244 12724 57296 12733
rect 55588 12656 55640 12708
rect 57980 12699 58032 12708
rect 57980 12665 57989 12699
rect 57989 12665 58023 12699
rect 58023 12665 58032 12699
rect 57980 12656 58032 12665
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 51172 12631 51224 12640
rect 51172 12597 51181 12631
rect 51181 12597 51215 12631
rect 51215 12597 51224 12631
rect 51172 12588 51224 12597
rect 51816 12588 51868 12640
rect 52460 12588 52512 12640
rect 52644 12588 52696 12640
rect 53104 12588 53156 12640
rect 53564 12588 53616 12640
rect 53656 12588 53708 12640
rect 54852 12588 54904 12640
rect 56692 12588 56744 12640
rect 57888 12588 57940 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 50326 12486 50378 12538
rect 50390 12486 50442 12538
rect 50454 12486 50506 12538
rect 50518 12486 50570 12538
rect 52000 12384 52052 12436
rect 52368 12384 52420 12436
rect 1768 12223 1820 12232
rect 1768 12189 1777 12223
rect 1777 12189 1811 12223
rect 1811 12189 1820 12223
rect 1768 12180 1820 12189
rect 2964 12248 3016 12300
rect 49884 12291 49936 12300
rect 49884 12257 49893 12291
rect 49893 12257 49927 12291
rect 49927 12257 49936 12291
rect 49884 12248 49936 12257
rect 50528 12291 50580 12300
rect 50528 12257 50537 12291
rect 50537 12257 50571 12291
rect 50571 12257 50580 12291
rect 50528 12248 50580 12257
rect 51172 12248 51224 12300
rect 51724 12291 51776 12300
rect 51724 12257 51733 12291
rect 51733 12257 51767 12291
rect 51767 12257 51776 12291
rect 52000 12291 52052 12300
rect 51724 12248 51776 12257
rect 52000 12257 52009 12291
rect 52009 12257 52043 12291
rect 52043 12257 52052 12291
rect 52000 12248 52052 12257
rect 50896 12180 50948 12232
rect 51080 12180 51132 12232
rect 51816 12180 51868 12232
rect 54300 12384 54352 12436
rect 55128 12384 55180 12436
rect 57980 12384 58032 12436
rect 52276 12248 52328 12300
rect 52920 12291 52972 12300
rect 52920 12257 52929 12291
rect 52929 12257 52963 12291
rect 52963 12257 52972 12291
rect 52920 12248 52972 12257
rect 53012 12291 53064 12300
rect 53012 12257 53021 12291
rect 53021 12257 53055 12291
rect 53055 12257 53064 12291
rect 53012 12248 53064 12257
rect 53196 12291 53248 12300
rect 53196 12257 53205 12291
rect 53205 12257 53239 12291
rect 53239 12257 53248 12291
rect 53196 12248 53248 12257
rect 54208 12248 54260 12300
rect 54944 12248 54996 12300
rect 56692 12291 56744 12300
rect 1860 12112 1912 12164
rect 53472 12112 53524 12164
rect 54760 12112 54812 12164
rect 56692 12257 56701 12291
rect 56701 12257 56735 12291
rect 56735 12257 56744 12291
rect 56692 12248 56744 12257
rect 57612 12180 57664 12232
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 49884 12044 49936 12096
rect 50804 12044 50856 12096
rect 50896 12044 50948 12096
rect 52920 12044 52972 12096
rect 54576 12044 54628 12096
rect 55404 12044 55456 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 1768 11840 1820 11892
rect 2872 11636 2924 11688
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 51080 11840 51132 11892
rect 51724 11840 51776 11892
rect 52000 11840 52052 11892
rect 52828 11840 52880 11892
rect 53564 11840 53616 11892
rect 55404 11840 55456 11892
rect 55588 11883 55640 11892
rect 55588 11849 55597 11883
rect 55597 11849 55631 11883
rect 55631 11849 55640 11883
rect 55588 11840 55640 11849
rect 53932 11772 53984 11824
rect 56692 11815 56744 11824
rect 56692 11781 56701 11815
rect 56701 11781 56735 11815
rect 56735 11781 56744 11815
rect 56692 11772 56744 11781
rect 53472 11704 53524 11756
rect 49424 11679 49476 11688
rect 49424 11645 49433 11679
rect 49433 11645 49467 11679
rect 49467 11645 49476 11679
rect 49424 11636 49476 11645
rect 49792 11636 49844 11688
rect 1860 11611 1912 11620
rect 1860 11577 1869 11611
rect 1869 11577 1903 11611
rect 1903 11577 1912 11611
rect 1860 11568 1912 11577
rect 2596 11611 2648 11620
rect 2596 11577 2605 11611
rect 2605 11577 2639 11611
rect 2639 11577 2648 11611
rect 2596 11568 2648 11577
rect 2780 11611 2832 11620
rect 2780 11577 2789 11611
rect 2789 11577 2823 11611
rect 2823 11577 2832 11611
rect 2780 11568 2832 11577
rect 49332 11611 49384 11620
rect 49332 11577 49341 11611
rect 49341 11577 49375 11611
rect 49375 11577 49384 11611
rect 49332 11568 49384 11577
rect 50620 11636 50672 11688
rect 51172 11636 51224 11688
rect 51540 11568 51592 11620
rect 52828 11636 52880 11688
rect 54760 11679 54812 11688
rect 54760 11645 54769 11679
rect 54769 11645 54803 11679
rect 54803 11645 54812 11679
rect 54760 11636 54812 11645
rect 54852 11679 54904 11688
rect 54852 11645 54861 11679
rect 54861 11645 54895 11679
rect 54895 11645 54904 11679
rect 55128 11679 55180 11688
rect 54852 11636 54904 11645
rect 55128 11645 55137 11679
rect 55137 11645 55171 11679
rect 55171 11645 55180 11679
rect 55128 11636 55180 11645
rect 55588 11679 55640 11688
rect 55588 11645 55597 11679
rect 55597 11645 55631 11679
rect 55631 11645 55640 11679
rect 55588 11636 55640 11645
rect 54668 11568 54720 11620
rect 56324 11636 56376 11688
rect 57152 11679 57204 11688
rect 57152 11645 57161 11679
rect 57161 11645 57195 11679
rect 57195 11645 57204 11679
rect 57152 11636 57204 11645
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 52460 11500 52512 11552
rect 52552 11500 52604 11552
rect 53012 11500 53064 11552
rect 57980 11500 58032 11552
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 50326 11398 50378 11450
rect 50390 11398 50442 11450
rect 50454 11398 50506 11450
rect 50518 11398 50570 11450
rect 2596 11296 2648 11348
rect 50712 11296 50764 11348
rect 51540 11339 51592 11348
rect 51540 11305 51549 11339
rect 51549 11305 51583 11339
rect 51583 11305 51592 11339
rect 51540 11296 51592 11305
rect 52736 11296 52788 11348
rect 53012 11296 53064 11348
rect 4068 11228 4120 11280
rect 2872 11160 2924 11212
rect 52368 11228 52420 11280
rect 52552 11228 52604 11280
rect 50620 11160 50672 11212
rect 51448 11203 51500 11212
rect 51448 11169 51457 11203
rect 51457 11169 51491 11203
rect 51491 11169 51500 11203
rect 51448 11160 51500 11169
rect 52000 11160 52052 11212
rect 52828 11160 52880 11212
rect 53012 11203 53064 11212
rect 53012 11169 53021 11203
rect 53021 11169 53055 11203
rect 53055 11169 53064 11203
rect 53012 11160 53064 11169
rect 53656 11228 53708 11280
rect 54208 11228 54260 11280
rect 52644 11092 52696 11144
rect 53196 11135 53248 11144
rect 53196 11101 53205 11135
rect 53205 11101 53239 11135
rect 53239 11101 53248 11135
rect 56692 11296 56744 11348
rect 54668 11271 54720 11280
rect 54668 11237 54677 11271
rect 54677 11237 54711 11271
rect 54711 11237 54720 11271
rect 54668 11228 54720 11237
rect 55588 11228 55640 11280
rect 57980 11271 58032 11280
rect 54576 11203 54628 11212
rect 54576 11169 54585 11203
rect 54585 11169 54619 11203
rect 54619 11169 54628 11203
rect 54576 11160 54628 11169
rect 55496 11203 55548 11212
rect 55496 11169 55505 11203
rect 55505 11169 55539 11203
rect 55539 11169 55548 11203
rect 55496 11160 55548 11169
rect 55680 11203 55732 11212
rect 55680 11169 55689 11203
rect 55689 11169 55723 11203
rect 55723 11169 55732 11203
rect 55680 11160 55732 11169
rect 57980 11237 57989 11271
rect 57989 11237 58023 11271
rect 58023 11237 58032 11271
rect 57980 11228 58032 11237
rect 58164 11271 58216 11280
rect 58164 11237 58173 11271
rect 58173 11237 58207 11271
rect 58207 11237 58216 11271
rect 58164 11228 58216 11237
rect 53196 11092 53248 11101
rect 52092 11024 52144 11076
rect 55588 11092 55640 11144
rect 55772 11092 55824 11144
rect 54668 11024 54720 11076
rect 55220 10956 55272 11008
rect 56692 10999 56744 11008
rect 56692 10965 56701 10999
rect 56701 10965 56735 10999
rect 56735 10965 56744 10999
rect 56692 10956 56744 10965
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 1860 10752 1912 10804
rect 54024 10752 54076 10804
rect 54944 10752 54996 10804
rect 55680 10752 55732 10804
rect 53104 10684 53156 10736
rect 53840 10684 53892 10736
rect 54300 10684 54352 10736
rect 54392 10616 54444 10668
rect 2504 10548 2556 10600
rect 50804 10591 50856 10600
rect 50804 10557 50813 10591
rect 50813 10557 50847 10591
rect 50847 10557 50856 10591
rect 50804 10548 50856 10557
rect 51908 10548 51960 10600
rect 52092 10548 52144 10600
rect 54760 10616 54812 10668
rect 3332 10480 3384 10532
rect 54668 10523 54720 10532
rect 54668 10489 54677 10523
rect 54677 10489 54711 10523
rect 54711 10489 54720 10523
rect 54668 10480 54720 10489
rect 51264 10455 51316 10464
rect 51264 10421 51273 10455
rect 51273 10421 51307 10455
rect 51307 10421 51316 10455
rect 51264 10412 51316 10421
rect 52920 10412 52972 10464
rect 53196 10412 53248 10464
rect 54484 10412 54536 10464
rect 54576 10412 54628 10464
rect 54944 10548 54996 10600
rect 56692 10548 56744 10600
rect 57520 10480 57572 10532
rect 57980 10523 58032 10532
rect 57980 10489 57989 10523
rect 57989 10489 58023 10523
rect 58023 10489 58032 10523
rect 57980 10480 58032 10489
rect 58164 10523 58216 10532
rect 58164 10489 58173 10523
rect 58173 10489 58207 10523
rect 58207 10489 58216 10523
rect 58164 10480 58216 10489
rect 55680 10412 55732 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 50326 10310 50378 10362
rect 50390 10310 50442 10362
rect 50454 10310 50506 10362
rect 50518 10310 50570 10362
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 50804 10208 50856 10260
rect 54300 10208 54352 10260
rect 54392 10208 54444 10260
rect 57980 10208 58032 10260
rect 50068 10140 50120 10192
rect 51264 10140 51316 10192
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 2872 10072 2924 10124
rect 3332 10115 3384 10124
rect 3332 10081 3341 10115
rect 3341 10081 3375 10115
rect 3375 10081 3384 10115
rect 3332 10072 3384 10081
rect 49976 10115 50028 10124
rect 49976 10081 49985 10115
rect 49985 10081 50019 10115
rect 50019 10081 50028 10115
rect 49976 10072 50028 10081
rect 51172 10072 51224 10124
rect 52460 10072 52512 10124
rect 50160 10004 50212 10056
rect 50988 10004 51040 10056
rect 53840 10072 53892 10124
rect 53932 10115 53984 10124
rect 53932 10081 53941 10115
rect 53941 10081 53975 10115
rect 53975 10081 53984 10115
rect 54576 10115 54628 10124
rect 53932 10072 53984 10081
rect 54576 10081 54585 10115
rect 54585 10081 54619 10115
rect 54619 10081 54628 10115
rect 54576 10072 54628 10081
rect 55220 10115 55272 10124
rect 55220 10081 55229 10115
rect 55229 10081 55263 10115
rect 55263 10081 55272 10115
rect 55220 10072 55272 10081
rect 54484 10004 54536 10056
rect 55496 10115 55548 10124
rect 55496 10081 55505 10115
rect 55505 10081 55539 10115
rect 55539 10081 55548 10115
rect 55496 10072 55548 10081
rect 55680 10072 55732 10124
rect 56876 10115 56928 10124
rect 56876 10081 56885 10115
rect 56885 10081 56919 10115
rect 56919 10081 56928 10115
rect 56876 10072 56928 10081
rect 55772 10004 55824 10056
rect 55496 9936 55548 9988
rect 57060 9979 57112 9988
rect 57060 9945 57069 9979
rect 57069 9945 57103 9979
rect 57103 9945 57112 9979
rect 57060 9936 57112 9945
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 50344 9911 50396 9920
rect 50344 9877 50353 9911
rect 50353 9877 50387 9911
rect 50387 9877 50396 9911
rect 50344 9868 50396 9877
rect 54116 9868 54168 9920
rect 54208 9868 54260 9920
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 1860 9664 1912 9716
rect 51172 9707 51224 9716
rect 51172 9673 51181 9707
rect 51181 9673 51215 9707
rect 51215 9673 51224 9707
rect 51172 9664 51224 9673
rect 50712 9596 50764 9648
rect 56876 9664 56928 9716
rect 50160 9528 50212 9580
rect 2872 9460 2924 9512
rect 48872 9392 48924 9444
rect 50344 9460 50396 9512
rect 51356 9503 51408 9512
rect 50988 9392 51040 9444
rect 51356 9469 51365 9503
rect 51365 9469 51399 9503
rect 51399 9469 51408 9503
rect 51356 9460 51408 9469
rect 51816 9460 51868 9512
rect 52460 9503 52512 9512
rect 52460 9469 52469 9503
rect 52469 9469 52503 9503
rect 52503 9469 52512 9503
rect 52460 9460 52512 9469
rect 53840 9460 53892 9512
rect 54024 9503 54076 9512
rect 54024 9469 54033 9503
rect 54033 9469 54067 9503
rect 54067 9469 54076 9503
rect 54024 9460 54076 9469
rect 54116 9460 54168 9512
rect 55588 9460 55640 9512
rect 56968 9503 57020 9512
rect 56968 9469 56977 9503
rect 56977 9469 57011 9503
rect 57011 9469 57020 9503
rect 56968 9460 57020 9469
rect 50160 9324 50212 9376
rect 55220 9392 55272 9444
rect 55312 9392 55364 9444
rect 57980 9435 58032 9444
rect 57980 9401 57989 9435
rect 57989 9401 58023 9435
rect 58023 9401 58032 9435
rect 57980 9392 58032 9401
rect 58164 9435 58216 9444
rect 58164 9401 58173 9435
rect 58173 9401 58207 9435
rect 58207 9401 58216 9435
rect 58164 9392 58216 9401
rect 52460 9324 52512 9376
rect 54208 9324 54260 9376
rect 54668 9324 54720 9376
rect 55956 9367 56008 9376
rect 55956 9333 55965 9367
rect 55965 9333 55999 9367
rect 55999 9333 56008 9367
rect 55956 9324 56008 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 50326 9222 50378 9274
rect 50390 9222 50442 9274
rect 50454 9222 50506 9274
rect 50518 9222 50570 9274
rect 49976 9163 50028 9172
rect 49976 9129 49985 9163
rect 49985 9129 50019 9163
rect 50019 9129 50028 9163
rect 49976 9120 50028 9129
rect 50712 9120 50764 9172
rect 52000 9120 52052 9172
rect 53932 9120 53984 9172
rect 54484 9163 54536 9172
rect 54484 9129 54493 9163
rect 54493 9129 54527 9163
rect 54527 9129 54536 9163
rect 54484 9120 54536 9129
rect 57704 9120 57756 9172
rect 57980 9120 58032 9172
rect 2872 8984 2924 9036
rect 48044 9027 48096 9036
rect 48044 8993 48053 9027
rect 48053 8993 48087 9027
rect 48087 8993 48096 9027
rect 48044 8984 48096 8993
rect 50896 9052 50948 9104
rect 51632 9052 51684 9104
rect 52920 9095 52972 9104
rect 52920 9061 52929 9095
rect 52929 9061 52963 9095
rect 52963 9061 52972 9095
rect 52920 9052 52972 9061
rect 53012 9052 53064 9104
rect 49516 9027 49568 9036
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 49516 8993 49525 9027
rect 49525 8993 49559 9027
rect 49559 8993 49568 9027
rect 49516 8984 49568 8993
rect 50160 9027 50212 9036
rect 50160 8993 50169 9027
rect 50169 8993 50203 9027
rect 50203 8993 50212 9027
rect 50160 8984 50212 8993
rect 50252 9027 50304 9036
rect 50252 8993 50261 9027
rect 50261 8993 50295 9027
rect 50295 8993 50304 9027
rect 50252 8984 50304 8993
rect 50804 8984 50856 9036
rect 49608 8916 49660 8968
rect 51448 8916 51500 8968
rect 52368 8984 52420 9036
rect 54392 9052 54444 9104
rect 54668 9027 54720 9036
rect 52828 8916 52880 8968
rect 54668 8993 54677 9027
rect 54677 8993 54711 9027
rect 54711 8993 54720 9027
rect 54668 8984 54720 8993
rect 54760 9027 54812 9036
rect 54760 8993 54769 9027
rect 54769 8993 54803 9027
rect 54803 8993 54812 9027
rect 54760 8984 54812 8993
rect 56784 8984 56836 9036
rect 57520 9027 57572 9036
rect 57520 8993 57529 9027
rect 57529 8993 57563 9027
rect 57563 8993 57572 9027
rect 57520 8984 57572 8993
rect 57704 8959 57756 8968
rect 57704 8925 57713 8959
rect 57713 8925 57747 8959
rect 57747 8925 57756 8959
rect 57704 8916 57756 8925
rect 56968 8848 57020 8900
rect 2596 8780 2648 8832
rect 48688 8823 48740 8832
rect 48688 8789 48697 8823
rect 48697 8789 48731 8823
rect 48731 8789 48740 8823
rect 48688 8780 48740 8789
rect 49884 8780 49936 8832
rect 54116 8780 54168 8832
rect 54944 8823 54996 8832
rect 54944 8789 54953 8823
rect 54953 8789 54987 8823
rect 54987 8789 54996 8823
rect 54944 8780 54996 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 1676 8576 1728 8628
rect 2780 8551 2832 8560
rect 2780 8517 2789 8551
rect 2789 8517 2823 8551
rect 2823 8517 2832 8551
rect 2780 8508 2832 8517
rect 3700 8508 3752 8560
rect 50252 8551 50304 8560
rect 50252 8517 50261 8551
rect 50261 8517 50295 8551
rect 50295 8517 50304 8551
rect 51448 8551 51500 8560
rect 50252 8508 50304 8517
rect 48872 8483 48924 8492
rect 2596 8415 2648 8424
rect 2596 8381 2605 8415
rect 2605 8381 2639 8415
rect 2639 8381 2648 8415
rect 2596 8372 2648 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 2044 8347 2096 8356
rect 2044 8313 2053 8347
rect 2053 8313 2087 8347
rect 2087 8313 2096 8347
rect 2044 8304 2096 8313
rect 48872 8449 48881 8483
rect 48881 8449 48915 8483
rect 48915 8449 48924 8483
rect 48872 8440 48924 8449
rect 50160 8440 50212 8492
rect 51448 8517 51457 8551
rect 51457 8517 51491 8551
rect 51491 8517 51500 8551
rect 51448 8508 51500 8517
rect 47032 8415 47084 8424
rect 47032 8381 47041 8415
rect 47041 8381 47075 8415
rect 47075 8381 47084 8415
rect 47032 8372 47084 8381
rect 47584 8304 47636 8356
rect 47768 8372 47820 8424
rect 50068 8304 50120 8356
rect 51816 8440 51868 8492
rect 51908 8372 51960 8424
rect 52460 8508 52512 8560
rect 53932 8440 53984 8492
rect 52828 8415 52880 8424
rect 52828 8381 52837 8415
rect 52837 8381 52871 8415
rect 52871 8381 52880 8415
rect 52828 8372 52880 8381
rect 52920 8415 52972 8424
rect 52920 8381 52929 8415
rect 52929 8381 52963 8415
rect 52963 8381 52972 8415
rect 52920 8372 52972 8381
rect 53840 8372 53892 8424
rect 54116 8372 54168 8424
rect 54760 8372 54812 8424
rect 55128 8372 55180 8424
rect 56600 8415 56652 8424
rect 56600 8381 56609 8415
rect 56609 8381 56643 8415
rect 56643 8381 56652 8415
rect 56600 8372 56652 8381
rect 46940 8236 46992 8288
rect 50620 8236 50672 8288
rect 50804 8279 50856 8288
rect 50804 8245 50813 8279
rect 50813 8245 50847 8279
rect 50847 8245 50856 8279
rect 50804 8236 50856 8245
rect 51264 8236 51316 8288
rect 52092 8279 52144 8288
rect 52092 8245 52101 8279
rect 52101 8245 52135 8279
rect 52135 8245 52144 8279
rect 52092 8236 52144 8245
rect 55956 8304 56008 8356
rect 58164 8347 58216 8356
rect 58164 8313 58173 8347
rect 58173 8313 58207 8347
rect 58207 8313 58216 8347
rect 58164 8304 58216 8313
rect 57428 8236 57480 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 50326 8134 50378 8186
rect 50390 8134 50442 8186
rect 50454 8134 50506 8186
rect 50518 8134 50570 8186
rect 49332 8075 49384 8084
rect 49332 8041 49341 8075
rect 49341 8041 49375 8075
rect 49375 8041 49384 8075
rect 49332 8032 49384 8041
rect 50068 8075 50120 8084
rect 50068 8041 50077 8075
rect 50077 8041 50111 8075
rect 50111 8041 50120 8075
rect 50068 8032 50120 8041
rect 2320 7896 2372 7948
rect 3148 7964 3200 8016
rect 47032 7964 47084 8016
rect 55220 8032 55272 8084
rect 57612 8032 57664 8084
rect 50620 7964 50672 8016
rect 51264 7964 51316 8016
rect 51356 7964 51408 8016
rect 2780 7896 2832 7948
rect 46940 7939 46992 7948
rect 46940 7905 46949 7939
rect 46949 7905 46983 7939
rect 46983 7905 46992 7939
rect 46940 7896 46992 7905
rect 47768 7896 47820 7948
rect 47952 7896 48004 7948
rect 48412 7896 48464 7948
rect 48964 7896 49016 7948
rect 49516 7939 49568 7948
rect 49516 7905 49525 7939
rect 49525 7905 49559 7939
rect 49559 7905 49568 7939
rect 49516 7896 49568 7905
rect 49884 7896 49936 7948
rect 50804 7896 50856 7948
rect 50988 7896 51040 7948
rect 52092 7964 52144 8016
rect 54944 7964 54996 8016
rect 52920 7896 52972 7948
rect 53196 7896 53248 7948
rect 51540 7828 51592 7880
rect 54760 7896 54812 7948
rect 55128 7939 55180 7948
rect 55128 7905 55137 7939
rect 55137 7905 55171 7939
rect 55171 7905 55180 7939
rect 55128 7896 55180 7905
rect 56784 7896 56836 7948
rect 56968 7828 57020 7880
rect 57336 7871 57388 7880
rect 57336 7837 57345 7871
rect 57345 7837 57379 7871
rect 57379 7837 57388 7871
rect 57336 7828 57388 7837
rect 1952 7735 2004 7744
rect 1952 7701 1961 7735
rect 1961 7701 1995 7735
rect 1995 7701 2004 7735
rect 1952 7692 2004 7701
rect 2780 7692 2832 7744
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 47768 7692 47820 7744
rect 51356 7692 51408 7744
rect 53472 7735 53524 7744
rect 53472 7701 53481 7735
rect 53481 7701 53515 7735
rect 53515 7701 53524 7735
rect 53472 7692 53524 7701
rect 53564 7735 53616 7744
rect 53564 7701 53573 7735
rect 53573 7701 53607 7735
rect 53607 7701 53616 7735
rect 53564 7692 53616 7701
rect 54760 7692 54812 7744
rect 55496 7692 55548 7744
rect 55864 7692 55916 7744
rect 56876 7692 56928 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 1860 7488 1912 7540
rect 47584 7488 47636 7540
rect 47952 7488 48004 7540
rect 49700 7488 49752 7540
rect 51448 7531 51500 7540
rect 49608 7420 49660 7472
rect 51448 7497 51457 7531
rect 51457 7497 51491 7531
rect 51491 7497 51500 7531
rect 51448 7488 51500 7497
rect 51540 7488 51592 7540
rect 51724 7463 51776 7472
rect 50160 7352 50212 7404
rect 51724 7429 51733 7463
rect 51733 7429 51767 7463
rect 51767 7429 51776 7463
rect 51724 7420 51776 7429
rect 52828 7420 52880 7472
rect 50804 7352 50856 7404
rect 51632 7352 51684 7404
rect 53656 7352 53708 7404
rect 54576 7352 54628 7404
rect 57704 7488 57756 7540
rect 3148 7284 3200 7336
rect 46572 7327 46624 7336
rect 46572 7293 46581 7327
rect 46581 7293 46615 7327
rect 46615 7293 46624 7327
rect 46572 7284 46624 7293
rect 47216 7327 47268 7336
rect 47216 7293 47225 7327
rect 47225 7293 47259 7327
rect 47259 7293 47268 7327
rect 47216 7284 47268 7293
rect 47860 7327 47912 7336
rect 47860 7293 47869 7327
rect 47869 7293 47903 7327
rect 47903 7293 47912 7327
rect 47860 7284 47912 7293
rect 48964 7327 49016 7336
rect 48964 7293 48973 7327
rect 48973 7293 49007 7327
rect 49007 7293 49016 7327
rect 48964 7284 49016 7293
rect 50620 7284 50672 7336
rect 52184 7284 52236 7336
rect 53288 7284 53340 7336
rect 53472 7284 53524 7336
rect 54392 7284 54444 7336
rect 56784 7352 56836 7404
rect 58164 7395 58216 7404
rect 58164 7361 58173 7395
rect 58173 7361 58207 7395
rect 58207 7361 58216 7395
rect 58164 7352 58216 7361
rect 57980 7259 58032 7268
rect 57980 7225 57989 7259
rect 57989 7225 58023 7259
rect 58023 7225 58032 7259
rect 57980 7216 58032 7225
rect 50160 7148 50212 7200
rect 50712 7191 50764 7200
rect 50712 7157 50721 7191
rect 50721 7157 50755 7191
rect 50755 7157 50764 7191
rect 50712 7148 50764 7157
rect 50896 7191 50948 7200
rect 50896 7157 50905 7191
rect 50905 7157 50939 7191
rect 50939 7157 50948 7191
rect 50896 7148 50948 7157
rect 52092 7148 52144 7200
rect 54760 7191 54812 7200
rect 54760 7157 54769 7191
rect 54769 7157 54803 7191
rect 54803 7157 54812 7191
rect 54760 7148 54812 7157
rect 57060 7191 57112 7200
rect 57060 7157 57069 7191
rect 57069 7157 57103 7191
rect 57103 7157 57112 7191
rect 57060 7148 57112 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 50326 7046 50378 7098
rect 50390 7046 50442 7098
rect 50454 7046 50506 7098
rect 50518 7046 50570 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 46572 6944 46624 6996
rect 52092 6987 52144 6996
rect 47860 6876 47912 6928
rect 51632 6876 51684 6928
rect 52092 6953 52101 6987
rect 52101 6953 52135 6987
rect 52135 6953 52144 6987
rect 52092 6944 52144 6953
rect 52736 6944 52788 6996
rect 57520 6944 57572 6996
rect 57980 6944 58032 6996
rect 54760 6876 54812 6928
rect 57060 6876 57112 6928
rect 45192 6808 45244 6860
rect 48780 6808 48832 6860
rect 50896 6808 50948 6860
rect 52092 6808 52144 6860
rect 53196 6851 53248 6860
rect 53196 6817 53205 6851
rect 53205 6817 53239 6851
rect 53239 6817 53248 6851
rect 53196 6808 53248 6817
rect 53380 6851 53432 6860
rect 53380 6817 53389 6851
rect 53389 6817 53423 6851
rect 53423 6817 53432 6851
rect 53380 6808 53432 6817
rect 2504 6740 2556 6792
rect 48688 6783 48740 6792
rect 48688 6749 48697 6783
rect 48697 6749 48731 6783
rect 48731 6749 48740 6783
rect 48688 6740 48740 6749
rect 49700 6740 49752 6792
rect 50804 6740 50856 6792
rect 52736 6740 52788 6792
rect 48596 6604 48648 6656
rect 51540 6672 51592 6724
rect 51908 6715 51960 6724
rect 51908 6681 51917 6715
rect 51917 6681 51951 6715
rect 51951 6681 51960 6715
rect 51908 6672 51960 6681
rect 55312 6808 55364 6860
rect 56968 6808 57020 6860
rect 53564 6740 53616 6792
rect 53840 6740 53892 6792
rect 57152 6740 57204 6792
rect 57428 6740 57480 6792
rect 49700 6604 49752 6656
rect 49976 6604 50028 6656
rect 50436 6604 50488 6656
rect 51172 6604 51224 6656
rect 53196 6604 53248 6656
rect 55220 6604 55272 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 51816 6400 51868 6452
rect 52368 6443 52420 6452
rect 52368 6409 52377 6443
rect 52377 6409 52411 6443
rect 52411 6409 52420 6443
rect 52368 6400 52420 6409
rect 53288 6400 53340 6452
rect 54208 6400 54260 6452
rect 2780 6196 2832 6248
rect 3332 6239 3384 6248
rect 3332 6205 3341 6239
rect 3341 6205 3375 6239
rect 3375 6205 3384 6239
rect 3332 6196 3384 6205
rect 45284 6239 45336 6248
rect 2320 6128 2372 6180
rect 45284 6205 45293 6239
rect 45293 6205 45327 6239
rect 45327 6205 45336 6239
rect 45284 6196 45336 6205
rect 46480 6196 46532 6248
rect 50896 6264 50948 6316
rect 51540 6264 51592 6316
rect 52460 6264 52512 6316
rect 52736 6307 52788 6316
rect 52736 6273 52745 6307
rect 52745 6273 52779 6307
rect 52779 6273 52788 6307
rect 52736 6264 52788 6273
rect 53564 6264 53616 6316
rect 57520 6307 57572 6316
rect 57520 6273 57529 6307
rect 57529 6273 57563 6307
rect 57563 6273 57572 6307
rect 57520 6264 57572 6273
rect 45376 6128 45428 6180
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 47768 6128 47820 6180
rect 48320 6196 48372 6248
rect 49516 6239 49568 6248
rect 49516 6205 49525 6239
rect 49525 6205 49559 6239
rect 49559 6205 49568 6239
rect 49516 6196 49568 6205
rect 49424 6128 49476 6180
rect 50436 6239 50488 6248
rect 50436 6205 50445 6239
rect 50445 6205 50479 6239
rect 50479 6205 50488 6239
rect 50436 6196 50488 6205
rect 50712 6196 50764 6248
rect 50068 6128 50120 6180
rect 51264 6196 51316 6248
rect 52092 6196 52144 6248
rect 52644 6239 52696 6248
rect 52644 6205 52653 6239
rect 52653 6205 52687 6239
rect 52687 6205 52696 6239
rect 52644 6196 52696 6205
rect 54024 6196 54076 6248
rect 54208 6239 54260 6248
rect 54208 6205 54217 6239
rect 54217 6205 54251 6239
rect 54251 6205 54260 6239
rect 54208 6196 54260 6205
rect 54300 6239 54352 6248
rect 54300 6205 54309 6239
rect 54309 6205 54343 6239
rect 54343 6205 54352 6239
rect 54300 6196 54352 6205
rect 54576 6196 54628 6248
rect 55220 6239 55272 6248
rect 55220 6205 55229 6239
rect 55229 6205 55263 6239
rect 55263 6205 55272 6239
rect 55220 6196 55272 6205
rect 51724 6171 51776 6180
rect 51724 6137 51733 6171
rect 51733 6137 51767 6171
rect 51767 6137 51776 6171
rect 51724 6128 51776 6137
rect 56508 6196 56560 6248
rect 58072 6196 58124 6248
rect 48688 6060 48740 6112
rect 48872 6103 48924 6112
rect 48872 6069 48881 6103
rect 48881 6069 48915 6103
rect 48915 6069 48924 6103
rect 48872 6060 48924 6069
rect 48964 6060 49016 6112
rect 49608 6060 49660 6112
rect 50620 6060 50672 6112
rect 50896 6060 50948 6112
rect 52460 6060 52512 6112
rect 53196 6060 53248 6112
rect 53748 6060 53800 6112
rect 57060 6103 57112 6112
rect 57060 6069 57069 6103
rect 57069 6069 57103 6103
rect 57103 6069 57112 6103
rect 57060 6060 57112 6069
rect 57980 6060 58032 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 50326 5958 50378 6010
rect 50390 5958 50442 6010
rect 50454 5958 50506 6010
rect 50518 5958 50570 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2780 5788 2832 5840
rect 3424 5720 3476 5772
rect 43812 5763 43864 5772
rect 43812 5729 43821 5763
rect 43821 5729 43855 5763
rect 43855 5729 43864 5763
rect 43812 5720 43864 5729
rect 49976 5788 50028 5840
rect 50068 5788 50120 5840
rect 51908 5856 51960 5908
rect 52000 5856 52052 5908
rect 52644 5856 52696 5908
rect 53196 5856 53248 5908
rect 55404 5856 55456 5908
rect 51356 5788 51408 5840
rect 47768 5763 47820 5772
rect 47768 5729 47777 5763
rect 47777 5729 47811 5763
rect 47811 5729 47820 5763
rect 47768 5720 47820 5729
rect 48412 5763 48464 5772
rect 48412 5729 48421 5763
rect 48421 5729 48455 5763
rect 48455 5729 48464 5763
rect 48412 5720 48464 5729
rect 49056 5763 49108 5772
rect 49056 5729 49065 5763
rect 49065 5729 49099 5763
rect 49099 5729 49108 5763
rect 49056 5720 49108 5729
rect 49608 5720 49660 5772
rect 50160 5763 50212 5772
rect 50160 5729 50169 5763
rect 50169 5729 50203 5763
rect 50203 5729 50212 5763
rect 50160 5720 50212 5729
rect 57980 5831 58032 5840
rect 57980 5797 57989 5831
rect 57989 5797 58023 5831
rect 58023 5797 58032 5831
rect 57980 5788 58032 5797
rect 52184 5763 52236 5772
rect 50896 5652 50948 5704
rect 50988 5652 51040 5704
rect 51632 5652 51684 5704
rect 52184 5729 52193 5763
rect 52193 5729 52227 5763
rect 52227 5729 52236 5763
rect 52184 5720 52236 5729
rect 52920 5763 52972 5772
rect 52920 5729 52929 5763
rect 52929 5729 52963 5763
rect 52963 5729 52972 5763
rect 52920 5720 52972 5729
rect 53288 5763 53340 5772
rect 52092 5652 52144 5704
rect 53288 5729 53297 5763
rect 53297 5729 53331 5763
rect 53331 5729 53340 5763
rect 53288 5720 53340 5729
rect 53748 5763 53800 5772
rect 53748 5729 53757 5763
rect 53757 5729 53791 5763
rect 53791 5729 53800 5763
rect 53748 5720 53800 5729
rect 54024 5720 54076 5772
rect 54760 5720 54812 5772
rect 56324 5720 56376 5772
rect 58164 5763 58216 5772
rect 58164 5729 58173 5763
rect 58173 5729 58207 5763
rect 58207 5729 58216 5763
rect 58164 5720 58216 5729
rect 56692 5695 56744 5704
rect 56692 5661 56701 5695
rect 56701 5661 56735 5695
rect 56735 5661 56744 5695
rect 56692 5652 56744 5661
rect 56784 5652 56836 5704
rect 48044 5584 48096 5636
rect 44640 5559 44692 5568
rect 44640 5525 44649 5559
rect 44649 5525 44683 5559
rect 44683 5525 44692 5559
rect 44640 5516 44692 5525
rect 44916 5559 44968 5568
rect 44916 5525 44925 5559
rect 44925 5525 44959 5559
rect 44959 5525 44968 5559
rect 44916 5516 44968 5525
rect 47124 5559 47176 5568
rect 47124 5525 47133 5559
rect 47133 5525 47167 5559
rect 47167 5525 47176 5559
rect 47124 5516 47176 5525
rect 48136 5516 48188 5568
rect 49332 5516 49384 5568
rect 56508 5584 56560 5636
rect 51172 5516 51224 5568
rect 51540 5559 51592 5568
rect 51540 5525 51549 5559
rect 51549 5525 51583 5559
rect 51583 5525 51592 5559
rect 51540 5516 51592 5525
rect 51908 5516 51960 5568
rect 52644 5516 52696 5568
rect 52828 5516 52880 5568
rect 54300 5516 54352 5568
rect 56416 5516 56468 5568
rect 56600 5516 56652 5568
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 49700 5312 49752 5364
rect 50712 5355 50764 5364
rect 50712 5321 50721 5355
rect 50721 5321 50755 5355
rect 50755 5321 50764 5355
rect 50712 5312 50764 5321
rect 51172 5312 51224 5364
rect 52184 5312 52236 5364
rect 53288 5312 53340 5364
rect 53380 5312 53432 5364
rect 55496 5312 55548 5364
rect 56968 5355 57020 5364
rect 56968 5321 56977 5355
rect 56977 5321 57011 5355
rect 57011 5321 57020 5355
rect 56968 5312 57020 5321
rect 43812 5244 43864 5296
rect 55772 5287 55824 5296
rect 2872 5176 2924 5228
rect 2964 5176 3016 5228
rect 49148 5176 49200 5228
rect 55772 5253 55781 5287
rect 55781 5253 55815 5287
rect 55815 5253 55824 5287
rect 55772 5244 55824 5253
rect 57152 5244 57204 5296
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 44088 5108 44140 5160
rect 45008 5151 45060 5160
rect 45008 5117 45017 5151
rect 45017 5117 45051 5151
rect 45051 5117 45060 5151
rect 45008 5108 45060 5117
rect 45652 5151 45704 5160
rect 45652 5117 45661 5151
rect 45661 5117 45695 5151
rect 45695 5117 45704 5151
rect 45652 5108 45704 5117
rect 46940 5108 46992 5160
rect 2320 5040 2372 5092
rect 2596 5083 2648 5092
rect 2596 5049 2605 5083
rect 2605 5049 2639 5083
rect 2639 5049 2648 5083
rect 2596 5040 2648 5049
rect 2780 4972 2832 5024
rect 47768 5108 47820 5160
rect 47860 5151 47912 5160
rect 47860 5117 47869 5151
rect 47869 5117 47903 5151
rect 47903 5117 47912 5151
rect 47860 5108 47912 5117
rect 48320 5108 48372 5160
rect 48780 5108 48832 5160
rect 49240 5108 49292 5160
rect 55312 5176 55364 5228
rect 50160 5108 50212 5160
rect 50712 5108 50764 5160
rect 51908 5151 51960 5160
rect 51908 5117 51917 5151
rect 51917 5117 51951 5151
rect 51951 5117 51960 5151
rect 51908 5108 51960 5117
rect 52092 5151 52144 5160
rect 52092 5117 52101 5151
rect 52101 5117 52135 5151
rect 52135 5117 52144 5151
rect 52092 5108 52144 5117
rect 52920 5151 52972 5160
rect 52920 5117 52929 5151
rect 52929 5117 52963 5151
rect 52963 5117 52972 5151
rect 52920 5108 52972 5117
rect 54024 5151 54076 5160
rect 54024 5117 54039 5151
rect 54039 5117 54073 5151
rect 54073 5117 54076 5151
rect 54208 5151 54260 5160
rect 54024 5108 54076 5117
rect 54208 5117 54217 5151
rect 54217 5117 54251 5151
rect 54251 5117 54260 5151
rect 54208 5108 54260 5117
rect 54392 5108 54444 5160
rect 55496 5108 55548 5160
rect 57060 5108 57112 5160
rect 49424 4972 49476 5024
rect 49976 5040 50028 5092
rect 56508 5040 56560 5092
rect 51080 4972 51132 5024
rect 51172 4972 51224 5024
rect 53380 4972 53432 5024
rect 53472 4972 53524 5024
rect 53840 4972 53892 5024
rect 54116 5015 54168 5024
rect 54116 4981 54125 5015
rect 54125 4981 54159 5015
rect 54159 4981 54168 5015
rect 54116 4972 54168 4981
rect 56232 4972 56284 5024
rect 57336 5015 57388 5024
rect 57336 4981 57345 5015
rect 57345 4981 57379 5015
rect 57379 4981 57388 5015
rect 57336 4972 57388 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 50326 4870 50378 4922
rect 50390 4870 50442 4922
rect 50454 4870 50506 4922
rect 50518 4870 50570 4922
rect 2596 4811 2648 4820
rect 2596 4777 2605 4811
rect 2605 4777 2639 4811
rect 2639 4777 2648 4811
rect 2596 4768 2648 4777
rect 45284 4768 45336 4820
rect 47768 4768 47820 4820
rect 47952 4768 48004 4820
rect 49056 4768 49108 4820
rect 49976 4811 50028 4820
rect 49976 4777 49985 4811
rect 49985 4777 50019 4811
rect 50019 4777 50028 4811
rect 49976 4768 50028 4777
rect 50160 4768 50212 4820
rect 55220 4768 55272 4820
rect 2780 4632 2832 4684
rect 3424 4632 3476 4684
rect 38108 4675 38160 4684
rect 38108 4641 38117 4675
rect 38117 4641 38151 4675
rect 38151 4641 38160 4675
rect 38108 4632 38160 4641
rect 46572 4632 46624 4684
rect 47860 4700 47912 4752
rect 50252 4700 50304 4752
rect 47308 4632 47360 4684
rect 47952 4632 48004 4684
rect 48780 4632 48832 4684
rect 49608 4632 49660 4684
rect 49884 4675 49936 4684
rect 49884 4641 49893 4675
rect 49893 4641 49927 4675
rect 49927 4641 49936 4675
rect 49884 4632 49936 4641
rect 50068 4675 50120 4684
rect 50068 4641 50077 4675
rect 50077 4641 50111 4675
rect 50111 4641 50120 4675
rect 50068 4632 50120 4641
rect 51540 4700 51592 4752
rect 54116 4700 54168 4752
rect 57152 4700 57204 4752
rect 3332 4564 3384 4616
rect 47400 4496 47452 4548
rect 47768 4496 47820 4548
rect 50712 4564 50764 4616
rect 50896 4564 50948 4616
rect 53380 4607 53432 4616
rect 53380 4573 53389 4607
rect 53389 4573 53423 4607
rect 53423 4573 53432 4607
rect 53380 4564 53432 4573
rect 57244 4564 57296 4616
rect 48136 4496 48188 4548
rect 51448 4496 51500 4548
rect 52920 4539 52972 4548
rect 52920 4505 52929 4539
rect 52929 4505 52963 4539
rect 52963 4505 52972 4539
rect 52920 4496 52972 4505
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 4620 4428 4672 4480
rect 34520 4471 34572 4480
rect 34520 4437 34529 4471
rect 34529 4437 34563 4471
rect 34563 4437 34572 4471
rect 34520 4428 34572 4437
rect 35900 4471 35952 4480
rect 35900 4437 35909 4471
rect 35909 4437 35943 4471
rect 35943 4437 35952 4471
rect 35900 4428 35952 4437
rect 36268 4428 36320 4480
rect 38476 4428 38528 4480
rect 38752 4471 38804 4480
rect 38752 4437 38761 4471
rect 38761 4437 38795 4471
rect 38795 4437 38804 4471
rect 38752 4428 38804 4437
rect 42800 4471 42852 4480
rect 42800 4437 42809 4471
rect 42809 4437 42843 4471
rect 42843 4437 42852 4471
rect 42800 4428 42852 4437
rect 43536 4471 43588 4480
rect 43536 4437 43545 4471
rect 43545 4437 43579 4471
rect 43579 4437 43588 4471
rect 43536 4428 43588 4437
rect 44180 4471 44232 4480
rect 44180 4437 44189 4471
rect 44189 4437 44223 4471
rect 44223 4437 44232 4471
rect 44180 4428 44232 4437
rect 45100 4471 45152 4480
rect 45100 4437 45109 4471
rect 45109 4437 45143 4471
rect 45143 4437 45152 4471
rect 45100 4428 45152 4437
rect 47676 4428 47728 4480
rect 47952 4471 48004 4480
rect 47952 4437 47961 4471
rect 47961 4437 47995 4471
rect 47995 4437 48004 4471
rect 47952 4428 48004 4437
rect 49240 4471 49292 4480
rect 49240 4437 49249 4471
rect 49249 4437 49283 4471
rect 49283 4437 49292 4471
rect 49240 4428 49292 4437
rect 49792 4428 49844 4480
rect 50896 4428 50948 4480
rect 51080 4428 51132 4480
rect 55588 4496 55640 4548
rect 54760 4471 54812 4480
rect 54760 4437 54769 4471
rect 54769 4437 54803 4471
rect 54803 4437 54812 4471
rect 54760 4428 54812 4437
rect 56968 4471 57020 4480
rect 56968 4437 56977 4471
rect 56977 4437 57011 4471
rect 57011 4437 57020 4471
rect 56968 4428 57020 4437
rect 57980 4471 58032 4480
rect 57980 4437 57989 4471
rect 57989 4437 58023 4471
rect 58023 4437 58032 4471
rect 57980 4428 58032 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 44640 4224 44692 4276
rect 40040 4156 40092 4208
rect 41604 4156 41656 4208
rect 42708 4156 42760 4208
rect 46388 4156 46440 4208
rect 46572 4199 46624 4208
rect 46572 4165 46581 4199
rect 46581 4165 46615 4199
rect 46615 4165 46624 4199
rect 46572 4156 46624 4165
rect 3056 4088 3108 4140
rect 4620 4088 4672 4140
rect 3700 4020 3752 4072
rect 4160 4020 4212 4072
rect 33416 4020 33468 4072
rect 33968 4063 34020 4072
rect 33968 4029 33977 4063
rect 33977 4029 34011 4063
rect 34011 4029 34020 4063
rect 33968 4020 34020 4029
rect 37188 4088 37240 4140
rect 43352 4088 43404 4140
rect 47492 4156 47544 4208
rect 50252 4156 50304 4208
rect 55588 4224 55640 4276
rect 56508 4224 56560 4276
rect 57336 4156 57388 4208
rect 37372 4020 37424 4072
rect 38108 4020 38160 4072
rect 39120 4063 39172 4072
rect 39120 4029 39129 4063
rect 39129 4029 39163 4063
rect 39163 4029 39172 4063
rect 39120 4020 39172 4029
rect 40500 4063 40552 4072
rect 40500 4029 40509 4063
rect 40509 4029 40543 4063
rect 40543 4029 40552 4063
rect 40500 4020 40552 4029
rect 44640 4020 44692 4072
rect 45744 4020 45796 4072
rect 49516 4088 49568 4140
rect 50344 4088 50396 4140
rect 56692 4131 56744 4140
rect 56692 4097 56701 4131
rect 56701 4097 56735 4131
rect 56735 4097 56744 4131
rect 56692 4088 56744 4097
rect 46388 4063 46440 4072
rect 46388 4029 46397 4063
rect 46397 4029 46431 4063
rect 46431 4029 46440 4063
rect 46388 4020 46440 4029
rect 46480 4020 46532 4072
rect 1400 3884 1452 3936
rect 2964 3884 3016 3936
rect 33784 3884 33836 3936
rect 34796 3884 34848 3936
rect 35532 3927 35584 3936
rect 35532 3893 35541 3927
rect 35541 3893 35575 3927
rect 35575 3893 35584 3927
rect 35532 3884 35584 3893
rect 36176 3927 36228 3936
rect 36176 3893 36185 3927
rect 36185 3893 36219 3927
rect 36219 3893 36228 3927
rect 36176 3884 36228 3893
rect 39028 3884 39080 3936
rect 42892 3884 42944 3936
rect 44364 3884 44416 3936
rect 45468 3884 45520 3936
rect 47032 3952 47084 4004
rect 47308 4020 47360 4072
rect 49608 4020 49660 4072
rect 50896 4063 50948 4072
rect 50344 3952 50396 4004
rect 50896 4029 50905 4063
rect 50905 4029 50939 4063
rect 50939 4029 50948 4063
rect 50896 4020 50948 4029
rect 51724 4063 51776 4072
rect 51724 4029 51733 4063
rect 51733 4029 51767 4063
rect 51767 4029 51776 4063
rect 51724 4020 51776 4029
rect 52736 4020 52788 4072
rect 48136 3884 48188 3936
rect 49424 3884 49476 3936
rect 50068 3884 50120 3936
rect 50988 3884 51040 3936
rect 53104 3995 53156 4004
rect 53104 3961 53113 3995
rect 53113 3961 53147 3995
rect 53147 3961 53156 3995
rect 53104 3952 53156 3961
rect 55036 3952 55088 4004
rect 55588 3952 55640 4004
rect 54208 3884 54260 3936
rect 54484 3927 54536 3936
rect 54484 3893 54493 3927
rect 54493 3893 54527 3927
rect 54527 3893 54536 3927
rect 54484 3884 54536 3893
rect 55680 3884 55732 3936
rect 57980 4063 58032 4072
rect 56048 3995 56100 4004
rect 56048 3961 56057 3995
rect 56057 3961 56091 3995
rect 56091 3961 56100 3995
rect 56048 3952 56100 3961
rect 57980 4029 57989 4063
rect 57989 4029 58023 4063
rect 58023 4029 58032 4063
rect 57980 4020 58032 4029
rect 56600 3952 56652 4004
rect 58164 3995 58216 4004
rect 58164 3961 58173 3995
rect 58173 3961 58207 3995
rect 58207 3961 58216 3995
rect 58164 3952 58216 3961
rect 57244 3884 57296 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 50326 3782 50378 3834
rect 50390 3782 50442 3834
rect 50454 3782 50506 3834
rect 50518 3782 50570 3834
rect 45560 3680 45612 3732
rect 47032 3680 47084 3732
rect 47216 3680 47268 3732
rect 48044 3680 48096 3732
rect 1676 3612 1728 3664
rect 2872 3544 2924 3596
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 3976 3476 4028 3528
rect 2320 3451 2372 3460
rect 2320 3417 2329 3451
rect 2329 3417 2363 3451
rect 2363 3417 2372 3451
rect 2320 3408 2372 3417
rect 2412 3408 2464 3460
rect 6092 3544 6144 3596
rect 28540 3587 28592 3596
rect 28540 3553 28549 3587
rect 28549 3553 28583 3587
rect 28583 3553 28592 3587
rect 28540 3544 28592 3553
rect 29460 3544 29512 3596
rect 31300 3544 31352 3596
rect 33324 3587 33376 3596
rect 33324 3553 33333 3587
rect 33333 3553 33367 3587
rect 33367 3553 33376 3587
rect 33324 3544 33376 3553
rect 34244 3587 34296 3596
rect 34244 3553 34253 3587
rect 34253 3553 34287 3587
rect 34287 3553 34296 3587
rect 34244 3544 34296 3553
rect 35808 3587 35860 3596
rect 35808 3553 35817 3587
rect 35817 3553 35851 3587
rect 35851 3553 35860 3587
rect 35808 3544 35860 3553
rect 37096 3587 37148 3596
rect 37096 3553 37105 3587
rect 37105 3553 37139 3587
rect 37139 3553 37148 3587
rect 37096 3544 37148 3553
rect 38660 3544 38712 3596
rect 38936 3587 38988 3596
rect 38936 3553 38945 3587
rect 38945 3553 38979 3587
rect 38979 3553 38988 3587
rect 38936 3544 38988 3553
rect 39764 3587 39816 3596
rect 39764 3553 39773 3587
rect 39773 3553 39807 3587
rect 39807 3553 39816 3587
rect 39764 3544 39816 3553
rect 46388 3612 46440 3664
rect 48780 3612 48832 3664
rect 51448 3612 51500 3664
rect 52368 3612 52420 3664
rect 52460 3612 52512 3664
rect 43076 3544 43128 3596
rect 43352 3587 43404 3596
rect 43352 3553 43353 3587
rect 43353 3553 43387 3587
rect 43387 3553 43404 3587
rect 43352 3544 43404 3553
rect 44640 3587 44692 3596
rect 44640 3553 44649 3587
rect 44649 3553 44683 3587
rect 44683 3553 44692 3587
rect 44640 3544 44692 3553
rect 45744 3544 45796 3596
rect 46296 3587 46348 3596
rect 46296 3553 46305 3587
rect 46305 3553 46339 3587
rect 46339 3553 46348 3587
rect 46296 3544 46348 3553
rect 47032 3587 47084 3596
rect 47032 3553 47041 3587
rect 47041 3553 47075 3587
rect 47075 3553 47084 3587
rect 47032 3544 47084 3553
rect 47768 3587 47820 3596
rect 47768 3553 47777 3587
rect 47777 3553 47811 3587
rect 47811 3553 47820 3587
rect 47768 3544 47820 3553
rect 47860 3544 47912 3596
rect 49608 3544 49660 3596
rect 50160 3544 50212 3596
rect 52644 3544 52696 3596
rect 53012 3587 53064 3596
rect 53012 3553 53021 3587
rect 53021 3553 53055 3587
rect 53055 3553 53064 3587
rect 53012 3544 53064 3553
rect 2872 3340 2924 3392
rect 4620 3340 4672 3392
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 31116 3340 31168 3392
rect 31392 3383 31444 3392
rect 31392 3349 31401 3383
rect 31401 3349 31435 3383
rect 31435 3349 31444 3383
rect 31392 3340 31444 3349
rect 32036 3383 32088 3392
rect 32036 3349 32045 3383
rect 32045 3349 32079 3383
rect 32079 3349 32088 3383
rect 32036 3340 32088 3349
rect 33140 3340 33192 3392
rect 33232 3340 33284 3392
rect 34152 3340 34204 3392
rect 35256 3340 35308 3392
rect 37004 3340 37056 3392
rect 37924 3340 37976 3392
rect 38844 3340 38896 3392
rect 40224 3340 40276 3392
rect 41788 3340 41840 3392
rect 41972 3383 42024 3392
rect 41972 3349 41981 3383
rect 41981 3349 42015 3383
rect 42015 3349 42024 3383
rect 41972 3340 42024 3349
rect 42616 3340 42668 3392
rect 47584 3476 47636 3528
rect 47952 3476 48004 3528
rect 55220 3544 55272 3596
rect 55772 3612 55824 3664
rect 56876 3655 56928 3664
rect 56876 3621 56885 3655
rect 56885 3621 56919 3655
rect 56919 3621 56928 3655
rect 56876 3612 56928 3621
rect 53656 3476 53708 3528
rect 56416 3544 56468 3596
rect 57612 3544 57664 3596
rect 48964 3408 49016 3460
rect 49056 3408 49108 3460
rect 55220 3408 55272 3460
rect 55772 3451 55824 3460
rect 55772 3417 55781 3451
rect 55781 3417 55815 3451
rect 55815 3417 55824 3451
rect 55772 3408 55824 3417
rect 45376 3340 45428 3392
rect 46480 3340 46532 3392
rect 47308 3340 47360 3392
rect 48228 3340 48280 3392
rect 49608 3383 49660 3392
rect 49608 3349 49617 3383
rect 49617 3349 49651 3383
rect 49651 3349 49660 3383
rect 49608 3340 49660 3349
rect 52000 3340 52052 3392
rect 52920 3340 52972 3392
rect 54392 3383 54444 3392
rect 54392 3349 54401 3383
rect 54401 3349 54435 3383
rect 54435 3349 54444 3383
rect 54392 3340 54444 3349
rect 55312 3340 55364 3392
rect 56416 3340 56468 3392
rect 57980 3383 58032 3392
rect 57980 3349 57989 3383
rect 57989 3349 58023 3383
rect 58023 3349 58032 3383
rect 57980 3340 58032 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 3148 3179 3200 3188
rect 3148 3145 3157 3179
rect 3157 3145 3191 3179
rect 3191 3145 3200 3179
rect 3148 3136 3200 3145
rect 3976 3136 4028 3188
rect 34244 3179 34296 3188
rect 34244 3145 34253 3179
rect 34253 3145 34287 3179
rect 34287 3145 34296 3179
rect 34244 3136 34296 3145
rect 37372 3179 37424 3188
rect 37372 3145 37381 3179
rect 37381 3145 37415 3179
rect 37415 3145 37424 3179
rect 37372 3136 37424 3145
rect 38660 3179 38712 3188
rect 38660 3145 38669 3179
rect 38669 3145 38703 3179
rect 38703 3145 38712 3179
rect 38660 3136 38712 3145
rect 43536 3136 43588 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 4068 3068 4120 3120
rect 4712 3068 4764 3120
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 480 2932 532 2984
rect 3700 2932 3752 2984
rect 5356 2932 5408 2984
rect 7012 2932 7064 2984
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 33968 3000 34020 3052
rect 35532 3043 35584 3052
rect 35532 3009 35541 3043
rect 35541 3009 35575 3043
rect 35575 3009 35584 3043
rect 35532 3000 35584 3009
rect 38476 3043 38528 3052
rect 38476 3009 38485 3043
rect 38485 3009 38519 3043
rect 38519 3009 38528 3043
rect 38476 3000 38528 3009
rect 40500 3000 40552 3052
rect 41972 3000 42024 3052
rect 31300 2975 31352 2984
rect 31300 2941 31309 2975
rect 31309 2941 31343 2975
rect 31343 2941 31352 2975
rect 31300 2932 31352 2941
rect 33416 2932 33468 2984
rect 3976 2907 4028 2916
rect 3976 2873 3985 2907
rect 3985 2873 4019 2907
rect 4019 2873 4028 2907
rect 3976 2864 4028 2873
rect 4160 2907 4212 2916
rect 4160 2873 4169 2907
rect 4169 2873 4203 2907
rect 4203 2873 4212 2907
rect 4160 2864 4212 2873
rect 3240 2796 3292 2848
rect 5632 2864 5684 2916
rect 31944 2907 31996 2916
rect 31944 2873 31953 2907
rect 31953 2873 31987 2907
rect 31987 2873 31996 2907
rect 31944 2864 31996 2873
rect 32312 2864 32364 2916
rect 4344 2796 4396 2848
rect 5080 2796 5132 2848
rect 5264 2839 5316 2848
rect 5264 2805 5273 2839
rect 5273 2805 5307 2839
rect 5307 2805 5316 2839
rect 5264 2796 5316 2805
rect 30564 2839 30616 2848
rect 30564 2805 30573 2839
rect 30573 2805 30607 2839
rect 30607 2805 30616 2839
rect 30564 2796 30616 2805
rect 32220 2796 32272 2848
rect 35900 2932 35952 2984
rect 37188 2975 37240 2984
rect 37188 2941 37197 2975
rect 37197 2941 37231 2975
rect 37231 2941 37240 2975
rect 37188 2932 37240 2941
rect 39120 2932 39172 2984
rect 37372 2864 37424 2916
rect 39764 2932 39816 2984
rect 36084 2796 36136 2848
rect 42800 2932 42852 2984
rect 45468 3068 45520 3120
rect 47032 3136 47084 3188
rect 47860 3179 47912 3188
rect 47860 3145 47869 3179
rect 47869 3145 47903 3179
rect 47903 3145 47912 3179
rect 47860 3136 47912 3145
rect 49240 3136 49292 3188
rect 51540 3136 51592 3188
rect 53012 3179 53064 3188
rect 53012 3145 53021 3179
rect 53021 3145 53055 3179
rect 53055 3145 53064 3179
rect 53012 3136 53064 3145
rect 53104 3136 53156 3188
rect 54852 3136 54904 3188
rect 55036 3136 55088 3188
rect 56232 3136 56284 3188
rect 57244 3111 57296 3120
rect 45652 3000 45704 3052
rect 47124 3000 47176 3052
rect 47400 3043 47452 3052
rect 47400 3009 47409 3043
rect 47409 3009 47443 3043
rect 47443 3009 47452 3043
rect 47400 3000 47452 3009
rect 48596 3000 48648 3052
rect 48964 3043 49016 3052
rect 48964 3009 48973 3043
rect 48973 3009 49007 3043
rect 49007 3009 49016 3043
rect 48964 3000 49016 3009
rect 41972 2907 42024 2916
rect 41972 2873 41981 2907
rect 41981 2873 42015 2907
rect 42015 2873 42024 2907
rect 41972 2864 42024 2873
rect 44732 2907 44784 2916
rect 44732 2873 44741 2907
rect 44741 2873 44775 2907
rect 44775 2873 44784 2907
rect 44732 2864 44784 2873
rect 40776 2796 40828 2848
rect 41696 2796 41748 2848
rect 44456 2796 44508 2848
rect 46756 2932 46808 2984
rect 49332 2932 49384 2984
rect 55496 3000 55548 3052
rect 57244 3077 57253 3111
rect 57253 3077 57287 3111
rect 57287 3077 57296 3111
rect 57244 3068 57296 3077
rect 58072 3136 58124 3188
rect 58532 3068 58584 3120
rect 57060 3043 57112 3052
rect 57060 3009 57069 3043
rect 57069 3009 57103 3043
rect 57103 3009 57112 3043
rect 57060 3000 57112 3009
rect 52368 2975 52420 2984
rect 52368 2941 52377 2975
rect 52377 2941 52411 2975
rect 52411 2941 52420 2975
rect 52368 2932 52420 2941
rect 45284 2864 45336 2916
rect 49056 2864 49108 2916
rect 50712 2907 50764 2916
rect 50712 2873 50721 2907
rect 50721 2873 50755 2907
rect 50755 2873 50764 2907
rect 50712 2864 50764 2873
rect 51448 2907 51500 2916
rect 51448 2873 51457 2907
rect 51457 2873 51491 2907
rect 51491 2873 51500 2907
rect 51448 2864 51500 2873
rect 51632 2864 51684 2916
rect 54116 2907 54168 2916
rect 54116 2873 54125 2907
rect 54125 2873 54159 2907
rect 54159 2873 54168 2907
rect 54116 2864 54168 2873
rect 54392 2932 54444 2984
rect 55956 2932 56008 2984
rect 55864 2864 55916 2916
rect 59452 2864 59504 2916
rect 48412 2796 48464 2848
rect 49148 2796 49200 2848
rect 50160 2796 50212 2848
rect 51080 2796 51132 2848
rect 53840 2796 53892 2848
rect 54760 2796 54812 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 50326 2694 50378 2746
rect 50390 2694 50442 2746
rect 50454 2694 50506 2746
rect 50518 2694 50570 2746
rect 3976 2592 4028 2644
rect 35808 2592 35860 2644
rect 37096 2592 37148 2644
rect 38936 2592 38988 2644
rect 44732 2592 44784 2644
rect 46296 2592 46348 2644
rect 47768 2592 47820 2644
rect 50712 2592 50764 2644
rect 51448 2592 51500 2644
rect 54116 2592 54168 2644
rect 55588 2635 55640 2644
rect 55588 2601 55597 2635
rect 55597 2601 55631 2635
rect 55631 2601 55640 2635
rect 55588 2592 55640 2601
rect 56324 2592 56376 2644
rect 5080 2524 5132 2576
rect 4620 2456 4672 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 5632 2456 5684 2508
rect 30564 2524 30616 2576
rect 46756 2524 46808 2576
rect 48872 2524 48924 2576
rect 7932 2456 7984 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 11704 2456 11756 2508
rect 12624 2456 12676 2508
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 14464 2456 14516 2508
rect 15476 2456 15528 2508
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 17316 2456 17368 2508
rect 18236 2499 18288 2508
rect 18236 2465 18245 2499
rect 18245 2465 18279 2499
rect 18279 2465 18288 2499
rect 18236 2456 18288 2465
rect 19156 2499 19208 2508
rect 19156 2465 19165 2499
rect 19165 2465 19199 2499
rect 19199 2465 19208 2499
rect 19156 2456 19208 2465
rect 20076 2456 20128 2508
rect 21088 2499 21140 2508
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 22008 2456 22060 2508
rect 22928 2499 22980 2508
rect 22928 2465 22937 2499
rect 22937 2465 22971 2499
rect 22971 2465 22980 2499
rect 22928 2456 22980 2465
rect 23848 2499 23900 2508
rect 23848 2465 23857 2499
rect 23857 2465 23891 2499
rect 23891 2465 23900 2499
rect 23848 2456 23900 2465
rect 24768 2456 24820 2508
rect 25780 2456 25832 2508
rect 26700 2456 26752 2508
rect 27620 2456 27672 2508
rect 4344 2388 4396 2440
rect 5264 2388 5316 2440
rect 30472 2320 30524 2372
rect 31392 2456 31444 2508
rect 32036 2499 32088 2508
rect 32036 2465 32045 2499
rect 32045 2465 32079 2499
rect 32079 2465 32088 2499
rect 32036 2456 32088 2465
rect 32220 2499 32272 2508
rect 32220 2465 32229 2499
rect 32229 2465 32263 2499
rect 32263 2465 32272 2499
rect 32220 2456 32272 2465
rect 33140 2456 33192 2508
rect 33784 2499 33836 2508
rect 33784 2465 33793 2499
rect 33793 2465 33827 2499
rect 33827 2465 33836 2499
rect 33784 2456 33836 2465
rect 34520 2456 34572 2508
rect 34796 2456 34848 2508
rect 36176 2456 36228 2508
rect 38752 2456 38804 2508
rect 39028 2456 39080 2508
rect 40040 2499 40092 2508
rect 40040 2465 40049 2499
rect 40049 2465 40083 2499
rect 40083 2465 40092 2499
rect 40040 2456 40092 2465
rect 40224 2499 40276 2508
rect 40224 2465 40233 2499
rect 40233 2465 40267 2499
rect 40267 2465 40276 2499
rect 40224 2456 40276 2465
rect 41604 2499 41656 2508
rect 41604 2465 41613 2499
rect 41613 2465 41647 2499
rect 41647 2465 41656 2499
rect 41604 2456 41656 2465
rect 41788 2499 41840 2508
rect 41788 2465 41797 2499
rect 41797 2465 41831 2499
rect 41831 2465 41840 2499
rect 41788 2456 41840 2465
rect 42708 2499 42760 2508
rect 42708 2465 42717 2499
rect 42717 2465 42751 2499
rect 42751 2465 42760 2499
rect 42708 2456 42760 2465
rect 42892 2499 42944 2508
rect 42892 2465 42901 2499
rect 42901 2465 42935 2499
rect 42935 2465 42944 2499
rect 42892 2456 42944 2465
rect 44180 2456 44232 2508
rect 44364 2456 44416 2508
rect 45100 2456 45152 2508
rect 45560 2499 45612 2508
rect 45560 2465 45569 2499
rect 45569 2465 45603 2499
rect 45603 2465 45612 2499
rect 46940 2499 46992 2508
rect 45560 2456 45612 2465
rect 46940 2465 46949 2499
rect 46949 2465 46983 2499
rect 46983 2465 46992 2499
rect 46940 2456 46992 2465
rect 47216 2456 47268 2508
rect 48780 2456 48832 2508
rect 49700 2456 49752 2508
rect 31116 2431 31168 2440
rect 31116 2397 31125 2431
rect 31125 2397 31159 2431
rect 31159 2397 31168 2431
rect 31116 2388 31168 2397
rect 36268 2431 36320 2440
rect 36268 2397 36277 2431
rect 36277 2397 36311 2431
rect 36311 2397 36320 2431
rect 36268 2388 36320 2397
rect 43536 2388 43588 2440
rect 31944 2320 31996 2372
rect 33324 2320 33376 2372
rect 39764 2320 39816 2372
rect 41972 2363 42024 2372
rect 41972 2329 41981 2363
rect 41981 2329 42015 2363
rect 42015 2329 42024 2363
rect 41972 2320 42024 2329
rect 43076 2363 43128 2372
rect 43076 2329 43085 2363
rect 43085 2329 43119 2363
rect 43119 2329 43128 2363
rect 43076 2320 43128 2329
rect 45192 2320 45244 2372
rect 50804 2388 50856 2440
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 31392 2252 31444 2304
rect 49516 2320 49568 2372
rect 51356 2456 51408 2508
rect 51816 2388 51868 2440
rect 51172 2320 51224 2372
rect 52644 2363 52696 2372
rect 52644 2329 52653 2363
rect 52653 2329 52687 2363
rect 52687 2329 52696 2363
rect 52644 2320 52696 2329
rect 55220 2524 55272 2576
rect 57980 2567 58032 2576
rect 57980 2533 57989 2567
rect 57989 2533 58023 2567
rect 58023 2533 58032 2567
rect 57980 2524 58032 2533
rect 55312 2456 55364 2508
rect 55128 2431 55180 2440
rect 54668 2252 54720 2304
rect 55128 2397 55137 2431
rect 55137 2397 55171 2431
rect 55171 2397 55180 2431
rect 55128 2388 55180 2397
rect 56232 2431 56284 2440
rect 56232 2397 56241 2431
rect 56241 2397 56275 2431
rect 56275 2397 56284 2431
rect 56232 2388 56284 2397
rect 57888 2252 57940 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 44916 2048 44968 2100
rect 54668 2048 54720 2100
rect 47676 1980 47728 2032
rect 51172 1980 51224 2032
rect 48136 1912 48188 1964
rect 55128 1912 55180 1964
rect 49424 1844 49476 1896
rect 56232 1844 56284 1896
rect 54484 1640 54536 1692
rect 56692 1640 56744 1692
rect 44088 1300 44140 1352
rect 55220 1300 55272 1352
<< metal2 >>
rect 386 59200 442 60000
rect 1122 59200 1178 60000
rect 1950 59200 2006 60000
rect 2686 59200 2742 60000
rect 2778 59528 2834 59537
rect 2778 59463 2834 59472
rect 400 56506 428 59200
rect 388 56500 440 56506
rect 388 56442 440 56448
rect 1136 56302 1164 59200
rect 1398 57624 1454 57633
rect 1398 57559 1454 57568
rect 1412 57390 1440 57559
rect 1400 57384 1452 57390
rect 1400 57326 1452 57332
rect 1400 56908 1452 56914
rect 1400 56850 1452 56856
rect 1412 56681 1440 56850
rect 1398 56672 1454 56681
rect 1398 56607 1454 56616
rect 1308 56500 1360 56506
rect 1308 56442 1360 56448
rect 1124 56296 1176 56302
rect 1124 56238 1176 56244
rect 1320 25974 1348 56442
rect 1964 56302 1992 59200
rect 2042 58576 2098 58585
rect 2042 58511 2098 58520
rect 2056 57390 2084 58511
rect 2044 57384 2096 57390
rect 2044 57326 2096 57332
rect 2700 56914 2728 59200
rect 2792 57390 2820 59463
rect 3514 59200 3570 60000
rect 4250 59200 4306 60000
rect 5078 59200 5134 60000
rect 5906 59200 5962 60000
rect 6642 59200 6698 60000
rect 7470 59200 7526 60000
rect 8206 59200 8262 60000
rect 9034 59200 9090 60000
rect 9770 59200 9826 60000
rect 10598 59200 10654 60000
rect 11426 59200 11482 60000
rect 12162 59200 12218 60000
rect 12990 59200 13046 60000
rect 13726 59200 13782 60000
rect 14554 59200 14610 60000
rect 15382 59200 15438 60000
rect 16118 59200 16174 60000
rect 16946 59200 17002 60000
rect 17682 59200 17738 60000
rect 18510 59200 18566 60000
rect 19246 59200 19302 60000
rect 20074 59200 20130 60000
rect 20902 59200 20958 60000
rect 21638 59200 21694 60000
rect 22466 59200 22522 60000
rect 23202 59200 23258 60000
rect 24030 59200 24086 60000
rect 24766 59200 24822 60000
rect 25594 59200 25650 60000
rect 26422 59200 26478 60000
rect 27158 59200 27214 60000
rect 27986 59200 28042 60000
rect 28722 59200 28778 60000
rect 29550 59200 29606 60000
rect 30378 59200 30434 60000
rect 31114 59200 31170 60000
rect 31942 59200 31998 60000
rect 32678 59200 32734 60000
rect 33506 59200 33562 60000
rect 34242 59200 34298 60000
rect 35070 59200 35126 60000
rect 35898 59200 35954 60000
rect 36634 59200 36690 60000
rect 37462 59200 37518 60000
rect 38198 59200 38254 60000
rect 39026 59200 39082 60000
rect 39762 59200 39818 60000
rect 40590 59200 40646 60000
rect 41418 59200 41474 60000
rect 42154 59200 42210 60000
rect 42982 59200 43038 60000
rect 43718 59200 43774 60000
rect 44546 59200 44602 60000
rect 45374 59200 45430 60000
rect 46110 59200 46166 60000
rect 46938 59200 46994 60000
rect 47674 59200 47730 60000
rect 48502 59200 48558 60000
rect 49238 59200 49294 60000
rect 50066 59200 50122 60000
rect 50894 59200 50950 60000
rect 51630 59200 51686 60000
rect 52458 59200 52514 60000
rect 53194 59200 53250 60000
rect 54022 59200 54078 60000
rect 54758 59200 54814 60000
rect 55586 59200 55642 60000
rect 56414 59200 56470 60000
rect 56506 59664 56562 59673
rect 56506 59599 56562 59608
rect 2780 57384 2832 57390
rect 2780 57326 2832 57332
rect 2688 56908 2740 56914
rect 2688 56850 2740 56856
rect 3332 56704 3384 56710
rect 3332 56646 3384 56652
rect 3344 56370 3372 56646
rect 3332 56364 3384 56370
rect 3332 56306 3384 56312
rect 1952 56296 2004 56302
rect 1952 56238 2004 56244
rect 3528 55826 3556 59200
rect 4264 58290 4292 59200
rect 4264 58262 4660 58290
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4632 57526 4660 58262
rect 4620 57520 4672 57526
rect 4620 57462 4672 57468
rect 5092 57390 5120 59200
rect 5920 57390 5948 59200
rect 6656 57458 6684 59200
rect 6644 57452 6696 57458
rect 6644 57394 6696 57400
rect 7484 57390 7512 59200
rect 8220 57390 8248 59200
rect 9048 57390 9076 59200
rect 9784 57390 9812 59200
rect 10612 57390 10640 59200
rect 11440 57390 11468 59200
rect 5080 57384 5132 57390
rect 5080 57326 5132 57332
rect 5908 57384 5960 57390
rect 5908 57326 5960 57332
rect 7472 57384 7524 57390
rect 7472 57326 7524 57332
rect 8208 57384 8260 57390
rect 8208 57326 8260 57332
rect 9036 57384 9088 57390
rect 9036 57326 9088 57332
rect 9772 57384 9824 57390
rect 9772 57326 9824 57332
rect 10600 57384 10652 57390
rect 10600 57326 10652 57332
rect 11428 57384 11480 57390
rect 12176 57372 12204 59200
rect 13004 57390 13032 59200
rect 12440 57384 12492 57390
rect 12176 57344 12440 57372
rect 11428 57326 11480 57332
rect 12440 57326 12492 57332
rect 12992 57384 13044 57390
rect 13740 57372 13768 59200
rect 14568 57458 14596 59200
rect 15396 57458 15424 59200
rect 14556 57452 14608 57458
rect 14556 57394 14608 57400
rect 15384 57452 15436 57458
rect 15384 57394 15436 57400
rect 13820 57384 13872 57390
rect 13740 57344 13820 57372
rect 12992 57326 13044 57332
rect 13820 57326 13872 57332
rect 4620 57316 4672 57322
rect 4620 57258 4672 57264
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4632 56506 4660 57258
rect 5080 57248 5132 57254
rect 5080 57190 5132 57196
rect 4712 56840 4764 56846
rect 4712 56782 4764 56788
rect 4724 56506 4752 56782
rect 4620 56500 4672 56506
rect 4620 56442 4672 56448
rect 4712 56500 4764 56506
rect 4712 56442 4764 56448
rect 3700 56228 3752 56234
rect 3700 56170 3752 56176
rect 1400 55820 1452 55826
rect 1400 55762 1452 55768
rect 3516 55820 3568 55826
rect 3516 55762 3568 55768
rect 1412 55729 1440 55762
rect 1398 55720 1454 55729
rect 1398 55655 1454 55664
rect 1398 54768 1454 54777
rect 1398 54703 1400 54712
rect 1452 54703 1454 54712
rect 1400 54674 1452 54680
rect 1398 53816 1454 53825
rect 1398 53751 1454 53760
rect 1412 53650 1440 53751
rect 1400 53644 1452 53650
rect 1400 53586 1452 53592
rect 1400 53032 1452 53038
rect 1400 52974 1452 52980
rect 1412 52873 1440 52974
rect 1398 52864 1454 52873
rect 1398 52799 1454 52808
rect 1400 51944 1452 51950
rect 1398 51912 1400 51921
rect 1452 51912 1454 51921
rect 1398 51847 1454 51856
rect 1398 51096 1454 51105
rect 1398 51031 1454 51040
rect 1412 50862 1440 51031
rect 1400 50856 1452 50862
rect 1400 50798 1452 50804
rect 1400 50380 1452 50386
rect 1400 50322 1452 50328
rect 1412 50153 1440 50322
rect 1398 50144 1454 50153
rect 1398 50079 1454 50088
rect 1400 49292 1452 49298
rect 1400 49234 1452 49240
rect 1412 49201 1440 49234
rect 1398 49192 1454 49201
rect 1398 49127 1454 49136
rect 1398 48240 1454 48249
rect 1398 48175 1400 48184
rect 1452 48175 1454 48184
rect 1400 48146 1452 48152
rect 1398 47288 1454 47297
rect 1398 47223 1454 47232
rect 1412 47122 1440 47223
rect 1400 47116 1452 47122
rect 1400 47058 1452 47064
rect 1400 46504 1452 46510
rect 1400 46446 1452 46452
rect 1412 46345 1440 46446
rect 1398 46336 1454 46345
rect 1398 46271 1454 46280
rect 1400 45416 1452 45422
rect 1398 45384 1400 45393
rect 1452 45384 1454 45393
rect 1398 45319 1454 45328
rect 1398 44432 1454 44441
rect 1398 44367 1454 44376
rect 1412 44334 1440 44367
rect 1400 44328 1452 44334
rect 1400 44270 1452 44276
rect 1398 43480 1454 43489
rect 1398 43415 1454 43424
rect 1412 43246 1440 43415
rect 1400 43240 1452 43246
rect 1400 43182 1452 43188
rect 1400 42764 1452 42770
rect 1400 42706 1452 42712
rect 1412 42673 1440 42706
rect 1398 42664 1454 42673
rect 1398 42599 1454 42608
rect 1398 41712 1454 41721
rect 1398 41647 1400 41656
rect 1452 41647 1454 41656
rect 1400 41618 1452 41624
rect 1398 40760 1454 40769
rect 1398 40695 1454 40704
rect 1412 40594 1440 40695
rect 1400 40588 1452 40594
rect 1400 40530 1452 40536
rect 1400 39976 1452 39982
rect 1400 39918 1452 39924
rect 1412 39817 1440 39918
rect 1398 39808 1454 39817
rect 1398 39743 1454 39752
rect 1400 38888 1452 38894
rect 1398 38856 1400 38865
rect 1452 38856 1454 38865
rect 1398 38791 1454 38800
rect 1398 37904 1454 37913
rect 1398 37839 1454 37848
rect 1412 37806 1440 37839
rect 1400 37800 1452 37806
rect 1400 37742 1452 37748
rect 1398 36952 1454 36961
rect 1398 36887 1454 36896
rect 1412 36718 1440 36887
rect 1400 36712 1452 36718
rect 1400 36654 1452 36660
rect 1400 36236 1452 36242
rect 1400 36178 1452 36184
rect 1412 36009 1440 36178
rect 1398 36000 1454 36009
rect 1398 35935 1454 35944
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 1412 35057 1440 35090
rect 1398 35048 1454 35057
rect 1398 34983 1454 34992
rect 1398 34232 1454 34241
rect 1398 34167 1454 34176
rect 1412 34066 1440 34167
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1412 33289 1440 33390
rect 1398 33280 1454 33289
rect 1398 33215 1454 33224
rect 1400 32360 1452 32366
rect 1398 32328 1400 32337
rect 1452 32328 1454 32337
rect 1398 32263 1454 32272
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1412 31278 1440 31311
rect 1400 31272 1452 31278
rect 1400 31214 1452 31220
rect 1400 30796 1452 30802
rect 1400 30738 1452 30744
rect 1412 30433 1440 30738
rect 1398 30424 1454 30433
rect 1398 30359 1454 30368
rect 1860 30116 1912 30122
rect 1860 30058 1912 30064
rect 1400 29504 1452 29510
rect 1400 29446 1452 29452
rect 1412 28529 1440 29446
rect 1872 29306 1900 30058
rect 1952 30048 2004 30054
rect 1952 29990 2004 29996
rect 1964 29481 1992 29990
rect 2136 29708 2188 29714
rect 2136 29650 2188 29656
rect 1950 29472 2006 29481
rect 1950 29407 2006 29416
rect 1860 29300 1912 29306
rect 1860 29242 1912 29248
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1398 28520 1454 28529
rect 1398 28455 1454 28464
rect 1780 28218 1808 29038
rect 2148 28490 2176 29650
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2700 29170 2728 29446
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 3148 28552 3200 28558
rect 3148 28494 3200 28500
rect 2136 28484 2188 28490
rect 2136 28426 2188 28432
rect 3160 28218 3188 28494
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 2688 28008 2740 28014
rect 2688 27950 2740 27956
rect 2044 27940 2096 27946
rect 2044 27882 2096 27888
rect 1952 27872 2004 27878
rect 1952 27814 2004 27820
rect 1964 27577 1992 27814
rect 1950 27568 2006 27577
rect 1950 27503 2006 27512
rect 2056 27402 2084 27882
rect 2504 27464 2556 27470
rect 2504 27406 2556 27412
rect 2044 27396 2096 27402
rect 2044 27338 2096 27344
rect 2516 27130 2544 27406
rect 2504 27124 2556 27130
rect 2504 27066 2556 27072
rect 2700 26926 2728 27950
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 3344 27130 3372 27474
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2320 26852 2372 26858
rect 2320 26794 2372 26800
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 1964 26625 1992 26726
rect 1950 26616 2006 26625
rect 2332 26586 2360 26794
rect 1950 26551 2006 26560
rect 2320 26580 2372 26586
rect 2320 26522 2372 26528
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1872 26042 1900 26318
rect 1860 26036 1912 26042
rect 1860 25978 1912 25984
rect 1308 25968 1360 25974
rect 1308 25910 1360 25916
rect 2780 25832 2832 25838
rect 2042 25800 2098 25809
rect 1860 25764 1912 25770
rect 2780 25774 2832 25780
rect 2042 25735 2044 25744
rect 1860 25706 1912 25712
rect 2096 25735 2098 25744
rect 2044 25706 2096 25712
rect 1872 25498 1900 25706
rect 1860 25492 1912 25498
rect 1860 25434 1912 25440
rect 2792 25362 2820 25774
rect 2780 25356 2832 25362
rect 2780 25298 2832 25304
rect 2778 24848 2834 24857
rect 2778 24783 2780 24792
rect 2832 24783 2834 24792
rect 2780 24754 2832 24760
rect 2044 24676 2096 24682
rect 2044 24618 2096 24624
rect 2596 24676 2648 24682
rect 2596 24618 2648 24624
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1964 23905 1992 24550
rect 1950 23896 2006 23905
rect 2056 23866 2084 24618
rect 2608 24410 2636 24618
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 1950 23831 2006 23840
rect 2044 23860 2096 23866
rect 2044 23802 2096 23808
rect 1860 23656 1912 23662
rect 1860 23598 1912 23604
rect 1872 23322 1900 23598
rect 1860 23316 1912 23322
rect 1860 23258 1912 23264
rect 1860 23180 1912 23186
rect 1860 23122 1912 23128
rect 1584 23044 1636 23050
rect 1584 22986 1636 22992
rect 1596 22642 1624 22986
rect 1872 22778 1900 23122
rect 1952 22976 2004 22982
rect 1950 22944 1952 22953
rect 2004 22944 2006 22953
rect 1950 22879 2006 22888
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1584 22636 1636 22642
rect 1584 22578 1636 22584
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1872 21690 1900 22034
rect 2884 22030 2912 26862
rect 3148 25764 3200 25770
rect 3148 25706 3200 25712
rect 3160 25362 3188 25706
rect 3148 25356 3200 25362
rect 3148 25298 3200 25304
rect 3160 24750 3188 25298
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3160 23186 3188 24686
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3252 24206 3280 24550
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3148 23180 3200 23186
rect 3148 23122 3200 23128
rect 3160 22778 3188 23122
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3160 22574 3188 22714
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 2976 22166 3004 22510
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 2872 22024 2924 22030
rect 2042 21992 2098 22001
rect 2872 21966 2924 21972
rect 2042 21927 2044 21936
rect 2096 21927 2098 21936
rect 2044 21898 2096 21904
rect 1860 21684 1912 21690
rect 1860 21626 1912 21632
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2778 21040 2834 21049
rect 1860 21004 1912 21010
rect 1860 20946 1912 20952
rect 2596 21004 2648 21010
rect 2778 20975 2780 20984
rect 2596 20946 2648 20952
rect 2832 20975 2834 20984
rect 2780 20946 2832 20952
rect 1872 20058 1900 20946
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1964 20097 1992 20742
rect 2608 20602 2636 20946
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2884 20466 2912 21286
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 1950 20088 2006 20097
rect 1860 20052 1912 20058
rect 1950 20023 2006 20032
rect 1860 19994 1912 20000
rect 2976 19922 3004 22102
rect 3148 21616 3200 21622
rect 3148 21558 3200 21564
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 3068 20398 3096 21422
rect 3160 20482 3188 21558
rect 3240 21412 3292 21418
rect 3240 21354 3292 21360
rect 3252 20602 3280 21354
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3160 20454 3280 20482
rect 3252 20398 3280 20454
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 1860 19236 1912 19242
rect 1860 19178 1912 19184
rect 2596 19236 2648 19242
rect 2596 19178 2648 19184
rect 2780 19236 2832 19242
rect 2780 19178 2832 19184
rect 1872 18426 1900 19178
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 1768 18216 1820 18222
rect 1964 18193 1992 19110
rect 2608 18970 2636 19178
rect 2792 19145 2820 19178
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2884 18834 2912 19246
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 1768 18158 1820 18164
rect 1950 18184 2006 18193
rect 1780 17882 1808 18158
rect 1950 18119 2006 18128
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1872 17338 1900 17682
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 17377 1992 17478
rect 1950 17368 2006 17377
rect 1860 17332 1912 17338
rect 1950 17303 2006 17312
rect 1860 17274 1912 17280
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2516 16794 2544 17070
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16250 1900 16594
rect 1952 16448 2004 16454
rect 1950 16416 1952 16425
rect 2004 16416 2006 16425
rect 1950 16351 2006 16360
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1860 15564 1912 15570
rect 1860 15506 1912 15512
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 1872 14618 1900 15506
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1964 14521 1992 15302
rect 2608 15162 2636 15506
rect 2778 15464 2834 15473
rect 2778 15399 2780 15408
rect 2832 15399 2834 15408
rect 2780 15370 2832 15376
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2976 14958 3004 19858
rect 3252 19718 3280 20334
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3252 18834 3280 19654
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3252 17746 3280 18770
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 3068 16046 3096 16594
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 16114 3188 16390
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3068 15162 3096 15982
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 1950 14512 2006 14521
rect 1950 14447 2006 14456
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2516 14074 2544 14350
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2044 13796 2096 13802
rect 2044 13738 2096 13744
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13569 1992 13670
rect 1950 13560 2006 13569
rect 1950 13495 2006 13504
rect 2056 13258 2084 13738
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2976 12986 3004 14894
rect 3068 13870 3096 15098
rect 3252 15026 3280 15846
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13326 3188 13670
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1780 11898 1808 12174
rect 1872 12170 1900 12650
rect 1952 12640 2004 12646
rect 1950 12608 1952 12617
rect 2004 12608 2006 12617
rect 1950 12543 2006 12552
rect 2976 12306 3004 12922
rect 2964 12300 3016 12306
rect 2964 12242 3016 12248
rect 1860 12164 1912 12170
rect 1860 12106 1912 12112
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 2884 11694 2912 12038
rect 2872 11688 2924 11694
rect 2778 11656 2834 11665
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 2596 11620 2648 11626
rect 2872 11630 2924 11636
rect 2778 11591 2780 11600
rect 2596 11562 2648 11568
rect 2832 11591 2834 11600
rect 2780 11562 2832 11568
rect 1872 10810 1900 11562
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1964 10713 1992 11494
rect 2608 11354 2636 11562
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2884 11218 2912 11630
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 1950 10704 2006 10713
rect 1950 10639 2006 10648
rect 2504 10600 2556 10606
rect 2504 10542 2556 10548
rect 2516 10266 2544 10542
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2884 10130 2912 11154
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3344 10130 3372 10474
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 3332 10124 3384 10130
rect 3332 10066 3384 10072
rect 1872 9722 1900 10066
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9761 1992 9862
rect 1950 9752 2006 9761
rect 1860 9716 1912 9722
rect 1950 9687 2006 9696
rect 1860 9658 1912 9664
rect 2884 9518 2912 10066
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9042 2912 9454
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 2778 8936 2834 8945
rect 1688 8634 1716 8910
rect 2778 8871 2834 8880
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 2608 8430 2636 8774
rect 2792 8566 2820 8871
rect 3712 8566 3740 56170
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 3976 28620 4028 28626
rect 3976 28562 4028 28568
rect 3988 28218 4016 28562
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 3976 28212 4028 28218
rect 3976 28154 4028 28160
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 19990 3924 20198
rect 3884 19984 3936 19990
rect 3884 19926 3936 19932
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4080 15094 4108 15982
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3976 14340 4028 14346
rect 3976 14282 4028 14288
rect 3988 14074 4016 14282
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 5092 13394 5120 57190
rect 16132 56914 16160 59200
rect 16960 57390 16988 59200
rect 17696 57390 17724 59200
rect 18524 57390 18552 59200
rect 16948 57384 17000 57390
rect 16948 57326 17000 57332
rect 17684 57384 17736 57390
rect 17684 57326 17736 57332
rect 18512 57384 18564 57390
rect 19260 57372 19288 59200
rect 20088 57458 20116 59200
rect 20076 57452 20128 57458
rect 20076 57394 20128 57400
rect 19340 57384 19392 57390
rect 19260 57344 19340 57372
rect 18512 57326 18564 57332
rect 20916 57372 20944 59200
rect 21652 57390 21680 59200
rect 22480 57458 22508 59200
rect 23216 57458 23244 59200
rect 24044 57526 24072 59200
rect 24032 57520 24084 57526
rect 24032 57462 24084 57468
rect 22468 57452 22520 57458
rect 22468 57394 22520 57400
rect 23204 57452 23256 57458
rect 23204 57394 23256 57400
rect 20996 57384 21048 57390
rect 20916 57344 20996 57372
rect 19340 57326 19392 57332
rect 20996 57326 21048 57332
rect 21640 57384 21692 57390
rect 21640 57326 21692 57332
rect 24780 57338 24808 59200
rect 25608 57474 25636 59200
rect 25608 57458 25728 57474
rect 25608 57452 25740 57458
rect 25608 57446 25688 57452
rect 25688 57394 25740 57400
rect 24780 57310 24900 57338
rect 24872 57254 24900 57310
rect 24860 57248 24912 57254
rect 24860 57190 24912 57196
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 26436 56914 26464 59200
rect 27172 57390 27200 59200
rect 28000 57458 28028 59200
rect 28736 57474 28764 59200
rect 29564 57474 29592 59200
rect 27988 57452 28040 57458
rect 28736 57446 29040 57474
rect 29564 57446 29684 57474
rect 30392 57458 30420 59200
rect 31128 57458 31156 59200
rect 31956 57526 31984 59200
rect 31944 57520 31996 57526
rect 31944 57462 31996 57468
rect 27988 57394 28040 57400
rect 29012 57390 29040 57446
rect 29656 57390 29684 57446
rect 30380 57452 30432 57458
rect 30380 57394 30432 57400
rect 31116 57452 31168 57458
rect 31116 57394 31168 57400
rect 27160 57384 27212 57390
rect 27160 57326 27212 57332
rect 29000 57384 29052 57390
rect 29000 57326 29052 57332
rect 29644 57384 29696 57390
rect 29644 57326 29696 57332
rect 32692 57322 32720 59200
rect 33520 57458 33548 59200
rect 33508 57452 33560 57458
rect 33508 57394 33560 57400
rect 32680 57316 32732 57322
rect 32680 57258 32732 57264
rect 34256 56914 34284 59200
rect 35084 57882 35112 59200
rect 35084 57854 35296 57882
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 35268 57390 35296 57854
rect 35256 57384 35308 57390
rect 35256 57326 35308 57332
rect 35912 57322 35940 59200
rect 36648 57458 36676 59200
rect 36636 57452 36688 57458
rect 36636 57394 36688 57400
rect 37476 57372 37504 59200
rect 37648 57384 37700 57390
rect 37476 57344 37648 57372
rect 37648 57326 37700 57332
rect 38212 57322 38240 59200
rect 39040 57458 39068 59200
rect 39028 57452 39080 57458
rect 39028 57394 39080 57400
rect 35900 57316 35952 57322
rect 35900 57258 35952 57264
rect 38200 57316 38252 57322
rect 38200 57258 38252 57264
rect 39776 56914 39804 59200
rect 40604 56914 40632 59200
rect 41432 56914 41460 59200
rect 42168 57390 42196 59200
rect 42996 57390 43024 59200
rect 43732 57390 43760 59200
rect 44560 57390 44588 59200
rect 45388 57458 45416 59200
rect 45376 57452 45428 57458
rect 45376 57394 45428 57400
rect 46124 57390 46152 59200
rect 42156 57384 42208 57390
rect 42156 57326 42208 57332
rect 42984 57384 43036 57390
rect 42984 57326 43036 57332
rect 43720 57384 43772 57390
rect 43720 57326 43772 57332
rect 44548 57384 44600 57390
rect 44548 57326 44600 57332
rect 46112 57384 46164 57390
rect 46952 57372 46980 59200
rect 47688 57390 47716 59200
rect 48516 57390 48544 59200
rect 49252 57458 49280 59200
rect 50080 57458 50108 59200
rect 49240 57452 49292 57458
rect 49240 57394 49292 57400
rect 50068 57452 50120 57458
rect 50068 57394 50120 57400
rect 47032 57384 47084 57390
rect 46952 57344 47032 57372
rect 46112 57326 46164 57332
rect 47032 57326 47084 57332
rect 47676 57384 47728 57390
rect 47676 57326 47728 57332
rect 48504 57384 48556 57390
rect 48504 57326 48556 57332
rect 50300 57148 50596 57168
rect 50356 57146 50380 57148
rect 50436 57146 50460 57148
rect 50516 57146 50540 57148
rect 50378 57094 50380 57146
rect 50442 57094 50454 57146
rect 50516 57094 50518 57146
rect 50356 57092 50380 57094
rect 50436 57092 50460 57094
rect 50516 57092 50540 57094
rect 50300 57072 50596 57092
rect 16120 56908 16172 56914
rect 16120 56850 16172 56856
rect 26424 56908 26476 56914
rect 26424 56850 26476 56856
rect 34244 56908 34296 56914
rect 34244 56850 34296 56856
rect 39764 56908 39816 56914
rect 39764 56850 39816 56856
rect 40592 56908 40644 56914
rect 40592 56850 40644 56856
rect 41420 56908 41472 56914
rect 50908 56896 50936 59200
rect 51644 56914 51672 59200
rect 52472 56914 52500 59200
rect 53104 57316 53156 57322
rect 53104 57258 53156 57264
rect 53116 57050 53144 57258
rect 53104 57044 53156 57050
rect 53104 56986 53156 56992
rect 51080 56908 51132 56914
rect 50908 56868 51080 56896
rect 41420 56850 41472 56856
rect 51080 56850 51132 56856
rect 51632 56908 51684 56914
rect 51632 56850 51684 56856
rect 52460 56908 52512 56914
rect 52460 56850 52512 56856
rect 5448 56772 5500 56778
rect 5448 56714 5500 56720
rect 5460 56506 5488 56714
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 5448 56500 5500 56506
rect 5448 56442 5500 56448
rect 53208 56302 53236 59200
rect 53840 57316 53892 57322
rect 53840 57258 53892 57264
rect 53852 56846 53880 57258
rect 53840 56840 53892 56846
rect 53840 56782 53892 56788
rect 53932 56500 53984 56506
rect 53932 56442 53984 56448
rect 53196 56296 53248 56302
rect 53196 56238 53248 56244
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 50300 56060 50596 56080
rect 50356 56058 50380 56060
rect 50436 56058 50460 56060
rect 50516 56058 50540 56060
rect 50378 56006 50380 56058
rect 50442 56006 50454 56058
rect 50516 56006 50518 56058
rect 50356 56004 50380 56006
rect 50436 56004 50460 56006
rect 50516 56004 50540 56006
rect 50300 55984 50596 56004
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 53944 55214 53972 56442
rect 54036 55826 54064 59200
rect 54772 56506 54800 59200
rect 55600 59106 55628 59200
rect 55324 59078 55628 59106
rect 56322 59120 56378 59129
rect 55034 58440 55090 58449
rect 55034 58375 55090 58384
rect 54942 58168 54998 58177
rect 54942 58103 54998 58112
rect 54956 57458 54984 58103
rect 55048 57526 55076 58375
rect 55220 58336 55272 58342
rect 55220 58278 55272 58284
rect 55036 57520 55088 57526
rect 55232 57474 55260 58278
rect 55036 57462 55088 57468
rect 54944 57452 54996 57458
rect 54944 57394 54996 57400
rect 55140 57446 55260 57474
rect 54760 56500 54812 56506
rect 54760 56442 54812 56448
rect 55140 56370 55168 57446
rect 55128 56364 55180 56370
rect 55128 56306 55180 56312
rect 54024 55820 54076 55826
rect 54024 55762 54076 55768
rect 55324 55758 55352 59078
rect 56322 59055 56378 59064
rect 55494 58576 55550 58585
rect 55494 58511 55550 58520
rect 55508 57526 55536 58511
rect 56336 58449 56364 59055
rect 56322 58440 56378 58449
rect 56322 58375 56378 58384
rect 56428 58342 56456 59200
rect 56416 58336 56468 58342
rect 56416 58278 56468 58284
rect 56520 58177 56548 59599
rect 57150 59200 57206 60000
rect 57978 59200 58034 60000
rect 58714 59200 58770 60000
rect 59542 59200 59598 60000
rect 56506 58168 56562 58177
rect 56506 58103 56562 58112
rect 56506 58032 56562 58041
rect 56506 57967 56562 57976
rect 55496 57520 55548 57526
rect 55496 57462 55548 57468
rect 55586 57488 55642 57497
rect 55586 57423 55642 57432
rect 55404 57384 55456 57390
rect 55404 57326 55456 57332
rect 55416 56438 55444 57326
rect 55600 56914 55628 57423
rect 55772 57316 55824 57322
rect 55772 57258 55824 57264
rect 55784 56914 55812 57258
rect 55588 56908 55640 56914
rect 55588 56850 55640 56856
rect 55772 56908 55824 56914
rect 55772 56850 55824 56856
rect 55404 56432 55456 56438
rect 55404 56374 55456 56380
rect 55784 56302 55812 56850
rect 56324 56840 56376 56846
rect 56324 56782 56376 56788
rect 56140 56772 56192 56778
rect 56140 56714 56192 56720
rect 56152 56302 56180 56714
rect 56336 56506 56364 56782
rect 56324 56500 56376 56506
rect 56324 56442 56376 56448
rect 56232 56432 56284 56438
rect 56232 56374 56284 56380
rect 55772 56296 55824 56302
rect 55772 56238 55824 56244
rect 56140 56296 56192 56302
rect 56140 56238 56192 56244
rect 55678 55992 55734 56001
rect 55678 55927 55734 55936
rect 55692 55826 55720 55927
rect 55784 55826 55812 56238
rect 55680 55820 55732 55826
rect 55680 55762 55732 55768
rect 55772 55820 55824 55826
rect 55772 55762 55824 55768
rect 55312 55752 55364 55758
rect 55312 55694 55364 55700
rect 55496 55616 55548 55622
rect 55496 55558 55548 55564
rect 53932 55208 53984 55214
rect 53932 55150 53984 55156
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 50300 54972 50596 54992
rect 50356 54970 50380 54972
rect 50436 54970 50460 54972
rect 50516 54970 50540 54972
rect 50378 54918 50380 54970
rect 50442 54918 50454 54970
rect 50516 54918 50518 54970
rect 50356 54916 50380 54918
rect 50436 54916 50460 54918
rect 50516 54916 50540 54918
rect 50300 54896 50596 54916
rect 55312 54732 55364 54738
rect 55312 54674 55364 54680
rect 54944 54528 54996 54534
rect 54944 54470 54996 54476
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 54956 54194 54984 54470
rect 54944 54188 54996 54194
rect 54944 54130 54996 54136
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 50300 53884 50596 53904
rect 50356 53882 50380 53884
rect 50436 53882 50460 53884
rect 50516 53882 50540 53884
rect 50378 53830 50380 53882
rect 50442 53830 50454 53882
rect 50516 53830 50518 53882
rect 50356 53828 50380 53830
rect 50436 53828 50460 53830
rect 50516 53828 50540 53830
rect 50300 53808 50596 53828
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 50300 52796 50596 52816
rect 50356 52794 50380 52796
rect 50436 52794 50460 52796
rect 50516 52794 50540 52796
rect 50378 52742 50380 52794
rect 50442 52742 50454 52794
rect 50516 52742 50518 52794
rect 50356 52740 50380 52742
rect 50436 52740 50460 52742
rect 50516 52740 50540 52742
rect 50300 52720 50596 52740
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 50300 51708 50596 51728
rect 50356 51706 50380 51708
rect 50436 51706 50460 51708
rect 50516 51706 50540 51708
rect 50378 51654 50380 51706
rect 50442 51654 50454 51706
rect 50516 51654 50518 51706
rect 50356 51652 50380 51654
rect 50436 51652 50460 51654
rect 50516 51652 50540 51654
rect 50300 51632 50596 51652
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 50300 50620 50596 50640
rect 50356 50618 50380 50620
rect 50436 50618 50460 50620
rect 50516 50618 50540 50620
rect 50378 50566 50380 50618
rect 50442 50566 50454 50618
rect 50516 50566 50518 50618
rect 50356 50564 50380 50566
rect 50436 50564 50460 50566
rect 50516 50564 50540 50566
rect 50300 50544 50596 50564
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 55220 49768 55272 49774
rect 55218 49736 55220 49745
rect 55272 49736 55274 49745
rect 55218 49671 55274 49680
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 50300 49532 50596 49552
rect 50356 49530 50380 49532
rect 50436 49530 50460 49532
rect 50516 49530 50540 49532
rect 50378 49478 50380 49530
rect 50442 49478 50454 49530
rect 50516 49478 50518 49530
rect 50356 49476 50380 49478
rect 50436 49476 50460 49478
rect 50516 49476 50540 49478
rect 50300 49456 50596 49476
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 50300 48444 50596 48464
rect 50356 48442 50380 48444
rect 50436 48442 50460 48444
rect 50516 48442 50540 48444
rect 50378 48390 50380 48442
rect 50442 48390 50454 48442
rect 50516 48390 50518 48442
rect 50356 48388 50380 48390
rect 50436 48388 50460 48390
rect 50516 48388 50540 48390
rect 50300 48368 50596 48388
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 50300 47356 50596 47376
rect 50356 47354 50380 47356
rect 50436 47354 50460 47356
rect 50516 47354 50540 47356
rect 50378 47302 50380 47354
rect 50442 47302 50454 47354
rect 50516 47302 50518 47354
rect 50356 47300 50380 47302
rect 50436 47300 50460 47302
rect 50516 47300 50540 47302
rect 50300 47280 50596 47300
rect 55220 47116 55272 47122
rect 55220 47058 55272 47064
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 55232 46753 55260 47058
rect 55218 46744 55274 46753
rect 55218 46679 55274 46688
rect 55036 46572 55088 46578
rect 55036 46514 55088 46520
rect 54760 46504 54812 46510
rect 54760 46446 54812 46452
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 50300 46268 50596 46288
rect 50356 46266 50380 46268
rect 50436 46266 50460 46268
rect 50516 46266 50540 46268
rect 50378 46214 50380 46266
rect 50442 46214 50454 46266
rect 50516 46214 50518 46266
rect 50356 46212 50380 46214
rect 50436 46212 50460 46214
rect 50516 46212 50540 46214
rect 50300 46192 50596 46212
rect 51540 45892 51592 45898
rect 51540 45834 51592 45840
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 50300 45180 50596 45200
rect 50356 45178 50380 45180
rect 50436 45178 50460 45180
rect 50516 45178 50540 45180
rect 50378 45126 50380 45178
rect 50442 45126 50454 45178
rect 50516 45126 50518 45178
rect 50356 45124 50380 45126
rect 50436 45124 50460 45126
rect 50516 45124 50540 45126
rect 50300 45104 50596 45124
rect 51264 44872 51316 44878
rect 51264 44814 51316 44820
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 51276 44538 51304 44814
rect 51080 44532 51132 44538
rect 51080 44474 51132 44480
rect 51264 44532 51316 44538
rect 51264 44474 51316 44480
rect 50712 44328 50764 44334
rect 50712 44270 50764 44276
rect 50620 44260 50672 44266
rect 50620 44202 50672 44208
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 50632 43994 50660 44202
rect 50620 43988 50672 43994
rect 50620 43930 50672 43936
rect 50724 43926 50752 44270
rect 50712 43920 50764 43926
rect 50712 43862 50764 43868
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 50620 43240 50672 43246
rect 50620 43182 50672 43188
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 50632 42906 50660 43182
rect 50620 42900 50672 42906
rect 50620 42842 50672 42848
rect 50528 42832 50580 42838
rect 50528 42774 50580 42780
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 50436 42288 50488 42294
rect 50434 42256 50436 42265
rect 50488 42256 50490 42265
rect 50540 42226 50568 42774
rect 50434 42191 50490 42200
rect 50528 42220 50580 42226
rect 50528 42162 50580 42168
rect 49424 42152 49476 42158
rect 49422 42120 49424 42129
rect 49476 42120 49478 42129
rect 49422 42055 49478 42064
rect 50160 42016 50212 42022
rect 50160 41958 50212 41964
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 50068 41676 50120 41682
rect 50068 41618 50120 41624
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 50080 39982 50108 41618
rect 50068 39976 50120 39982
rect 50068 39918 50120 39924
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 49700 38412 49752 38418
rect 49700 38354 49752 38360
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 49056 37664 49108 37670
rect 49056 37606 49108 37612
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 49068 37330 49096 37606
rect 49712 37330 49740 38354
rect 50068 38208 50120 38214
rect 50068 38150 50120 38156
rect 50080 37806 50108 38150
rect 50068 37800 50120 37806
rect 50068 37742 50120 37748
rect 49056 37324 49108 37330
rect 49056 37266 49108 37272
rect 49700 37324 49752 37330
rect 49700 37266 49752 37272
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 49712 35154 49740 37266
rect 49792 37256 49844 37262
rect 49790 37224 49792 37233
rect 49844 37224 49846 37233
rect 49790 37159 49846 37168
rect 50172 36718 50200 41958
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 50620 40996 50672 41002
rect 50620 40938 50672 40944
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 50632 40662 50660 40938
rect 50620 40656 50672 40662
rect 50620 40598 50672 40604
rect 50620 40520 50672 40526
rect 50724 40474 50752 43862
rect 50988 42764 51040 42770
rect 50988 42706 51040 42712
rect 51000 42362 51028 42706
rect 51092 42566 51120 44474
rect 51448 44192 51500 44198
rect 51448 44134 51500 44140
rect 51460 43858 51488 44134
rect 51552 43994 51580 45834
rect 53932 45416 53984 45422
rect 53932 45358 53984 45364
rect 54208 45416 54260 45422
rect 54208 45358 54260 45364
rect 52920 45348 52972 45354
rect 52920 45290 52972 45296
rect 52736 45076 52788 45082
rect 52736 45018 52788 45024
rect 52092 44940 52144 44946
rect 52092 44882 52144 44888
rect 52104 44538 52132 44882
rect 52092 44532 52144 44538
rect 52092 44474 52144 44480
rect 52552 44396 52604 44402
rect 52552 44338 52604 44344
rect 52460 44328 52512 44334
rect 52460 44270 52512 44276
rect 51540 43988 51592 43994
rect 51540 43930 51592 43936
rect 51172 43852 51224 43858
rect 51172 43794 51224 43800
rect 51448 43852 51500 43858
rect 51448 43794 51500 43800
rect 51184 43314 51212 43794
rect 51172 43308 51224 43314
rect 51172 43250 51224 43256
rect 51552 43178 51580 43930
rect 51632 43240 51684 43246
rect 51632 43182 51684 43188
rect 52092 43240 52144 43246
rect 52092 43182 52144 43188
rect 51540 43172 51592 43178
rect 51540 43114 51592 43120
rect 51172 43104 51224 43110
rect 51172 43046 51224 43052
rect 51448 43104 51500 43110
rect 51448 43046 51500 43052
rect 51184 42838 51212 43046
rect 51172 42832 51224 42838
rect 51172 42774 51224 42780
rect 51080 42560 51132 42566
rect 51080 42502 51132 42508
rect 51172 42560 51224 42566
rect 51172 42502 51224 42508
rect 50988 42356 51040 42362
rect 50988 42298 51040 42304
rect 51092 41070 51120 42502
rect 51184 42158 51212 42502
rect 51172 42152 51224 42158
rect 51172 42094 51224 42100
rect 51337 42152 51389 42158
rect 51460 42140 51488 43046
rect 51552 42770 51580 43114
rect 51644 42906 51672 43182
rect 52104 42906 52132 43182
rect 51632 42900 51684 42906
rect 51632 42842 51684 42848
rect 52092 42900 52144 42906
rect 52092 42842 52144 42848
rect 51540 42764 51592 42770
rect 51540 42706 51592 42712
rect 51632 42560 51684 42566
rect 51632 42502 51684 42508
rect 51389 42112 51488 42140
rect 51337 42094 51389 42100
rect 51460 41682 51488 42112
rect 51644 41682 51672 42502
rect 52184 42288 52236 42294
rect 52182 42256 52184 42265
rect 52236 42256 52238 42265
rect 52182 42191 52238 42200
rect 52092 42152 52144 42158
rect 52092 42094 52144 42100
rect 52472 42106 52500 44270
rect 52564 43994 52592 44338
rect 52552 43988 52604 43994
rect 52552 43930 52604 43936
rect 52644 43920 52696 43926
rect 52644 43862 52696 43868
rect 52656 43450 52684 43862
rect 52748 43858 52776 45018
rect 52932 44334 52960 45290
rect 53944 44878 53972 45358
rect 54116 45280 54168 45286
rect 54116 45222 54168 45228
rect 54128 44946 54156 45222
rect 54220 45014 54248 45358
rect 54208 45008 54260 45014
rect 54208 44950 54260 44956
rect 54116 44940 54168 44946
rect 54116 44882 54168 44888
rect 54300 44940 54352 44946
rect 54300 44882 54352 44888
rect 53932 44872 53984 44878
rect 53932 44814 53984 44820
rect 52920 44328 52972 44334
rect 52920 44270 52972 44276
rect 54312 43858 54340 44882
rect 54392 44804 54444 44810
rect 54392 44746 54444 44752
rect 54404 44334 54432 44746
rect 54392 44328 54444 44334
rect 54392 44270 54444 44276
rect 54484 44328 54536 44334
rect 54484 44270 54536 44276
rect 54404 43858 54432 44270
rect 52736 43852 52788 43858
rect 52736 43794 52788 43800
rect 53196 43852 53248 43858
rect 53196 43794 53248 43800
rect 54116 43852 54168 43858
rect 54116 43794 54168 43800
rect 54300 43852 54352 43858
rect 54300 43794 54352 43800
rect 54392 43852 54444 43858
rect 54392 43794 54444 43800
rect 52644 43444 52696 43450
rect 52644 43386 52696 43392
rect 52748 43382 52776 43794
rect 52736 43376 52788 43382
rect 52736 43318 52788 43324
rect 52644 43308 52696 43314
rect 52644 43250 52696 43256
rect 52656 43194 52684 43250
rect 52656 43166 52776 43194
rect 52748 42634 52776 43166
rect 52920 43172 52972 43178
rect 52920 43114 52972 43120
rect 52828 42832 52880 42838
rect 52828 42774 52880 42780
rect 52736 42628 52788 42634
rect 52736 42570 52788 42576
rect 52748 42158 52776 42570
rect 52736 42152 52788 42158
rect 52104 41818 52132 42094
rect 52472 42078 52592 42106
rect 52736 42094 52788 42100
rect 52840 42090 52868 42774
rect 52932 42770 52960 43114
rect 52920 42764 52972 42770
rect 52920 42706 52972 42712
rect 52932 42158 52960 42706
rect 52920 42152 52972 42158
rect 52920 42094 52972 42100
rect 52092 41812 52144 41818
rect 52092 41754 52144 41760
rect 51448 41676 51500 41682
rect 51448 41618 51500 41624
rect 51632 41676 51684 41682
rect 51632 41618 51684 41624
rect 52460 41540 52512 41546
rect 52460 41482 52512 41488
rect 51080 41064 51132 41070
rect 51080 41006 51132 41012
rect 51448 41064 51500 41070
rect 51448 41006 51500 41012
rect 50672 40468 50752 40474
rect 50620 40462 50752 40468
rect 50632 40446 50752 40462
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 50632 37806 50660 40446
rect 51172 39976 51224 39982
rect 51172 39918 51224 39924
rect 50712 39908 50764 39914
rect 50712 39850 50764 39856
rect 50724 38962 50752 39850
rect 51184 39098 51212 39918
rect 51172 39092 51224 39098
rect 51172 39034 51224 39040
rect 50712 38956 50764 38962
rect 50712 38898 50764 38904
rect 51184 38894 51212 39034
rect 51172 38888 51224 38894
rect 51172 38830 51224 38836
rect 50710 38584 50766 38593
rect 50710 38519 50712 38528
rect 50764 38519 50766 38528
rect 50712 38490 50764 38496
rect 50620 37800 50672 37806
rect 50620 37742 50672 37748
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 50160 36712 50212 36718
rect 50160 36654 50212 36660
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 50632 35562 50660 37742
rect 51184 37330 51212 38830
rect 51460 38654 51488 41006
rect 51908 40656 51960 40662
rect 51908 40598 51960 40604
rect 51816 40520 51868 40526
rect 51816 40462 51868 40468
rect 51828 39982 51856 40462
rect 51920 40186 51948 40598
rect 52472 40594 52500 41482
rect 52460 40588 52512 40594
rect 52460 40530 52512 40536
rect 51908 40180 51960 40186
rect 51908 40122 51960 40128
rect 51540 39976 51592 39982
rect 51540 39918 51592 39924
rect 51816 39976 51868 39982
rect 51816 39918 51868 39924
rect 52368 39976 52420 39982
rect 52368 39918 52420 39924
rect 51552 39574 51580 39918
rect 52380 39642 52408 39918
rect 52564 39794 52592 42078
rect 52828 42084 52880 42090
rect 52828 42026 52880 42032
rect 52472 39766 52592 39794
rect 52368 39636 52420 39642
rect 52368 39578 52420 39584
rect 51540 39568 51592 39574
rect 51540 39510 51592 39516
rect 52368 39432 52420 39438
rect 52368 39374 52420 39380
rect 51908 39364 51960 39370
rect 51908 39306 51960 39312
rect 51920 38894 51948 39306
rect 52380 39098 52408 39374
rect 52368 39092 52420 39098
rect 52368 39034 52420 39040
rect 52472 38978 52500 39766
rect 52564 39506 52684 39522
rect 52552 39500 52684 39506
rect 52604 39494 52684 39500
rect 52552 39442 52604 39448
rect 52656 39098 52684 39494
rect 52736 39500 52788 39506
rect 52840 39488 52868 42026
rect 52788 39460 52868 39488
rect 52736 39442 52788 39448
rect 52644 39092 52696 39098
rect 52644 39034 52696 39040
rect 52550 38992 52606 39001
rect 52472 38950 52550 38978
rect 52550 38927 52552 38936
rect 52604 38927 52606 38936
rect 52644 38956 52696 38962
rect 52552 38898 52604 38904
rect 52644 38898 52696 38904
rect 51908 38888 51960 38894
rect 51908 38830 51960 38836
rect 52460 38888 52512 38894
rect 52460 38830 52512 38836
rect 52000 38752 52052 38758
rect 52000 38694 52052 38700
rect 51368 38626 51488 38654
rect 51368 37806 51396 38626
rect 52012 38418 52040 38694
rect 52472 38457 52500 38830
rect 52552 38480 52604 38486
rect 52458 38448 52514 38457
rect 52000 38412 52052 38418
rect 52552 38422 52604 38428
rect 52458 38383 52514 38392
rect 52000 38354 52052 38360
rect 51356 37800 51408 37806
rect 51356 37742 51408 37748
rect 51172 37324 51224 37330
rect 51172 37266 51224 37272
rect 51080 36576 51132 36582
rect 51080 36518 51132 36524
rect 50896 35624 50948 35630
rect 50896 35566 50948 35572
rect 50620 35556 50672 35562
rect 50620 35498 50672 35504
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 49882 35184 49938 35193
rect 49700 35148 49752 35154
rect 49882 35119 49884 35128
rect 49700 35090 49752 35096
rect 49936 35119 49938 35128
rect 49884 35090 49936 35096
rect 50068 35080 50120 35086
rect 50068 35022 50120 35028
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 50080 34066 50108 35022
rect 50344 35012 50396 35018
rect 50344 34954 50396 34960
rect 50160 34944 50212 34950
rect 50160 34886 50212 34892
rect 50172 34746 50200 34886
rect 50160 34740 50212 34746
rect 50160 34682 50212 34688
rect 50068 34060 50120 34066
rect 50068 34002 50120 34008
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 50080 33454 50108 34002
rect 50068 33448 50120 33454
rect 50068 33390 50120 33396
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 49700 32972 49752 32978
rect 49700 32914 49752 32920
rect 49516 32836 49568 32842
rect 49516 32778 49568 32784
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 48320 31884 48372 31890
rect 48320 31826 48372 31832
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 47860 30184 47912 30190
rect 47860 30126 47912 30132
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 47872 29102 47900 30126
rect 48332 29306 48360 31826
rect 48872 31272 48924 31278
rect 48872 31214 48924 31220
rect 48780 30252 48832 30258
rect 48780 30194 48832 30200
rect 48320 29300 48372 29306
rect 48320 29242 48372 29248
rect 47860 29096 47912 29102
rect 47860 29038 47912 29044
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 47872 28762 47900 29038
rect 47860 28756 47912 28762
rect 47860 28698 47912 28704
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 48332 27538 48360 29242
rect 48792 28422 48820 30194
rect 48884 30054 48912 31214
rect 49056 30864 49108 30870
rect 49056 30806 49108 30812
rect 49068 30394 49096 30806
rect 49056 30388 49108 30394
rect 49056 30330 49108 30336
rect 48872 30048 48924 30054
rect 48872 29990 48924 29996
rect 48964 30048 49016 30054
rect 48964 29990 49016 29996
rect 48884 28558 48912 29990
rect 48976 29714 49004 29990
rect 48964 29708 49016 29714
rect 48964 29650 49016 29656
rect 49068 29102 49096 30330
rect 49528 30258 49556 32778
rect 49712 32745 49740 32914
rect 49698 32736 49754 32745
rect 49698 32671 49754 32680
rect 50172 31754 50200 34682
rect 50356 34649 50384 34954
rect 50908 34746 50936 35566
rect 50896 34740 50948 34746
rect 50896 34682 50948 34688
rect 50342 34640 50398 34649
rect 50342 34575 50398 34584
rect 50618 34504 50674 34513
rect 50908 34490 50936 34682
rect 50988 34536 51040 34542
rect 50908 34484 50988 34490
rect 50908 34478 51040 34484
rect 50618 34439 50674 34448
rect 50804 34468 50856 34474
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 50632 34202 50660 34439
rect 50804 34410 50856 34416
rect 50908 34462 51028 34478
rect 51092 34474 51120 36518
rect 51184 35698 51212 37266
rect 51368 37126 51396 37742
rect 51908 37324 51960 37330
rect 51908 37266 51960 37272
rect 52092 37324 52144 37330
rect 52092 37266 52144 37272
rect 52460 37324 52512 37330
rect 52460 37266 52512 37272
rect 51356 37120 51408 37126
rect 51920 37097 51948 37266
rect 52000 37188 52052 37194
rect 52000 37130 52052 37136
rect 51356 37062 51408 37068
rect 51906 37088 51962 37097
rect 51368 36650 51396 37062
rect 51906 37023 51962 37032
rect 51356 36644 51408 36650
rect 51356 36586 51408 36592
rect 51264 36236 51316 36242
rect 51264 36178 51316 36184
rect 51172 35692 51224 35698
rect 51172 35634 51224 35640
rect 51184 35154 51212 35634
rect 51276 35494 51304 36178
rect 51264 35488 51316 35494
rect 51264 35430 51316 35436
rect 51172 35148 51224 35154
rect 51172 35090 51224 35096
rect 51080 34468 51132 34474
rect 50712 34400 50764 34406
rect 50712 34342 50764 34348
rect 50620 34196 50672 34202
rect 50620 34138 50672 34144
rect 50724 33658 50752 34342
rect 50816 34105 50844 34410
rect 50802 34096 50858 34105
rect 50802 34031 50858 34040
rect 50712 33652 50764 33658
rect 50712 33594 50764 33600
rect 50712 33448 50764 33454
rect 50712 33390 50764 33396
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 50724 32230 50752 33390
rect 50712 32224 50764 32230
rect 50712 32166 50764 32172
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 50080 31726 50200 31754
rect 49516 30252 49568 30258
rect 49516 30194 49568 30200
rect 49424 30116 49476 30122
rect 49424 30058 49476 30064
rect 49884 30116 49936 30122
rect 49884 30058 49936 30064
rect 49436 29850 49464 30058
rect 49424 29844 49476 29850
rect 49424 29786 49476 29792
rect 49896 29306 49924 30058
rect 49976 29640 50028 29646
rect 49976 29582 50028 29588
rect 49988 29306 50016 29582
rect 49884 29300 49936 29306
rect 49884 29242 49936 29248
rect 49976 29300 50028 29306
rect 49976 29242 50028 29248
rect 49514 29200 49570 29209
rect 49514 29135 49516 29144
rect 49568 29135 49570 29144
rect 49516 29106 49568 29112
rect 49056 29096 49108 29102
rect 49056 29038 49108 29044
rect 49068 28626 49096 29038
rect 49240 28960 49292 28966
rect 49240 28902 49292 28908
rect 49252 28626 49280 28902
rect 49424 28756 49476 28762
rect 49424 28698 49476 28704
rect 49056 28620 49108 28626
rect 49056 28562 49108 28568
rect 49240 28620 49292 28626
rect 49240 28562 49292 28568
rect 48872 28552 48924 28558
rect 48872 28494 48924 28500
rect 48780 28416 48832 28422
rect 48780 28358 48832 28364
rect 48792 28014 48820 28358
rect 48780 28008 48832 28014
rect 48780 27950 48832 27956
rect 49068 27538 49096 28562
rect 49240 27872 49292 27878
rect 49240 27814 49292 27820
rect 48320 27532 48372 27538
rect 48320 27474 48372 27480
rect 49056 27532 49108 27538
rect 49056 27474 49108 27480
rect 48412 27328 48464 27334
rect 48412 27270 48464 27276
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 48424 26489 48452 27270
rect 48410 26480 48466 26489
rect 48410 26415 48466 26424
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 46204 26036 46256 26042
rect 46204 25978 46256 25984
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 46216 25430 46244 25978
rect 46204 25424 46256 25430
rect 46204 25366 46256 25372
rect 49068 25362 49096 27474
rect 49252 26926 49280 27814
rect 49240 26920 49292 26926
rect 49240 26862 49292 26868
rect 49252 26042 49280 26862
rect 49436 26246 49464 28698
rect 49988 28626 50016 29242
rect 49700 28620 49752 28626
rect 49700 28562 49752 28568
rect 49976 28620 50028 28626
rect 49976 28562 50028 28568
rect 49712 27674 49740 28562
rect 49700 27668 49752 27674
rect 49700 27610 49752 27616
rect 49884 27668 49936 27674
rect 49884 27610 49936 27616
rect 49608 27328 49660 27334
rect 49608 27270 49660 27276
rect 49424 26240 49476 26246
rect 49424 26182 49476 26188
rect 49240 26036 49292 26042
rect 49240 25978 49292 25984
rect 49056 25356 49108 25362
rect 49056 25298 49108 25304
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 49332 22094 49384 22098
rect 49436 22094 49464 26182
rect 49620 25401 49648 27270
rect 49896 27130 49924 27610
rect 49976 27532 50028 27538
rect 49976 27474 50028 27480
rect 49884 27124 49936 27130
rect 49884 27066 49936 27072
rect 49988 26450 50016 27474
rect 49976 26444 50028 26450
rect 49976 26386 50028 26392
rect 49606 25392 49662 25401
rect 49606 25327 49662 25336
rect 49988 24614 50016 26386
rect 50080 24682 50108 31726
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 50710 30968 50766 30977
rect 50710 30903 50712 30912
rect 50764 30903 50766 30912
rect 50712 30874 50764 30880
rect 50526 30832 50582 30841
rect 50526 30767 50528 30776
rect 50580 30767 50582 30776
rect 50620 30796 50672 30802
rect 50528 30738 50580 30744
rect 50620 30738 50672 30744
rect 50632 30054 50660 30738
rect 50160 30048 50212 30054
rect 50160 29990 50212 29996
rect 50620 30048 50672 30054
rect 50620 29990 50672 29996
rect 50172 27538 50200 29990
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50436 29640 50488 29646
rect 50436 29582 50488 29588
rect 50448 29306 50476 29582
rect 50436 29300 50488 29306
rect 50436 29242 50488 29248
rect 50620 29232 50672 29238
rect 50620 29174 50672 29180
rect 50300 28860 50596 28880
rect 50356 28858 50380 28860
rect 50436 28858 50460 28860
rect 50516 28858 50540 28860
rect 50378 28806 50380 28858
rect 50442 28806 50454 28858
rect 50516 28806 50518 28858
rect 50356 28804 50380 28806
rect 50436 28804 50460 28806
rect 50516 28804 50540 28806
rect 50300 28784 50596 28804
rect 50632 28626 50660 29174
rect 50712 29164 50764 29170
rect 50712 29106 50764 29112
rect 50724 28665 50752 29106
rect 50710 28656 50766 28665
rect 50620 28620 50672 28626
rect 50710 28591 50766 28600
rect 50620 28562 50672 28568
rect 50632 28218 50660 28562
rect 50620 28212 50672 28218
rect 50620 28154 50672 28160
rect 50724 28014 50752 28591
rect 50712 28008 50764 28014
rect 50712 27950 50764 27956
rect 50300 27772 50596 27792
rect 50356 27770 50380 27772
rect 50436 27770 50460 27772
rect 50516 27770 50540 27772
rect 50378 27718 50380 27770
rect 50442 27718 50454 27770
rect 50516 27718 50518 27770
rect 50356 27716 50380 27718
rect 50436 27716 50460 27718
rect 50516 27716 50540 27718
rect 50300 27696 50596 27716
rect 50252 27600 50304 27606
rect 50250 27568 50252 27577
rect 50304 27568 50306 27577
rect 50160 27532 50212 27538
rect 50250 27503 50306 27512
rect 50160 27474 50212 27480
rect 50816 26874 50844 34031
rect 50908 33522 50936 34462
rect 51080 34410 51132 34416
rect 50896 33516 50948 33522
rect 50896 33458 50948 33464
rect 51276 31754 51304 35430
rect 51368 35000 51396 36586
rect 52012 36310 52040 37130
rect 52104 36854 52132 37266
rect 52368 37256 52420 37262
rect 52368 37198 52420 37204
rect 52092 36848 52144 36854
rect 52092 36790 52144 36796
rect 52000 36304 52052 36310
rect 52000 36246 52052 36252
rect 52380 36174 52408 37198
rect 52472 36922 52500 37266
rect 52460 36916 52512 36922
rect 52460 36858 52512 36864
rect 52564 36378 52592 38422
rect 52656 38418 52684 38898
rect 52644 38412 52696 38418
rect 52644 38354 52696 38360
rect 52656 37097 52684 38354
rect 52642 37088 52698 37097
rect 52642 37023 52698 37032
rect 52656 36582 52684 37023
rect 52748 36718 52776 39442
rect 52828 38548 52880 38554
rect 52932 38536 52960 42094
rect 53208 41682 53236 43794
rect 53932 43648 53984 43654
rect 53932 43590 53984 43596
rect 53840 43240 53892 43246
rect 53840 43182 53892 43188
rect 53852 42702 53880 43182
rect 53944 42770 53972 43590
rect 54128 43314 54156 43794
rect 54208 43716 54260 43722
rect 54208 43658 54260 43664
rect 54220 43382 54248 43658
rect 54208 43376 54260 43382
rect 54208 43318 54260 43324
rect 54116 43308 54168 43314
rect 54116 43250 54168 43256
rect 54208 43240 54260 43246
rect 54208 43182 54260 43188
rect 54024 43172 54076 43178
rect 54024 43114 54076 43120
rect 53932 42764 53984 42770
rect 53932 42706 53984 42712
rect 53840 42696 53892 42702
rect 53840 42638 53892 42644
rect 54036 42158 54064 43114
rect 54220 42838 54248 43182
rect 54496 43178 54524 44270
rect 54772 43625 54800 46446
rect 55048 46170 55076 46514
rect 55036 46164 55088 46170
rect 55036 46106 55088 46112
rect 54944 46028 54996 46034
rect 54944 45970 54996 45976
rect 54956 45422 54984 45970
rect 55036 45960 55088 45966
rect 55036 45902 55088 45908
rect 54944 45416 54996 45422
rect 54944 45358 54996 45364
rect 55048 45121 55076 45902
rect 55128 45416 55180 45422
rect 55128 45358 55180 45364
rect 55034 45112 55090 45121
rect 55034 45047 55090 45056
rect 55140 44962 55168 45358
rect 55048 44934 55168 44962
rect 54944 44736 54996 44742
rect 54944 44678 54996 44684
rect 54956 43926 54984 44678
rect 54944 43920 54996 43926
rect 54944 43862 54996 43868
rect 54852 43784 54904 43790
rect 54852 43726 54904 43732
rect 54758 43616 54814 43625
rect 54758 43551 54814 43560
rect 54484 43172 54536 43178
rect 54484 43114 54536 43120
rect 54208 42832 54260 42838
rect 54208 42774 54260 42780
rect 54116 42560 54168 42566
rect 54116 42502 54168 42508
rect 54128 42158 54156 42502
rect 54220 42362 54248 42774
rect 54208 42356 54260 42362
rect 54208 42298 54260 42304
rect 54864 42158 54892 43726
rect 55048 43382 55076 44934
rect 55128 44260 55180 44266
rect 55128 44202 55180 44208
rect 55140 43994 55168 44202
rect 55128 43988 55180 43994
rect 55128 43930 55180 43936
rect 55036 43376 55088 43382
rect 55036 43318 55088 43324
rect 54944 43308 54996 43314
rect 54944 43250 54996 43256
rect 54956 42752 54984 43250
rect 55128 43240 55180 43246
rect 55128 43182 55180 43188
rect 55036 42764 55088 42770
rect 54956 42724 55036 42752
rect 55036 42706 55088 42712
rect 55048 42634 55076 42706
rect 55036 42628 55088 42634
rect 55036 42570 55088 42576
rect 55048 42226 55076 42570
rect 55140 42566 55168 43182
rect 55128 42560 55180 42566
rect 55128 42502 55180 42508
rect 55036 42220 55088 42226
rect 55036 42162 55088 42168
rect 54024 42152 54076 42158
rect 54024 42094 54076 42100
rect 54116 42152 54168 42158
rect 54116 42094 54168 42100
rect 54852 42152 54904 42158
rect 54852 42094 54904 42100
rect 54036 41970 54064 42094
rect 54036 41942 54156 41970
rect 53196 41676 53248 41682
rect 53196 41618 53248 41624
rect 53380 41676 53432 41682
rect 53380 41618 53432 41624
rect 53932 41676 53984 41682
rect 53932 41618 53984 41624
rect 53392 41274 53420 41618
rect 53840 41608 53892 41614
rect 53840 41550 53892 41556
rect 53852 41274 53880 41550
rect 53380 41268 53432 41274
rect 53380 41210 53432 41216
rect 53840 41268 53892 41274
rect 53840 41210 53892 41216
rect 53840 40928 53892 40934
rect 53840 40870 53892 40876
rect 53852 40594 53880 40870
rect 53472 40588 53524 40594
rect 53472 40530 53524 40536
rect 53840 40588 53892 40594
rect 53840 40530 53892 40536
rect 53104 40384 53156 40390
rect 53104 40326 53156 40332
rect 53012 39636 53064 39642
rect 53012 39578 53064 39584
rect 53024 39506 53052 39578
rect 53012 39500 53064 39506
rect 53012 39442 53064 39448
rect 53012 38888 53064 38894
rect 53012 38830 53064 38836
rect 52880 38508 52960 38536
rect 52828 38490 52880 38496
rect 53024 38010 53052 38830
rect 53116 38350 53144 40326
rect 53286 38992 53342 39001
rect 53196 38956 53248 38962
rect 53286 38927 53288 38936
rect 53196 38898 53248 38904
rect 53340 38927 53342 38936
rect 53288 38898 53340 38904
rect 53208 38758 53236 38898
rect 53196 38752 53248 38758
rect 53196 38694 53248 38700
rect 53208 38486 53236 38694
rect 53196 38480 53248 38486
rect 53196 38422 53248 38428
rect 53378 38448 53434 38457
rect 53378 38383 53434 38392
rect 53392 38350 53420 38383
rect 53104 38344 53156 38350
rect 53104 38286 53156 38292
rect 53380 38344 53432 38350
rect 53380 38286 53432 38292
rect 53012 38004 53064 38010
rect 53012 37946 53064 37952
rect 53392 37274 53420 38286
rect 53484 38010 53512 40530
rect 53564 40520 53616 40526
rect 53564 40462 53616 40468
rect 53576 39846 53604 40462
rect 53852 39982 53880 40530
rect 53944 40526 53972 41618
rect 54024 41540 54076 41546
rect 54024 41482 54076 41488
rect 54036 40934 54064 41482
rect 54128 41070 54156 41942
rect 54864 41682 54892 42094
rect 54852 41676 54904 41682
rect 54852 41618 54904 41624
rect 54864 41562 54892 41618
rect 54864 41534 55168 41562
rect 54852 41472 54904 41478
rect 54852 41414 54904 41420
rect 54864 41070 54892 41414
rect 54116 41064 54168 41070
rect 54116 41006 54168 41012
rect 54668 41064 54720 41070
rect 54668 41006 54720 41012
rect 54852 41064 54904 41070
rect 54852 41006 54904 41012
rect 54024 40928 54076 40934
rect 54024 40870 54076 40876
rect 54680 40712 54708 41006
rect 54680 40684 54892 40712
rect 53932 40520 53984 40526
rect 53932 40462 53984 40468
rect 54300 40520 54352 40526
rect 54300 40462 54352 40468
rect 54024 40452 54076 40458
rect 54024 40394 54076 40400
rect 54036 40118 54064 40394
rect 54024 40112 54076 40118
rect 54024 40054 54076 40060
rect 54312 39982 54340 40462
rect 54864 40050 54892 40684
rect 55140 40594 55168 41534
rect 55220 40656 55272 40662
rect 55220 40598 55272 40604
rect 55128 40588 55180 40594
rect 55128 40530 55180 40536
rect 55036 40452 55088 40458
rect 55036 40394 55088 40400
rect 54852 40044 54904 40050
rect 54852 39986 54904 39992
rect 53748 39976 53800 39982
rect 53748 39918 53800 39924
rect 53840 39976 53892 39982
rect 53840 39918 53892 39924
rect 54300 39976 54352 39982
rect 54300 39918 54352 39924
rect 54484 39976 54536 39982
rect 54484 39918 54536 39924
rect 53760 39846 53788 39918
rect 54496 39846 54524 39918
rect 53564 39840 53616 39846
rect 53564 39782 53616 39788
rect 53748 39840 53800 39846
rect 53748 39782 53800 39788
rect 54484 39840 54536 39846
rect 54484 39782 54536 39788
rect 53576 38894 53604 39782
rect 54864 39642 54892 39986
rect 55048 39982 55076 40394
rect 55036 39976 55088 39982
rect 55036 39918 55088 39924
rect 53840 39636 53892 39642
rect 53840 39578 53892 39584
rect 54852 39636 54904 39642
rect 54852 39578 54904 39584
rect 53748 39432 53800 39438
rect 53852 39386 53880 39578
rect 53800 39380 53880 39386
rect 53748 39374 53880 39380
rect 53760 39358 53880 39374
rect 53564 38888 53616 38894
rect 53564 38830 53616 38836
rect 54116 38752 54168 38758
rect 54116 38694 54168 38700
rect 54128 38554 54156 38694
rect 54206 38584 54262 38593
rect 54116 38548 54168 38554
rect 54206 38519 54208 38528
rect 54116 38490 54168 38496
rect 54260 38519 54262 38528
rect 54208 38490 54260 38496
rect 54024 38412 54076 38418
rect 54024 38354 54076 38360
rect 54760 38412 54812 38418
rect 54760 38354 54812 38360
rect 53472 38004 53524 38010
rect 53472 37946 53524 37952
rect 53484 37806 53512 37946
rect 54036 37874 54064 38354
rect 54772 37874 54800 38354
rect 54024 37868 54076 37874
rect 54024 37810 54076 37816
rect 54760 37868 54812 37874
rect 54760 37810 54812 37816
rect 53472 37800 53524 37806
rect 53472 37742 53524 37748
rect 54668 37800 54720 37806
rect 54668 37742 54720 37748
rect 54680 37398 54708 37742
rect 54668 37392 54720 37398
rect 54668 37334 54720 37340
rect 54772 37330 54800 37810
rect 54864 37806 54892 39578
rect 55036 39364 55088 39370
rect 55036 39306 55088 39312
rect 55048 38894 55076 39306
rect 55036 38888 55088 38894
rect 55036 38830 55088 38836
rect 54852 37800 54904 37806
rect 54852 37742 54904 37748
rect 54576 37324 54628 37330
rect 53392 37246 53788 37274
rect 54576 37266 54628 37272
rect 54760 37324 54812 37330
rect 54760 37266 54812 37272
rect 53760 36854 53788 37246
rect 53840 37256 53892 37262
rect 53840 37198 53892 37204
rect 53852 36922 53880 37198
rect 54588 37126 54616 37266
rect 54024 37120 54076 37126
rect 54024 37062 54076 37068
rect 54576 37120 54628 37126
rect 54576 37062 54628 37068
rect 53840 36916 53892 36922
rect 53840 36858 53892 36864
rect 53748 36848 53800 36854
rect 53748 36790 53800 36796
rect 52736 36712 52788 36718
rect 52736 36654 52788 36660
rect 53012 36712 53064 36718
rect 53012 36654 53064 36660
rect 52644 36576 52696 36582
rect 52644 36518 52696 36524
rect 52656 36378 52684 36518
rect 52552 36372 52604 36378
rect 52552 36314 52604 36320
rect 52644 36372 52696 36378
rect 52644 36314 52696 36320
rect 52368 36168 52420 36174
rect 52368 36110 52420 36116
rect 52748 36038 52776 36654
rect 53024 36310 53052 36654
rect 53012 36304 53064 36310
rect 53012 36246 53064 36252
rect 52828 36168 52880 36174
rect 52828 36110 52880 36116
rect 52840 36038 52868 36110
rect 52736 36032 52788 36038
rect 52736 35974 52788 35980
rect 52828 36032 52880 36038
rect 52828 35974 52880 35980
rect 51724 35624 51776 35630
rect 51724 35566 51776 35572
rect 52092 35624 52144 35630
rect 52092 35566 52144 35572
rect 53104 35624 53156 35630
rect 53104 35566 53156 35572
rect 51448 35012 51500 35018
rect 51368 34972 51448 35000
rect 51448 34954 51500 34960
rect 51356 33312 51408 33318
rect 51356 33254 51408 33260
rect 51184 31726 51304 31754
rect 51184 31210 51212 31726
rect 51264 31476 51316 31482
rect 51264 31418 51316 31424
rect 51172 31204 51224 31210
rect 51172 31146 51224 31152
rect 51276 30598 51304 31418
rect 51264 30592 51316 30598
rect 51264 30534 51316 30540
rect 50896 30048 50948 30054
rect 50896 29990 50948 29996
rect 50908 29714 50936 29990
rect 51264 29776 51316 29782
rect 51264 29718 51316 29724
rect 50896 29708 50948 29714
rect 50896 29650 50948 29656
rect 50908 29102 50936 29650
rect 51000 29158 51120 29186
rect 50896 29096 50948 29102
rect 50896 29038 50948 29044
rect 51000 28966 51028 29158
rect 51092 29050 51120 29158
rect 51092 29034 51212 29050
rect 51092 29028 51224 29034
rect 51092 29022 51172 29028
rect 51172 28970 51224 28976
rect 50988 28960 51040 28966
rect 50988 28902 51040 28908
rect 51080 28008 51132 28014
rect 51080 27950 51132 27956
rect 50988 26920 51040 26926
rect 50816 26846 50936 26874
rect 50988 26862 51040 26868
rect 50620 26784 50672 26790
rect 50620 26726 50672 26732
rect 50300 26684 50596 26704
rect 50356 26682 50380 26684
rect 50436 26682 50460 26684
rect 50516 26682 50540 26684
rect 50378 26630 50380 26682
rect 50442 26630 50454 26682
rect 50516 26630 50518 26682
rect 50356 26628 50380 26630
rect 50436 26628 50460 26630
rect 50516 26628 50540 26630
rect 50300 26608 50596 26628
rect 50632 26450 50660 26726
rect 50620 26444 50672 26450
rect 50620 26386 50672 26392
rect 50160 26376 50212 26382
rect 50160 26318 50212 26324
rect 50172 25838 50200 26318
rect 50620 26036 50672 26042
rect 50620 25978 50672 25984
rect 50632 25838 50660 25978
rect 50160 25832 50212 25838
rect 50160 25774 50212 25780
rect 50620 25832 50672 25838
rect 50620 25774 50672 25780
rect 50300 25596 50596 25616
rect 50356 25594 50380 25596
rect 50436 25594 50460 25596
rect 50516 25594 50540 25596
rect 50378 25542 50380 25594
rect 50442 25542 50454 25594
rect 50516 25542 50518 25594
rect 50356 25540 50380 25542
rect 50436 25540 50460 25542
rect 50516 25540 50540 25542
rect 50300 25520 50596 25540
rect 50632 24750 50660 25774
rect 50804 24948 50856 24954
rect 50804 24890 50856 24896
rect 50160 24744 50212 24750
rect 50160 24686 50212 24692
rect 50620 24744 50672 24750
rect 50620 24686 50672 24692
rect 50068 24676 50120 24682
rect 50068 24618 50120 24624
rect 49976 24608 50028 24614
rect 49976 24550 50028 24556
rect 50172 23730 50200 24686
rect 50300 24508 50596 24528
rect 50356 24506 50380 24508
rect 50436 24506 50460 24508
rect 50516 24506 50540 24508
rect 50378 24454 50380 24506
rect 50442 24454 50454 24506
rect 50516 24454 50518 24506
rect 50356 24452 50380 24454
rect 50436 24452 50460 24454
rect 50516 24452 50540 24454
rect 50300 24432 50596 24452
rect 50816 23866 50844 24890
rect 50804 23860 50856 23866
rect 50804 23802 50856 23808
rect 50160 23724 50212 23730
rect 50160 23666 50212 23672
rect 50804 23724 50856 23730
rect 50804 23666 50856 23672
rect 50712 23656 50764 23662
rect 50712 23598 50764 23604
rect 50724 23526 50752 23598
rect 49884 23520 49936 23526
rect 49884 23462 49936 23468
rect 50712 23520 50764 23526
rect 50712 23462 50764 23468
rect 49896 23322 49924 23462
rect 50300 23420 50596 23440
rect 50356 23418 50380 23420
rect 50436 23418 50460 23420
rect 50516 23418 50540 23420
rect 50378 23366 50380 23418
rect 50442 23366 50454 23418
rect 50516 23366 50518 23418
rect 50356 23364 50380 23366
rect 50436 23364 50460 23366
rect 50516 23364 50540 23366
rect 50300 23344 50596 23364
rect 49884 23316 49936 23322
rect 49884 23258 49936 23264
rect 50436 23248 50488 23254
rect 50434 23216 50436 23225
rect 50488 23216 50490 23225
rect 49884 23180 49936 23186
rect 50434 23151 50490 23160
rect 49884 23122 49936 23128
rect 49792 22976 49844 22982
rect 49792 22918 49844 22924
rect 49332 22092 49464 22094
rect 49384 22066 49464 22092
rect 49332 22034 49384 22040
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 49056 21888 49108 21894
rect 49056 21830 49108 21836
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 5092 12782 5120 13126
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11286 4108 11630
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 3700 8560 3752 8566
rect 3700 8502 3752 8508
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1872 7546 1900 8298
rect 2056 7993 2084 8298
rect 3160 8022 3188 8366
rect 3148 8016 3200 8022
rect 2042 7984 2098 7993
rect 3148 7958 3200 7964
rect 2042 7919 2098 7928
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1964 7041 1992 7686
rect 1950 7032 2006 7041
rect 2332 7002 2360 7890
rect 2792 7750 2820 7890
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 1950 6967 2006 6976
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2516 6458 2544 6734
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2792 6254 2820 7686
rect 3160 7342 3188 7686
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 1952 6112 2004 6118
rect 1950 6080 1952 6089
rect 2004 6080 2006 6089
rect 1950 6015 2006 6024
rect 2332 5914 2360 6122
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2792 5846 2820 6190
rect 2780 5840 2832 5846
rect 2780 5782 2832 5788
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2780 5160 2832 5166
rect 2778 5128 2780 5137
rect 2832 5128 2834 5137
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2596 5092 2648 5098
rect 2778 5063 2834 5072
rect 2596 5034 2648 5040
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1412 800 1440 3878
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1688 3058 1716 3606
rect 2332 3466 2360 5034
rect 2608 4826 2636 5034
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2596 4820 2648 4826
rect 2596 4762 2648 4768
rect 2792 4690 2820 4966
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2884 4434 2912 5170
rect 2792 4406 2912 4434
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 2424 1850 2452 3402
rect 2792 3233 2820 4406
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2884 4185 2912 4218
rect 2870 4176 2926 4185
rect 2870 4111 2926 4120
rect 2976 4026 3004 5170
rect 3344 4622 3372 6190
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3436 5166 3464 5714
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3436 4690 3464 5102
rect 3424 4684 3476 4690
rect 3424 4626 3476 4632
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4146 3096 4422
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3712 4078 3740 8502
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 4632 4146 4660 4422
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 2884 3998 3004 4026
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 2884 3602 2912 3998
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2332 1822 2452 1850
rect 2332 800 2360 1822
rect 2884 1329 2912 3334
rect 2976 3058 3004 3878
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3160 3194 3188 3538
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3712 2990 3740 4014
rect 3976 3528 4028 3534
rect 4172 3482 4200 4014
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 31312 3602 31340 21830
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 49068 21010 49096 21830
rect 49804 21010 49832 22918
rect 49896 22574 49924 23122
rect 49976 23112 50028 23118
rect 49976 23054 50028 23060
rect 49884 22568 49936 22574
rect 49884 22510 49936 22516
rect 49896 21486 49924 22510
rect 49884 21480 49936 21486
rect 49884 21422 49936 21428
rect 49988 21434 50016 23054
rect 50724 22574 50752 23462
rect 50620 22568 50672 22574
rect 50620 22510 50672 22516
rect 50712 22568 50764 22574
rect 50712 22510 50764 22516
rect 50300 22332 50596 22352
rect 50356 22330 50380 22332
rect 50436 22330 50460 22332
rect 50516 22330 50540 22332
rect 50378 22278 50380 22330
rect 50442 22278 50454 22330
rect 50516 22278 50518 22330
rect 50356 22276 50380 22278
rect 50436 22276 50460 22278
rect 50516 22276 50540 22278
rect 50300 22256 50596 22276
rect 50632 22234 50660 22510
rect 50620 22228 50672 22234
rect 50620 22170 50672 22176
rect 50160 21480 50212 21486
rect 47860 21004 47912 21010
rect 47860 20946 47912 20952
rect 49056 21004 49108 21010
rect 49056 20946 49108 20952
rect 49792 21004 49844 21010
rect 49792 20946 49844 20952
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 47872 19310 47900 20946
rect 48412 20800 48464 20806
rect 48412 20742 48464 20748
rect 48424 19961 48452 20742
rect 48410 19952 48466 19961
rect 49068 19922 49096 20946
rect 48410 19887 48466 19896
rect 49056 19916 49108 19922
rect 49056 19858 49108 19864
rect 49056 19712 49108 19718
rect 49056 19654 49108 19660
rect 49068 19310 49096 19654
rect 49804 19310 49832 20946
rect 47860 19304 47912 19310
rect 47860 19246 47912 19252
rect 49056 19304 49108 19310
rect 49056 19246 49108 19252
rect 49792 19304 49844 19310
rect 49792 19246 49844 19252
rect 49068 18834 49096 19246
rect 49700 19168 49752 19174
rect 49700 19110 49752 19116
rect 49056 18828 49108 18834
rect 49056 18770 49108 18776
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 49712 17202 49740 19110
rect 49804 18086 49832 19246
rect 49896 18834 49924 21422
rect 49988 21406 50108 21434
rect 50160 21422 50212 21428
rect 49976 21344 50028 21350
rect 49976 21286 50028 21292
rect 49988 21146 50016 21286
rect 49976 21140 50028 21146
rect 49976 21082 50028 21088
rect 50080 20482 50108 21406
rect 49988 20454 50108 20482
rect 49988 19310 50016 20454
rect 50068 20392 50120 20398
rect 50068 20334 50120 20340
rect 50080 19854 50108 20334
rect 50068 19848 50120 19854
rect 50068 19790 50120 19796
rect 50068 19712 50120 19718
rect 50068 19654 50120 19660
rect 49976 19304 50028 19310
rect 49976 19246 50028 19252
rect 49988 18970 50016 19246
rect 49976 18964 50028 18970
rect 49976 18906 50028 18912
rect 49884 18828 49936 18834
rect 49884 18770 49936 18776
rect 49792 18080 49844 18086
rect 49792 18022 49844 18028
rect 49804 17746 49832 18022
rect 49792 17740 49844 17746
rect 49792 17682 49844 17688
rect 49700 17196 49752 17202
rect 49700 17138 49752 17144
rect 49712 17082 49740 17138
rect 49882 17096 49938 17105
rect 49712 17054 49832 17082
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 49698 15600 49754 15609
rect 49698 15535 49700 15544
rect 49752 15535 49754 15544
rect 49700 15506 49752 15512
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 49804 15026 49832 17054
rect 49882 17031 49938 17040
rect 49896 16794 49924 17031
rect 49884 16788 49936 16794
rect 49884 16730 49936 16736
rect 50080 16674 50108 19654
rect 50172 19174 50200 21422
rect 50620 21412 50672 21418
rect 50620 21354 50672 21360
rect 50300 21244 50596 21264
rect 50356 21242 50380 21244
rect 50436 21242 50460 21244
rect 50516 21242 50540 21244
rect 50378 21190 50380 21242
rect 50442 21190 50454 21242
rect 50516 21190 50518 21242
rect 50356 21188 50380 21190
rect 50436 21188 50460 21190
rect 50516 21188 50540 21190
rect 50300 21168 50596 21188
rect 50632 21078 50660 21354
rect 50620 21072 50672 21078
rect 50620 21014 50672 21020
rect 50724 20398 50752 22510
rect 50712 20392 50764 20398
rect 50712 20334 50764 20340
rect 50620 20256 50672 20262
rect 50620 20198 50672 20204
rect 50300 20156 50596 20176
rect 50356 20154 50380 20156
rect 50436 20154 50460 20156
rect 50516 20154 50540 20156
rect 50378 20102 50380 20154
rect 50442 20102 50454 20154
rect 50516 20102 50518 20154
rect 50356 20100 50380 20102
rect 50436 20100 50460 20102
rect 50516 20100 50540 20102
rect 50300 20080 50596 20100
rect 50632 19786 50660 20198
rect 50724 19922 50752 20334
rect 50712 19916 50764 19922
rect 50712 19858 50764 19864
rect 50620 19780 50672 19786
rect 50620 19722 50672 19728
rect 50712 19712 50764 19718
rect 50712 19654 50764 19660
rect 50160 19168 50212 19174
rect 50160 19110 50212 19116
rect 50300 19068 50596 19088
rect 50356 19066 50380 19068
rect 50436 19066 50460 19068
rect 50516 19066 50540 19068
rect 50378 19014 50380 19066
rect 50442 19014 50454 19066
rect 50516 19014 50518 19066
rect 50356 19012 50380 19014
rect 50436 19012 50460 19014
rect 50516 19012 50540 19014
rect 50300 18992 50596 19012
rect 50724 18970 50752 19654
rect 50712 18964 50764 18970
rect 50712 18906 50764 18912
rect 50618 18864 50674 18873
rect 50618 18799 50674 18808
rect 50632 18766 50660 18799
rect 50620 18760 50672 18766
rect 50620 18702 50672 18708
rect 50158 18456 50214 18465
rect 50158 18391 50214 18400
rect 50172 18222 50200 18391
rect 50160 18216 50212 18222
rect 50160 18158 50212 18164
rect 50300 17980 50596 18000
rect 50356 17978 50380 17980
rect 50436 17978 50460 17980
rect 50516 17978 50540 17980
rect 50378 17926 50380 17978
rect 50442 17926 50454 17978
rect 50516 17926 50518 17978
rect 50356 17924 50380 17926
rect 50436 17924 50460 17926
rect 50516 17924 50540 17926
rect 50300 17904 50596 17924
rect 50528 17740 50580 17746
rect 50528 17682 50580 17688
rect 50540 17377 50568 17682
rect 50526 17368 50582 17377
rect 50526 17303 50582 17312
rect 50160 17060 50212 17066
rect 50160 17002 50212 17008
rect 50172 16794 50200 17002
rect 50300 16892 50596 16912
rect 50356 16890 50380 16892
rect 50436 16890 50460 16892
rect 50516 16890 50540 16892
rect 50378 16838 50380 16890
rect 50442 16838 50454 16890
rect 50516 16838 50518 16890
rect 50356 16836 50380 16838
rect 50436 16836 50460 16838
rect 50516 16836 50540 16838
rect 50300 16816 50596 16836
rect 50160 16788 50212 16794
rect 50160 16730 50212 16736
rect 49976 16652 50028 16658
rect 50080 16646 50200 16674
rect 49976 16594 50028 16600
rect 49988 15910 50016 16594
rect 49976 15904 50028 15910
rect 49976 15846 50028 15852
rect 49792 15020 49844 15026
rect 49792 14962 49844 14968
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 49146 14104 49202 14113
rect 49146 14039 49202 14048
rect 49700 14068 49752 14074
rect 49160 13870 49188 14039
rect 49700 14010 49752 14016
rect 49148 13864 49200 13870
rect 49148 13806 49200 13812
rect 49424 13796 49476 13802
rect 49424 13738 49476 13744
rect 47492 13388 47544 13394
rect 47492 13330 47544 13336
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 47032 8424 47084 8430
rect 47032 8366 47084 8372
rect 46940 8288 46992 8294
rect 46940 8230 46992 8236
rect 46952 7954 46980 8230
rect 47044 8022 47072 8366
rect 47032 8016 47084 8022
rect 47032 7958 47084 7964
rect 46940 7948 46992 7954
rect 46940 7890 46992 7896
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 46572 7336 46624 7342
rect 46572 7278 46624 7284
rect 47216 7336 47268 7342
rect 47216 7278 47268 7284
rect 46584 7002 46612 7278
rect 46572 6996 46624 7002
rect 46572 6938 46624 6944
rect 45192 6860 45244 6866
rect 45192 6802 45244 6808
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 43812 5772 43864 5778
rect 43812 5714 43864 5720
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 43824 5302 43852 5714
rect 44640 5568 44692 5574
rect 44640 5510 44692 5516
rect 44916 5568 44968 5574
rect 44916 5510 44968 5516
rect 43812 5296 43864 5302
rect 43812 5238 43864 5244
rect 44088 5160 44140 5166
rect 44088 5102 44140 5108
rect 38108 4684 38160 4690
rect 38108 4626 38160 4632
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33968 4072 34020 4078
rect 33968 4014 34020 4020
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 31300 3596 31352 3602
rect 31300 3538 31352 3544
rect 33324 3596 33376 3602
rect 33324 3538 33376 3544
rect 3976 3470 4028 3476
rect 3988 3194 4016 3470
rect 4080 3454 4200 3482
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4080 3126 4108 3454
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2870 1320 2926 1329
rect 2870 1255 2926 1264
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2976 513 3004 2246
rect 3252 800 3280 2790
rect 3988 2650 4016 2858
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4172 2394 4200 2858
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4356 2446 4384 2790
rect 4632 2514 4660 3334
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4080 2366 4200 2394
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4080 2281 4108 2366
rect 4066 2272 4122 2281
rect 4066 2207 4122 2216
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4724 1578 4752 3062
rect 5092 2854 5120 3334
rect 5356 2984 5408 2990
rect 5408 2944 5580 2972
rect 5356 2926 5408 2932
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4172 1550 4752 1578
rect 4172 800 4200 1550
rect 5092 800 5120 2518
rect 5276 2446 5304 2790
rect 5552 2514 5580 2944
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5644 2514 5672 2858
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6104 800 6132 3538
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 7024 800 7052 2926
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 7944 800 7972 2450
rect 8864 800 8892 2926
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 19156 2508 19208 2514
rect 19156 2450 19208 2456
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 23848 2508 23900 2514
rect 23848 2450 23900 2456
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 26700 2508 26752 2514
rect 26700 2450 26752 2456
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 9784 800 9812 2450
rect 10796 800 10824 2450
rect 11716 800 11744 2450
rect 12636 800 12664 2450
rect 13556 800 13584 2450
rect 14476 800 14504 2450
rect 15488 800 15516 2450
rect 16408 800 16436 2450
rect 17328 800 17356 2450
rect 18248 800 18276 2450
rect 19168 800 19196 2450
rect 20088 800 20116 2450
rect 21100 800 21128 2450
rect 22020 800 22048 2450
rect 22940 800 22968 2450
rect 23860 800 23888 2450
rect 24780 800 24808 2450
rect 25792 800 25820 2450
rect 26712 800 26740 2450
rect 27632 800 27660 2450
rect 28552 800 28580 3538
rect 29472 800 29500 3538
rect 31116 3392 31168 3398
rect 31116 3334 31168 3340
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 30576 2582 30604 2790
rect 30564 2576 30616 2582
rect 30564 2518 30616 2524
rect 31128 2446 31156 3334
rect 31312 2990 31340 3538
rect 31392 3392 31444 3398
rect 31392 3334 31444 3340
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 33140 3392 33192 3398
rect 33140 3334 33192 3340
rect 33232 3392 33284 3398
rect 33232 3334 33284 3340
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31404 2514 31432 3334
rect 31944 2916 31996 2922
rect 31944 2858 31996 2864
rect 31392 2508 31444 2514
rect 31392 2450 31444 2456
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31956 2378 31984 2858
rect 32048 2514 32076 3334
rect 32312 2916 32364 2922
rect 32312 2858 32364 2864
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 32232 2514 32260 2790
rect 32036 2508 32088 2514
rect 32036 2450 32088 2456
rect 32220 2508 32272 2514
rect 32220 2450 32272 2456
rect 30472 2372 30524 2378
rect 30472 2314 30524 2320
rect 31944 2372 31996 2378
rect 31944 2314 31996 2320
rect 30484 800 30512 2314
rect 31392 2304 31444 2310
rect 31392 2246 31444 2252
rect 31404 800 31432 2246
rect 32324 800 32352 2858
rect 33152 2514 33180 3334
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 33244 800 33272 3334
rect 33336 2378 33364 3538
rect 33428 2990 33456 4014
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 33416 2984 33468 2990
rect 33416 2926 33468 2932
rect 33796 2514 33824 3878
rect 33980 3058 34008 4014
rect 34244 3596 34296 3602
rect 34244 3538 34296 3544
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 33968 3052 34020 3058
rect 33968 2994 34020 3000
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 33324 2372 33376 2378
rect 33324 2314 33376 2320
rect 34164 800 34192 3334
rect 34256 3194 34284 3538
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34532 2514 34560 4422
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34796 3936 34848 3942
rect 34796 3878 34848 3884
rect 35532 3936 35584 3942
rect 35532 3878 35584 3884
rect 34808 2514 34836 3878
rect 35256 3392 35308 3398
rect 35256 3334 35308 3340
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34520 2508 34572 2514
rect 34520 2450 34572 2456
rect 34796 2508 34848 2514
rect 34796 2450 34848 2456
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35268 1714 35296 3334
rect 35544 3058 35572 3878
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35532 3052 35584 3058
rect 35532 2994 35584 3000
rect 35820 2650 35848 3538
rect 35912 2990 35940 4422
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 35900 2984 35952 2990
rect 35900 2926 35952 2932
rect 36084 2848 36136 2854
rect 36084 2790 36136 2796
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 35084 1686 35296 1714
rect 35084 800 35112 1686
rect 36096 800 36124 2790
rect 36188 2514 36216 3878
rect 36176 2508 36228 2514
rect 36176 2450 36228 2456
rect 36280 2446 36308 4422
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37004 3392 37056 3398
rect 37004 3334 37056 3340
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 37016 800 37044 3334
rect 37108 2650 37136 3538
rect 37200 2990 37228 4082
rect 38120 4078 38148 4626
rect 38476 4480 38528 4486
rect 38476 4422 38528 4428
rect 38752 4480 38804 4486
rect 38752 4422 38804 4428
rect 42800 4480 42852 4486
rect 42800 4422 42852 4428
rect 43536 4480 43588 4486
rect 43536 4422 43588 4428
rect 37372 4072 37424 4078
rect 37372 4014 37424 4020
rect 38108 4072 38160 4078
rect 38108 4014 38160 4020
rect 37384 3194 37412 4014
rect 37924 3392 37976 3398
rect 37924 3334 37976 3340
rect 37372 3188 37424 3194
rect 37372 3130 37424 3136
rect 37188 2984 37240 2990
rect 37188 2926 37240 2932
rect 37384 2922 37412 3130
rect 37372 2916 37424 2922
rect 37372 2858 37424 2864
rect 37096 2644 37148 2650
rect 37096 2586 37148 2592
rect 37936 800 37964 3334
rect 38488 3058 38516 4422
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38672 3194 38700 3538
rect 38660 3188 38712 3194
rect 38660 3130 38712 3136
rect 38476 3052 38528 3058
rect 38476 2994 38528 3000
rect 38764 2514 38792 4422
rect 40040 4208 40092 4214
rect 40040 4150 40092 4156
rect 41604 4208 41656 4214
rect 41604 4150 41656 4156
rect 42708 4208 42760 4214
rect 42708 4150 42760 4156
rect 39120 4072 39172 4078
rect 39120 4014 39172 4020
rect 39028 3936 39080 3942
rect 39028 3878 39080 3884
rect 38936 3596 38988 3602
rect 38936 3538 38988 3544
rect 38844 3392 38896 3398
rect 38844 3334 38896 3340
rect 38752 2508 38804 2514
rect 38752 2450 38804 2456
rect 38856 800 38884 3334
rect 38948 2650 38976 3538
rect 38936 2644 38988 2650
rect 38936 2586 38988 2592
rect 39040 2514 39068 3878
rect 39132 2990 39160 4014
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39776 2990 39804 3538
rect 39120 2984 39172 2990
rect 39120 2926 39172 2932
rect 39764 2984 39816 2990
rect 39764 2926 39816 2932
rect 40052 2514 40080 4150
rect 40500 4072 40552 4078
rect 40500 4014 40552 4020
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 40236 2514 40264 3334
rect 40512 3058 40540 4014
rect 40500 3052 40552 3058
rect 40500 2994 40552 3000
rect 40776 2848 40828 2854
rect 40776 2790 40828 2796
rect 39028 2508 39080 2514
rect 39028 2450 39080 2456
rect 40040 2508 40092 2514
rect 40040 2450 40092 2456
rect 40224 2508 40276 2514
rect 40224 2450 40276 2456
rect 39764 2372 39816 2378
rect 39764 2314 39816 2320
rect 39776 800 39804 2314
rect 40788 800 40816 2790
rect 41616 2514 41644 4150
rect 41788 3392 41840 3398
rect 41788 3334 41840 3340
rect 41972 3392 42024 3398
rect 41972 3334 42024 3340
rect 42616 3392 42668 3398
rect 42616 3334 42668 3340
rect 41696 2848 41748 2854
rect 41696 2790 41748 2796
rect 41604 2508 41656 2514
rect 41604 2450 41656 2456
rect 41708 800 41736 2790
rect 41800 2514 41828 3334
rect 41984 3058 42012 3334
rect 41972 3052 42024 3058
rect 41972 2994 42024 3000
rect 41972 2916 42024 2922
rect 41972 2858 42024 2864
rect 41788 2508 41840 2514
rect 41788 2450 41840 2456
rect 41984 2378 42012 2858
rect 41972 2372 42024 2378
rect 41972 2314 42024 2320
rect 42628 800 42656 3334
rect 42720 2514 42748 4150
rect 42812 2990 42840 4422
rect 43352 4140 43404 4146
rect 43352 4082 43404 4088
rect 42892 3936 42944 3942
rect 42892 3878 42944 3884
rect 42800 2984 42852 2990
rect 42800 2926 42852 2932
rect 42904 2514 42932 3878
rect 43364 3602 43392 4082
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 42708 2508 42760 2514
rect 42708 2450 42760 2456
rect 42892 2508 42944 2514
rect 42892 2450 42944 2456
rect 43088 2378 43116 3538
rect 43548 3194 43576 4422
rect 43536 3188 43588 3194
rect 43536 3130 43588 3136
rect 43536 2440 43588 2446
rect 43536 2382 43588 2388
rect 43076 2372 43128 2378
rect 43076 2314 43128 2320
rect 43548 800 43576 2382
rect 44100 1358 44128 5102
rect 44180 4480 44232 4486
rect 44180 4422 44232 4428
rect 44192 2514 44220 4422
rect 44652 4282 44680 5510
rect 44640 4276 44692 4282
rect 44640 4218 44692 4224
rect 44640 4072 44692 4078
rect 44640 4014 44692 4020
rect 44364 3936 44416 3942
rect 44364 3878 44416 3884
rect 44376 2514 44404 3878
rect 44652 3602 44680 4014
rect 44640 3596 44692 3602
rect 44640 3538 44692 3544
rect 44732 2916 44784 2922
rect 44732 2858 44784 2864
rect 44456 2848 44508 2854
rect 44456 2790 44508 2796
rect 44180 2508 44232 2514
rect 44180 2450 44232 2456
rect 44364 2508 44416 2514
rect 44364 2450 44416 2456
rect 44088 1352 44140 1358
rect 44088 1294 44140 1300
rect 44468 800 44496 2790
rect 44744 2650 44772 2858
rect 44732 2644 44784 2650
rect 44732 2586 44784 2592
rect 44928 2106 44956 5510
rect 45008 5160 45060 5166
rect 45008 5102 45060 5108
rect 45020 4593 45048 5102
rect 45006 4584 45062 4593
rect 45006 4519 45062 4528
rect 45100 4480 45152 4486
rect 45100 4422 45152 4428
rect 45112 2514 45140 4422
rect 45100 2508 45152 2514
rect 45100 2450 45152 2456
rect 45204 2378 45232 6802
rect 45284 6248 45336 6254
rect 45284 6190 45336 6196
rect 46480 6248 46532 6254
rect 46480 6190 46532 6196
rect 45296 4826 45324 6190
rect 45376 6180 45428 6186
rect 45376 6122 45428 6128
rect 45284 4820 45336 4826
rect 45284 4762 45336 4768
rect 45388 3482 45416 6122
rect 45652 5160 45704 5166
rect 45652 5102 45704 5108
rect 45468 3936 45520 3942
rect 45468 3878 45520 3884
rect 45296 3454 45416 3482
rect 45296 2922 45324 3454
rect 45376 3392 45428 3398
rect 45376 3334 45428 3340
rect 45284 2916 45336 2922
rect 45284 2858 45336 2864
rect 45388 2774 45416 3334
rect 45480 3126 45508 3878
rect 45560 3732 45612 3738
rect 45560 3674 45612 3680
rect 45468 3120 45520 3126
rect 45468 3062 45520 3068
rect 45388 2746 45508 2774
rect 45192 2372 45244 2378
rect 45192 2314 45244 2320
rect 44916 2100 44968 2106
rect 44916 2042 44968 2048
rect 45480 800 45508 2746
rect 45572 2514 45600 3674
rect 45664 3058 45692 5102
rect 46388 4208 46440 4214
rect 46388 4150 46440 4156
rect 46400 4078 46428 4150
rect 46492 4078 46520 6190
rect 47124 5568 47176 5574
rect 47124 5510 47176 5516
rect 46940 5160 46992 5166
rect 46940 5102 46992 5108
rect 46572 4684 46624 4690
rect 46572 4626 46624 4632
rect 46584 4214 46612 4626
rect 46572 4208 46624 4214
rect 46572 4150 46624 4156
rect 45744 4072 45796 4078
rect 45744 4014 45796 4020
rect 46388 4072 46440 4078
rect 46388 4014 46440 4020
rect 46480 4072 46532 4078
rect 46480 4014 46532 4020
rect 45756 3602 45784 4014
rect 46400 3670 46428 4014
rect 46388 3664 46440 3670
rect 46388 3606 46440 3612
rect 45744 3596 45796 3602
rect 45744 3538 45796 3544
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 45652 3052 45704 3058
rect 45652 2994 45704 3000
rect 46308 2650 46336 3538
rect 46480 3392 46532 3398
rect 46480 3334 46532 3340
rect 46492 2774 46520 3334
rect 46756 2984 46808 2990
rect 46756 2926 46808 2932
rect 46400 2746 46520 2774
rect 46296 2644 46348 2650
rect 46296 2586 46348 2592
rect 45560 2508 45612 2514
rect 45560 2450 45612 2456
rect 46400 800 46428 2746
rect 46768 2582 46796 2926
rect 46756 2576 46808 2582
rect 46756 2518 46808 2524
rect 46952 2514 46980 5102
rect 47032 4004 47084 4010
rect 47032 3946 47084 3952
rect 47044 3738 47072 3946
rect 47032 3732 47084 3738
rect 47032 3674 47084 3680
rect 47032 3596 47084 3602
rect 47032 3538 47084 3544
rect 47044 3194 47072 3538
rect 47032 3188 47084 3194
rect 47032 3130 47084 3136
rect 47136 3058 47164 5510
rect 47228 4049 47256 7278
rect 47308 4684 47360 4690
rect 47308 4626 47360 4632
rect 47320 4078 47348 4626
rect 47400 4548 47452 4554
rect 47400 4490 47452 4496
rect 47308 4072 47360 4078
rect 47214 4040 47270 4049
rect 47308 4014 47360 4020
rect 47214 3975 47270 3984
rect 47216 3732 47268 3738
rect 47216 3674 47268 3680
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 47228 2514 47256 3674
rect 47308 3392 47360 3398
rect 47308 3334 47360 3340
rect 46940 2508 46992 2514
rect 46940 2450 46992 2456
rect 47216 2508 47268 2514
rect 47216 2450 47268 2456
rect 47320 800 47348 3334
rect 47412 3058 47440 4490
rect 47504 4214 47532 13330
rect 47584 13184 47636 13190
rect 47584 13126 47636 13132
rect 47596 8362 47624 13126
rect 49436 11694 49464 13738
rect 49424 11688 49476 11694
rect 49330 11656 49386 11665
rect 49424 11630 49476 11636
rect 49330 11591 49332 11600
rect 49384 11591 49386 11600
rect 49332 11562 49384 11568
rect 48872 9444 48924 9450
rect 48872 9386 48924 9392
rect 48044 9036 48096 9042
rect 48044 8978 48096 8984
rect 47768 8424 47820 8430
rect 47768 8366 47820 8372
rect 47584 8356 47636 8362
rect 47584 8298 47636 8304
rect 47780 7954 47808 8366
rect 47768 7948 47820 7954
rect 47768 7890 47820 7896
rect 47952 7948 48004 7954
rect 47952 7890 48004 7896
rect 47780 7750 47808 7890
rect 47768 7744 47820 7750
rect 47768 7686 47820 7692
rect 47584 7540 47636 7546
rect 47584 7482 47636 7488
rect 47492 4208 47544 4214
rect 47492 4150 47544 4156
rect 47596 3534 47624 7482
rect 47780 6186 47808 7686
rect 47964 7546 47992 7890
rect 47952 7540 48004 7546
rect 47952 7482 48004 7488
rect 47860 7336 47912 7342
rect 47860 7278 47912 7284
rect 47872 6934 47900 7278
rect 47860 6928 47912 6934
rect 47860 6870 47912 6876
rect 47768 6180 47820 6186
rect 47768 6122 47820 6128
rect 47780 5778 47808 6122
rect 47768 5772 47820 5778
rect 47768 5714 47820 5720
rect 47780 5166 47808 5714
rect 48056 5642 48084 8978
rect 48688 8832 48740 8838
rect 48688 8774 48740 8780
rect 48412 7948 48464 7954
rect 48412 7890 48464 7896
rect 48424 7721 48452 7890
rect 48700 7857 48728 8774
rect 48884 8498 48912 9386
rect 49516 9036 49568 9042
rect 49516 8978 49568 8984
rect 48872 8492 48924 8498
rect 48872 8434 48924 8440
rect 48686 7848 48742 7857
rect 48686 7783 48742 7792
rect 48410 7712 48466 7721
rect 48410 7647 48466 7656
rect 48320 6248 48372 6254
rect 48320 6190 48372 6196
rect 48044 5636 48096 5642
rect 48044 5578 48096 5584
rect 48136 5568 48188 5574
rect 48136 5510 48188 5516
rect 47768 5160 47820 5166
rect 47768 5102 47820 5108
rect 47860 5160 47912 5166
rect 47860 5102 47912 5108
rect 47768 4820 47820 4826
rect 47768 4762 47820 4768
rect 47780 4554 47808 4762
rect 47872 4758 47900 5102
rect 48148 4978 48176 5510
rect 48332 5166 48360 6190
rect 48424 5778 48452 7647
rect 48778 6896 48834 6905
rect 48778 6831 48780 6840
rect 48832 6831 48834 6840
rect 48780 6802 48832 6808
rect 48688 6792 48740 6798
rect 48686 6760 48688 6769
rect 48740 6760 48742 6769
rect 48686 6695 48742 6704
rect 48596 6656 48648 6662
rect 48596 6598 48648 6604
rect 48412 5772 48464 5778
rect 48412 5714 48464 5720
rect 48320 5160 48372 5166
rect 48320 5102 48372 5108
rect 48056 4950 48176 4978
rect 47952 4820 48004 4826
rect 47952 4762 48004 4768
rect 47860 4752 47912 4758
rect 47860 4694 47912 4700
rect 47964 4690 47992 4762
rect 47952 4684 48004 4690
rect 47952 4626 48004 4632
rect 47768 4548 47820 4554
rect 47768 4490 47820 4496
rect 47676 4480 47728 4486
rect 47676 4422 47728 4428
rect 47952 4480 48004 4486
rect 47952 4422 48004 4428
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47400 3052 47452 3058
rect 47400 2994 47452 3000
rect 47688 2038 47716 4422
rect 47768 3596 47820 3602
rect 47768 3538 47820 3544
rect 47860 3596 47912 3602
rect 47860 3538 47912 3544
rect 47780 2650 47808 3538
rect 47872 3194 47900 3538
rect 47964 3534 47992 4422
rect 48056 3738 48084 4950
rect 48134 4584 48190 4593
rect 48134 4519 48136 4528
rect 48188 4519 48190 4528
rect 48136 4490 48188 4496
rect 48136 3936 48188 3942
rect 48136 3878 48188 3884
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 47952 3528 48004 3534
rect 47952 3470 48004 3476
rect 47860 3188 47912 3194
rect 47860 3130 47912 3136
rect 47768 2644 47820 2650
rect 47768 2586 47820 2592
rect 47676 2032 47728 2038
rect 47676 1974 47728 1980
rect 48148 1970 48176 3878
rect 48228 3392 48280 3398
rect 48228 3334 48280 3340
rect 48136 1964 48188 1970
rect 48136 1906 48188 1912
rect 48240 800 48268 3334
rect 48424 2854 48452 5714
rect 48608 3058 48636 6598
rect 48884 6202 48912 8434
rect 49332 8084 49384 8090
rect 49332 8026 49384 8032
rect 49344 7993 49372 8026
rect 49330 7984 49386 7993
rect 48964 7948 49016 7954
rect 49528 7954 49556 8978
rect 49608 8968 49660 8974
rect 49608 8910 49660 8916
rect 49330 7919 49386 7928
rect 49516 7948 49568 7954
rect 48964 7890 49016 7896
rect 49516 7890 49568 7896
rect 48976 7342 49004 7890
rect 49620 7478 49648 8910
rect 49712 7546 49740 14010
rect 49804 11694 49832 14962
rect 49988 14482 50016 15846
rect 49976 14476 50028 14482
rect 49896 14436 49976 14464
rect 49896 13394 49924 14436
rect 49976 14418 50028 14424
rect 50172 13784 50200 16646
rect 50300 15804 50596 15824
rect 50356 15802 50380 15804
rect 50436 15802 50460 15804
rect 50516 15802 50540 15804
rect 50378 15750 50380 15802
rect 50442 15750 50454 15802
rect 50516 15750 50518 15802
rect 50356 15748 50380 15750
rect 50436 15748 50460 15750
rect 50516 15748 50540 15750
rect 50300 15728 50596 15748
rect 50300 14716 50596 14736
rect 50356 14714 50380 14716
rect 50436 14714 50460 14716
rect 50516 14714 50540 14716
rect 50378 14662 50380 14714
rect 50442 14662 50454 14714
rect 50516 14662 50518 14714
rect 50356 14660 50380 14662
rect 50436 14660 50460 14662
rect 50516 14660 50540 14662
rect 50300 14640 50596 14660
rect 50434 14512 50490 14521
rect 50434 14447 50490 14456
rect 50252 14408 50304 14414
rect 50252 14350 50304 14356
rect 50264 13802 50292 14350
rect 50448 13870 50476 14447
rect 50436 13864 50488 13870
rect 50436 13806 50488 13812
rect 50080 13756 50200 13784
rect 50252 13796 50304 13802
rect 49884 13388 49936 13394
rect 49884 13330 49936 13336
rect 49896 12306 49924 13330
rect 49884 12300 49936 12306
rect 49884 12242 49936 12248
rect 49884 12096 49936 12102
rect 49884 12038 49936 12044
rect 49792 11688 49844 11694
rect 49792 11630 49844 11636
rect 49700 7540 49752 7546
rect 49700 7482 49752 7488
rect 49608 7472 49660 7478
rect 49608 7414 49660 7420
rect 48964 7336 49016 7342
rect 48964 7278 49016 7284
rect 48792 6174 48912 6202
rect 48688 6112 48740 6118
rect 48688 6054 48740 6060
rect 48596 3052 48648 3058
rect 48596 2994 48648 3000
rect 48412 2848 48464 2854
rect 48412 2790 48464 2796
rect 48700 2774 48728 6054
rect 48792 5166 48820 6174
rect 48976 6118 49004 7278
rect 49698 6896 49754 6905
rect 49698 6831 49754 6840
rect 49712 6798 49740 6831
rect 49700 6792 49752 6798
rect 49804 6769 49832 11630
rect 49896 8922 49924 12038
rect 50080 10198 50108 13756
rect 50252 13738 50304 13744
rect 50300 13628 50596 13648
rect 50356 13626 50380 13628
rect 50436 13626 50460 13628
rect 50516 13626 50540 13628
rect 50378 13574 50380 13626
rect 50442 13574 50454 13626
rect 50516 13574 50518 13626
rect 50356 13572 50380 13574
rect 50436 13572 50460 13574
rect 50516 13572 50540 13574
rect 50300 13552 50596 13572
rect 50436 13320 50488 13326
rect 50436 13262 50488 13268
rect 50448 12782 50476 13262
rect 50436 12776 50488 12782
rect 50436 12718 50488 12724
rect 50300 12540 50596 12560
rect 50356 12538 50380 12540
rect 50436 12538 50460 12540
rect 50516 12538 50540 12540
rect 50378 12486 50380 12538
rect 50442 12486 50454 12538
rect 50516 12486 50518 12538
rect 50356 12484 50380 12486
rect 50436 12484 50460 12486
rect 50516 12484 50540 12486
rect 50300 12464 50596 12484
rect 50632 12434 50660 18702
rect 50710 18592 50766 18601
rect 50710 18527 50766 18536
rect 50724 18222 50752 18527
rect 50712 18216 50764 18222
rect 50712 18158 50764 18164
rect 50724 18086 50752 18158
rect 50712 18080 50764 18086
rect 50712 18022 50764 18028
rect 50712 16992 50764 16998
rect 50712 16934 50764 16940
rect 50724 16726 50752 16934
rect 50712 16720 50764 16726
rect 50712 16662 50764 16668
rect 50816 16046 50844 23666
rect 50908 20040 50936 26846
rect 51000 26586 51028 26862
rect 50988 26580 51040 26586
rect 50988 26522 51040 26528
rect 51092 25770 51120 27950
rect 51276 27674 51304 29718
rect 51264 27668 51316 27674
rect 51264 27610 51316 27616
rect 51172 27464 51224 27470
rect 51172 27406 51224 27412
rect 51184 26994 51212 27406
rect 51172 26988 51224 26994
rect 51172 26930 51224 26936
rect 51080 25764 51132 25770
rect 51080 25706 51132 25712
rect 51092 24682 51120 25706
rect 50988 24676 51040 24682
rect 50988 24618 51040 24624
rect 51080 24676 51132 24682
rect 51080 24618 51132 24624
rect 51000 20262 51028 24618
rect 51368 22166 51396 33254
rect 51460 31482 51488 34954
rect 51736 34746 51764 35566
rect 51816 35488 51868 35494
rect 51816 35430 51868 35436
rect 51828 35222 51856 35430
rect 51816 35216 51868 35222
rect 51816 35158 51868 35164
rect 52104 34746 52132 35566
rect 53012 35556 53064 35562
rect 53012 35498 53064 35504
rect 53024 34950 53052 35498
rect 53116 35494 53144 35566
rect 53104 35488 53156 35494
rect 53104 35430 53156 35436
rect 53012 34944 53064 34950
rect 53012 34886 53064 34892
rect 51724 34740 51776 34746
rect 51724 34682 51776 34688
rect 52092 34740 52144 34746
rect 52092 34682 52144 34688
rect 51908 34536 51960 34542
rect 53116 34524 53144 35430
rect 53196 35012 53248 35018
rect 53196 34954 53248 34960
rect 51908 34478 51960 34484
rect 52840 34496 53144 34524
rect 51920 34202 51948 34478
rect 52368 34468 52420 34474
rect 52368 34410 52420 34416
rect 51908 34196 51960 34202
rect 51908 34138 51960 34144
rect 52184 34060 52236 34066
rect 52184 34002 52236 34008
rect 51540 32972 51592 32978
rect 51540 32914 51592 32920
rect 51552 32570 51580 32914
rect 51540 32564 51592 32570
rect 51540 32506 51592 32512
rect 52196 32502 52224 34002
rect 52380 33538 52408 34410
rect 52736 34400 52788 34406
rect 52736 34342 52788 34348
rect 52748 34202 52776 34342
rect 52736 34196 52788 34202
rect 52736 34138 52788 34144
rect 52840 34082 52868 34496
rect 52920 34400 52972 34406
rect 52920 34342 52972 34348
rect 52748 34054 52868 34082
rect 52460 33992 52512 33998
rect 52460 33934 52512 33940
rect 52472 33658 52500 33934
rect 52460 33652 52512 33658
rect 52460 33594 52512 33600
rect 52288 33510 52408 33538
rect 52550 33552 52606 33561
rect 52288 33318 52316 33510
rect 52550 33487 52606 33496
rect 52564 33454 52592 33487
rect 52552 33448 52604 33454
rect 52552 33390 52604 33396
rect 52276 33312 52328 33318
rect 52748 33266 52776 34054
rect 52932 33590 52960 34342
rect 53012 33924 53064 33930
rect 53012 33866 53064 33872
rect 52920 33584 52972 33590
rect 52920 33526 52972 33532
rect 52828 33448 52880 33454
rect 52828 33390 52880 33396
rect 52276 33254 52328 33260
rect 52656 33238 52776 33266
rect 52656 33114 52684 33238
rect 52840 33114 52868 33390
rect 52644 33108 52696 33114
rect 52644 33050 52696 33056
rect 52828 33108 52880 33114
rect 52828 33050 52880 33056
rect 52368 33040 52420 33046
rect 52368 32982 52420 32988
rect 52184 32496 52236 32502
rect 52184 32438 52236 32444
rect 52196 32366 52224 32438
rect 52000 32360 52052 32366
rect 52000 32302 52052 32308
rect 52184 32360 52236 32366
rect 52184 32302 52236 32308
rect 51724 32292 51776 32298
rect 51724 32234 51776 32240
rect 51736 32026 51764 32234
rect 51724 32020 51776 32026
rect 51724 31962 51776 31968
rect 51814 31920 51870 31929
rect 51814 31855 51816 31864
rect 51868 31855 51870 31864
rect 51816 31826 51868 31832
rect 51908 31816 51960 31822
rect 51908 31758 51960 31764
rect 51448 31476 51500 31482
rect 51448 31418 51500 31424
rect 51540 31408 51592 31414
rect 51540 31350 51592 31356
rect 51552 31142 51580 31350
rect 51920 31260 51948 31758
rect 52012 31414 52040 32302
rect 52276 32292 52328 32298
rect 52276 32234 52328 32240
rect 52184 31680 52236 31686
rect 52184 31622 52236 31628
rect 52000 31408 52052 31414
rect 52000 31350 52052 31356
rect 52000 31272 52052 31278
rect 51920 31232 52000 31260
rect 52000 31214 52052 31220
rect 51724 31204 51776 31210
rect 51724 31146 51776 31152
rect 51540 31136 51592 31142
rect 51540 31078 51592 31084
rect 51448 30660 51500 30666
rect 51448 30602 51500 30608
rect 51460 29238 51488 30602
rect 51552 30394 51580 31078
rect 51736 30802 51764 31146
rect 52012 30870 52040 31214
rect 52092 31136 52144 31142
rect 52092 31078 52144 31084
rect 52000 30864 52052 30870
rect 52000 30806 52052 30812
rect 51724 30796 51776 30802
rect 51724 30738 51776 30744
rect 51540 30388 51592 30394
rect 51540 30330 51592 30336
rect 52012 29782 52040 30806
rect 52000 29776 52052 29782
rect 52000 29718 52052 29724
rect 51540 29504 51592 29510
rect 51540 29446 51592 29452
rect 51552 29306 51580 29446
rect 51540 29300 51592 29306
rect 51540 29242 51592 29248
rect 51448 29232 51500 29238
rect 51448 29174 51500 29180
rect 51448 29096 51500 29102
rect 51724 29096 51776 29102
rect 51500 29056 51672 29084
rect 51448 29038 51500 29044
rect 51460 28762 51488 29038
rect 51448 28756 51500 28762
rect 51448 28698 51500 28704
rect 51644 28694 51672 29056
rect 52000 29096 52052 29102
rect 51776 29056 51856 29084
rect 51724 29038 51776 29044
rect 51724 28960 51776 28966
rect 51724 28902 51776 28908
rect 51632 28688 51684 28694
rect 51632 28630 51684 28636
rect 51736 28626 51764 28902
rect 51724 28620 51776 28626
rect 51724 28562 51776 28568
rect 51540 28008 51592 28014
rect 51540 27950 51592 27956
rect 51356 22160 51408 22166
rect 51356 22102 51408 22108
rect 51264 20936 51316 20942
rect 51264 20878 51316 20884
rect 51276 20602 51304 20878
rect 51264 20596 51316 20602
rect 51264 20538 51316 20544
rect 50988 20256 51040 20262
rect 50988 20198 51040 20204
rect 50908 20012 51028 20040
rect 50896 19916 50948 19922
rect 50896 19858 50948 19864
rect 50908 19786 50936 19858
rect 50896 19780 50948 19786
rect 50896 19722 50948 19728
rect 50896 19168 50948 19174
rect 50896 19110 50948 19116
rect 50804 16040 50856 16046
rect 50804 15982 50856 15988
rect 50712 15564 50764 15570
rect 50712 15506 50764 15512
rect 50724 13870 50752 15506
rect 50712 13864 50764 13870
rect 50712 13806 50764 13812
rect 50724 13705 50752 13806
rect 50710 13696 50766 13705
rect 50710 13631 50766 13640
rect 50632 12406 50752 12434
rect 50526 12336 50582 12345
rect 50526 12271 50528 12280
rect 50580 12271 50582 12280
rect 50528 12242 50580 12248
rect 50620 11688 50672 11694
rect 50620 11630 50672 11636
rect 50724 11642 50752 12406
rect 50816 12102 50844 15982
rect 50908 13954 50936 19110
rect 51000 14249 51028 20012
rect 51078 19000 51134 19009
rect 51078 18935 51134 18944
rect 51092 18698 51120 18935
rect 51080 18692 51132 18698
rect 51080 18634 51132 18640
rect 51264 18692 51316 18698
rect 51264 18634 51316 18640
rect 51276 18601 51304 18634
rect 51262 18592 51318 18601
rect 51262 18527 51318 18536
rect 51172 18216 51224 18222
rect 51172 18158 51224 18164
rect 51184 17746 51212 18158
rect 51368 17762 51396 22102
rect 51552 22094 51580 27950
rect 51828 27538 51856 29056
rect 52000 29038 52052 29044
rect 51908 29028 51960 29034
rect 51908 28970 51960 28976
rect 51920 28626 51948 28970
rect 51908 28620 51960 28626
rect 51908 28562 51960 28568
rect 51724 27532 51776 27538
rect 51724 27474 51776 27480
rect 51816 27532 51868 27538
rect 51816 27474 51868 27480
rect 51632 27328 51684 27334
rect 51632 27270 51684 27276
rect 51644 27130 51672 27270
rect 51632 27124 51684 27130
rect 51632 27066 51684 27072
rect 51736 26926 51764 27474
rect 51724 26920 51776 26926
rect 51724 26862 51776 26868
rect 51724 26444 51776 26450
rect 51828 26432 51856 27474
rect 52012 27334 52040 29038
rect 52104 27826 52132 31078
rect 52196 30938 52224 31622
rect 52184 30932 52236 30938
rect 52184 30874 52236 30880
rect 52288 30326 52316 32234
rect 52380 31890 52408 32982
rect 52552 32836 52604 32842
rect 52552 32778 52604 32784
rect 52368 31884 52420 31890
rect 52368 31826 52420 31832
rect 52460 31884 52512 31890
rect 52460 31826 52512 31832
rect 52380 31278 52408 31826
rect 52472 31686 52500 31826
rect 52564 31754 52592 32778
rect 52736 32768 52788 32774
rect 52736 32710 52788 32716
rect 52748 32570 52776 32710
rect 52736 32564 52788 32570
rect 52736 32506 52788 32512
rect 53024 32434 53052 33866
rect 53208 33318 53236 34954
rect 53564 34536 53616 34542
rect 53564 34478 53616 34484
rect 53380 34060 53432 34066
rect 53380 34002 53432 34008
rect 53288 33856 53340 33862
rect 53286 33824 53288 33833
rect 53340 33824 53342 33833
rect 53286 33759 53342 33768
rect 53300 33454 53328 33759
rect 53392 33522 53420 34002
rect 53380 33516 53432 33522
rect 53380 33458 53432 33464
rect 53288 33448 53340 33454
rect 53288 33390 53340 33396
rect 53472 33448 53524 33454
rect 53472 33390 53524 33396
rect 53196 33312 53248 33318
rect 53196 33254 53248 33260
rect 53012 32428 53064 32434
rect 53012 32370 53064 32376
rect 53288 32360 53340 32366
rect 53288 32302 53340 32308
rect 52736 31816 52788 31822
rect 52736 31758 52788 31764
rect 52552 31748 52604 31754
rect 52552 31690 52604 31696
rect 52460 31680 52512 31686
rect 52460 31622 52512 31628
rect 52748 31482 52776 31758
rect 52736 31476 52788 31482
rect 52736 31418 52788 31424
rect 52368 31272 52420 31278
rect 52368 31214 52420 31220
rect 52380 30938 52408 31214
rect 52828 31136 52880 31142
rect 52828 31078 52880 31084
rect 52920 31136 52972 31142
rect 52920 31078 52972 31084
rect 52368 30932 52420 30938
rect 52368 30874 52420 30880
rect 52380 30802 52408 30874
rect 52840 30802 52868 31078
rect 52368 30796 52420 30802
rect 52368 30738 52420 30744
rect 52644 30796 52696 30802
rect 52644 30738 52696 30744
rect 52828 30796 52880 30802
rect 52828 30738 52880 30744
rect 52380 30326 52408 30738
rect 52656 30546 52684 30738
rect 52932 30666 52960 31078
rect 52920 30660 52972 30666
rect 52920 30602 52972 30608
rect 52656 30518 53052 30546
rect 52656 30394 52684 30518
rect 52644 30388 52696 30394
rect 52644 30330 52696 30336
rect 52276 30320 52328 30326
rect 52276 30262 52328 30268
rect 52368 30320 52420 30326
rect 52368 30262 52420 30268
rect 52368 30184 52420 30190
rect 52368 30126 52420 30132
rect 52460 30184 52512 30190
rect 52460 30126 52512 30132
rect 52380 29714 52408 30126
rect 52472 29714 52500 30126
rect 52828 29776 52880 29782
rect 52828 29718 52880 29724
rect 52368 29708 52420 29714
rect 52368 29650 52420 29656
rect 52460 29708 52512 29714
rect 52460 29650 52512 29656
rect 52276 29640 52328 29646
rect 52276 29582 52328 29588
rect 52182 28656 52238 28665
rect 52182 28591 52184 28600
rect 52236 28591 52238 28600
rect 52184 28562 52236 28568
rect 52184 28484 52236 28490
rect 52184 28426 52236 28432
rect 52196 27946 52224 28426
rect 52288 28014 52316 29582
rect 52380 29170 52408 29650
rect 52368 29164 52420 29170
rect 52368 29106 52420 29112
rect 52472 28762 52500 29650
rect 52840 29186 52868 29718
rect 52748 29158 52868 29186
rect 52644 29096 52696 29102
rect 52644 29038 52696 29044
rect 52460 28756 52512 28762
rect 52460 28698 52512 28704
rect 52460 28620 52512 28626
rect 52460 28562 52512 28568
rect 52472 28218 52500 28562
rect 52460 28212 52512 28218
rect 52460 28154 52512 28160
rect 52276 28008 52328 28014
rect 52276 27950 52328 27956
rect 52184 27940 52236 27946
rect 52184 27882 52236 27888
rect 52104 27798 52224 27826
rect 52000 27328 52052 27334
rect 52000 27270 52052 27276
rect 51908 26444 51960 26450
rect 51828 26404 51908 26432
rect 51724 26386 51776 26392
rect 51908 26386 51960 26392
rect 51736 26042 51764 26386
rect 52012 26246 52040 27270
rect 51816 26240 51868 26246
rect 51816 26182 51868 26188
rect 52000 26240 52052 26246
rect 52000 26182 52052 26188
rect 51724 26036 51776 26042
rect 51724 25978 51776 25984
rect 51632 25764 51684 25770
rect 51632 25706 51684 25712
rect 51644 25362 51672 25706
rect 51828 25498 51856 26182
rect 52012 26058 52040 26182
rect 52012 26042 52132 26058
rect 52012 26036 52144 26042
rect 52012 26030 52092 26036
rect 52092 25978 52144 25984
rect 51906 25936 51962 25945
rect 51906 25871 51962 25880
rect 52092 25900 52144 25906
rect 51816 25492 51868 25498
rect 51816 25434 51868 25440
rect 51632 25356 51684 25362
rect 51632 25298 51684 25304
rect 51920 24410 51948 25871
rect 52092 25842 52144 25848
rect 52000 25356 52052 25362
rect 52000 25298 52052 25304
rect 52012 24970 52040 25298
rect 52104 25158 52132 25842
rect 52092 25152 52144 25158
rect 52092 25094 52144 25100
rect 52012 24942 52132 24970
rect 51908 24404 51960 24410
rect 51908 24346 51960 24352
rect 52104 24274 52132 24942
rect 52092 24268 52144 24274
rect 52092 24210 52144 24216
rect 52104 23730 52132 24210
rect 52092 23724 52144 23730
rect 52092 23666 52144 23672
rect 52092 23180 52144 23186
rect 52092 23122 52144 23128
rect 52000 22976 52052 22982
rect 52000 22918 52052 22924
rect 51722 22808 51778 22817
rect 51722 22743 51724 22752
rect 51776 22743 51778 22752
rect 51724 22714 51776 22720
rect 52012 22438 52040 22918
rect 52104 22778 52132 23122
rect 52092 22772 52144 22778
rect 52092 22714 52144 22720
rect 52000 22432 52052 22438
rect 52000 22374 52052 22380
rect 51552 22066 51856 22094
rect 51828 21690 51856 22066
rect 51816 21684 51868 21690
rect 51816 21626 51868 21632
rect 51724 21616 51776 21622
rect 51724 21558 51776 21564
rect 51632 21344 51684 21350
rect 51632 21286 51684 21292
rect 51644 20913 51672 21286
rect 51630 20904 51686 20913
rect 51736 20874 51764 21558
rect 51630 20839 51686 20848
rect 51724 20868 51776 20874
rect 51724 20810 51776 20816
rect 52000 20800 52052 20806
rect 52000 20742 52052 20748
rect 52012 20505 52040 20742
rect 51998 20496 52054 20505
rect 51998 20431 52054 20440
rect 51448 20392 51500 20398
rect 51448 20334 51500 20340
rect 51460 20262 51488 20334
rect 51448 20256 51500 20262
rect 51448 20198 51500 20204
rect 51460 20058 51488 20198
rect 51448 20052 51500 20058
rect 51448 19994 51500 20000
rect 51448 19780 51500 19786
rect 51448 19722 51500 19728
rect 51460 18834 51488 19722
rect 51540 19712 51592 19718
rect 51540 19654 51592 19660
rect 51552 19417 51580 19654
rect 51538 19408 51594 19417
rect 51538 19343 51594 19352
rect 51448 18828 51500 18834
rect 51448 18770 51500 18776
rect 51448 18624 51500 18630
rect 51448 18566 51500 18572
rect 51460 18358 51488 18566
rect 51448 18352 51500 18358
rect 51448 18294 51500 18300
rect 51460 18086 51488 18294
rect 51552 18222 51580 19343
rect 52092 19304 52144 19310
rect 52092 19246 52144 19252
rect 51908 19236 51960 19242
rect 51908 19178 51960 19184
rect 51632 19168 51684 19174
rect 51632 19110 51684 19116
rect 51644 18834 51672 19110
rect 51814 18864 51870 18873
rect 51632 18828 51684 18834
rect 51814 18799 51870 18808
rect 51632 18770 51684 18776
rect 51644 18578 51672 18770
rect 51828 18630 51856 18799
rect 51816 18624 51868 18630
rect 51644 18550 51764 18578
rect 51816 18566 51868 18572
rect 51540 18216 51592 18222
rect 51540 18158 51592 18164
rect 51448 18080 51500 18086
rect 51448 18022 51500 18028
rect 51172 17740 51224 17746
rect 51172 17682 51224 17688
rect 51276 17734 51396 17762
rect 51184 17270 51212 17682
rect 51172 17264 51224 17270
rect 51172 17206 51224 17212
rect 51172 16584 51224 16590
rect 51172 16526 51224 16532
rect 51184 15706 51212 16526
rect 51276 16046 51304 17734
rect 51460 17678 51488 18022
rect 51736 17746 51764 18550
rect 51920 18358 51948 19178
rect 51908 18352 51960 18358
rect 51908 18294 51960 18300
rect 52000 18284 52052 18290
rect 52000 18226 52052 18232
rect 52012 17746 52040 18226
rect 51724 17740 51776 17746
rect 51724 17682 51776 17688
rect 52000 17740 52052 17746
rect 52000 17682 52052 17688
rect 51356 17672 51408 17678
rect 51354 17640 51356 17649
rect 51448 17672 51500 17678
rect 51408 17640 51410 17649
rect 51448 17614 51500 17620
rect 51354 17575 51410 17584
rect 51356 17536 51408 17542
rect 51356 17478 51408 17484
rect 51632 17536 51684 17542
rect 52104 17513 52132 19246
rect 51632 17478 51684 17484
rect 52090 17504 52146 17513
rect 51368 17270 51396 17478
rect 51446 17368 51502 17377
rect 51446 17303 51502 17312
rect 51356 17264 51408 17270
rect 51356 17206 51408 17212
rect 51460 16658 51488 17303
rect 51644 17202 51672 17478
rect 52090 17439 52146 17448
rect 51632 17196 51684 17202
rect 51632 17138 51684 17144
rect 51644 16658 51672 17138
rect 51356 16652 51408 16658
rect 51356 16594 51408 16600
rect 51448 16652 51500 16658
rect 51448 16594 51500 16600
rect 51632 16652 51684 16658
rect 51632 16594 51684 16600
rect 51264 16040 51316 16046
rect 51264 15982 51316 15988
rect 51368 15978 51396 16594
rect 51632 16040 51684 16046
rect 51632 15982 51684 15988
rect 52000 16040 52052 16046
rect 52000 15982 52052 15988
rect 51356 15972 51408 15978
rect 51356 15914 51408 15920
rect 51172 15700 51224 15706
rect 51172 15642 51224 15648
rect 51264 15360 51316 15366
rect 51264 15302 51316 15308
rect 51276 14482 51304 15302
rect 51264 14476 51316 14482
rect 51264 14418 51316 14424
rect 51368 14414 51396 15914
rect 51448 14884 51500 14890
rect 51448 14826 51500 14832
rect 51356 14408 51408 14414
rect 51356 14350 51408 14356
rect 50986 14240 51042 14249
rect 50986 14175 51042 14184
rect 51000 14074 51028 14175
rect 50988 14068 51040 14074
rect 50988 14010 51040 14016
rect 50986 13968 51042 13977
rect 50908 13926 50986 13954
rect 50986 13903 51042 13912
rect 51000 12986 51028 13903
rect 51264 13864 51316 13870
rect 51264 13806 51316 13812
rect 51080 13728 51132 13734
rect 51080 13670 51132 13676
rect 51092 13462 51120 13670
rect 51080 13456 51132 13462
rect 51080 13398 51132 13404
rect 50988 12980 51040 12986
rect 50988 12922 51040 12928
rect 50896 12232 50948 12238
rect 50896 12174 50948 12180
rect 50908 12102 50936 12174
rect 50804 12096 50856 12102
rect 50804 12038 50856 12044
rect 50896 12096 50948 12102
rect 50896 12038 50948 12044
rect 50300 11452 50596 11472
rect 50356 11450 50380 11452
rect 50436 11450 50460 11452
rect 50516 11450 50540 11452
rect 50378 11398 50380 11450
rect 50442 11398 50454 11450
rect 50516 11398 50518 11450
rect 50356 11396 50380 11398
rect 50436 11396 50460 11398
rect 50516 11396 50540 11398
rect 50300 11376 50596 11396
rect 50632 11218 50660 11630
rect 50724 11614 50936 11642
rect 50712 11348 50764 11354
rect 50712 11290 50764 11296
rect 50620 11212 50672 11218
rect 50620 11154 50672 11160
rect 50300 10364 50596 10384
rect 50356 10362 50380 10364
rect 50436 10362 50460 10364
rect 50516 10362 50540 10364
rect 50378 10310 50380 10362
rect 50442 10310 50454 10362
rect 50516 10310 50518 10362
rect 50356 10308 50380 10310
rect 50436 10308 50460 10310
rect 50516 10308 50540 10310
rect 50300 10288 50596 10308
rect 50068 10192 50120 10198
rect 50068 10134 50120 10140
rect 49976 10124 50028 10130
rect 49976 10066 50028 10072
rect 49988 9178 50016 10066
rect 50160 10056 50212 10062
rect 50160 9998 50212 10004
rect 50172 9586 50200 9998
rect 50344 9920 50396 9926
rect 50344 9862 50396 9868
rect 50160 9580 50212 9586
rect 50160 9522 50212 9528
rect 50356 9518 50384 9862
rect 50724 9654 50752 11290
rect 50804 10600 50856 10606
rect 50804 10542 50856 10548
rect 50816 10266 50844 10542
rect 50804 10260 50856 10266
rect 50804 10202 50856 10208
rect 50712 9648 50764 9654
rect 50712 9590 50764 9596
rect 50344 9512 50396 9518
rect 50344 9454 50396 9460
rect 50160 9376 50212 9382
rect 50160 9318 50212 9324
rect 49976 9172 50028 9178
rect 49976 9114 50028 9120
rect 50172 9042 50200 9318
rect 50300 9276 50596 9296
rect 50356 9274 50380 9276
rect 50436 9274 50460 9276
rect 50516 9274 50540 9276
rect 50378 9222 50380 9274
rect 50442 9222 50454 9274
rect 50516 9222 50518 9274
rect 50356 9220 50380 9222
rect 50436 9220 50460 9222
rect 50516 9220 50540 9222
rect 50300 9200 50596 9220
rect 50712 9172 50764 9178
rect 50712 9114 50764 9120
rect 50160 9036 50212 9042
rect 50160 8978 50212 8984
rect 50252 9036 50304 9042
rect 50252 8978 50304 8984
rect 49896 8894 50016 8922
rect 49884 8832 49936 8838
rect 49884 8774 49936 8780
rect 49896 7954 49924 8774
rect 49884 7948 49936 7954
rect 49884 7890 49936 7896
rect 49700 6734 49752 6740
rect 49790 6760 49846 6769
rect 49790 6695 49846 6704
rect 49700 6656 49752 6662
rect 49700 6598 49752 6604
rect 49516 6248 49568 6254
rect 49712 6236 49740 6598
rect 49568 6208 49832 6236
rect 49516 6190 49568 6196
rect 49424 6180 49476 6186
rect 49424 6122 49476 6128
rect 48872 6112 48924 6118
rect 48872 6054 48924 6060
rect 48964 6112 49016 6118
rect 48964 6054 49016 6060
rect 48780 5160 48832 5166
rect 48780 5102 48832 5108
rect 48780 4684 48832 4690
rect 48780 4626 48832 4632
rect 48792 3670 48820 4626
rect 48780 3664 48832 3670
rect 48780 3606 48832 3612
rect 48700 2746 48820 2774
rect 48792 2514 48820 2746
rect 48884 2582 48912 6054
rect 49056 5772 49108 5778
rect 49056 5714 49108 5720
rect 49068 4826 49096 5714
rect 49332 5568 49384 5574
rect 49332 5510 49384 5516
rect 49148 5228 49200 5234
rect 49148 5170 49200 5176
rect 49056 4820 49108 4826
rect 49056 4762 49108 4768
rect 48964 3460 49016 3466
rect 48964 3402 49016 3408
rect 49056 3460 49108 3466
rect 49056 3402 49108 3408
rect 48976 3058 49004 3402
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 49068 2922 49096 3402
rect 49160 3369 49188 5170
rect 49240 5160 49292 5166
rect 49238 5128 49240 5137
rect 49292 5128 49294 5137
rect 49238 5063 49294 5072
rect 49240 4480 49292 4486
rect 49240 4422 49292 4428
rect 49146 3360 49202 3369
rect 49146 3295 49202 3304
rect 49252 3194 49280 4422
rect 49240 3188 49292 3194
rect 49240 3130 49292 3136
rect 49344 2990 49372 5510
rect 49436 5273 49464 6122
rect 49608 6112 49660 6118
rect 49608 6054 49660 6060
rect 49620 5817 49648 6054
rect 49606 5808 49662 5817
rect 49606 5743 49608 5752
rect 49660 5743 49662 5752
rect 49608 5714 49660 5720
rect 49700 5364 49752 5370
rect 49700 5306 49752 5312
rect 49422 5264 49478 5273
rect 49422 5199 49478 5208
rect 49436 5030 49464 5199
rect 49424 5024 49476 5030
rect 49424 4966 49476 4972
rect 49608 4684 49660 4690
rect 49608 4626 49660 4632
rect 49516 4140 49568 4146
rect 49516 4082 49568 4088
rect 49424 3936 49476 3942
rect 49424 3878 49476 3884
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 49056 2916 49108 2922
rect 49056 2858 49108 2864
rect 49148 2848 49200 2854
rect 49148 2790 49200 2796
rect 48872 2576 48924 2582
rect 48872 2518 48924 2524
rect 48780 2508 48832 2514
rect 48780 2450 48832 2456
rect 49160 800 49188 2790
rect 49436 1902 49464 3878
rect 49528 2378 49556 4082
rect 49620 4078 49648 4626
rect 49608 4072 49660 4078
rect 49608 4014 49660 4020
rect 49620 3602 49648 4014
rect 49608 3596 49660 3602
rect 49608 3538 49660 3544
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 49620 3097 49648 3334
rect 49606 3088 49662 3097
rect 49606 3023 49662 3032
rect 49712 2514 49740 5306
rect 49804 4486 49832 6208
rect 49896 4690 49924 7890
rect 49988 6662 50016 8894
rect 50172 8498 50200 8978
rect 50264 8566 50292 8978
rect 50252 8560 50304 8566
rect 50252 8502 50304 8508
rect 50160 8492 50212 8498
rect 50160 8434 50212 8440
rect 50068 8356 50120 8362
rect 50068 8298 50120 8304
rect 50080 8090 50108 8298
rect 50620 8288 50672 8294
rect 50620 8230 50672 8236
rect 50300 8188 50596 8208
rect 50356 8186 50380 8188
rect 50436 8186 50460 8188
rect 50516 8186 50540 8188
rect 50378 8134 50380 8186
rect 50442 8134 50454 8186
rect 50516 8134 50518 8186
rect 50356 8132 50380 8134
rect 50436 8132 50460 8134
rect 50516 8132 50540 8134
rect 50300 8112 50596 8132
rect 50068 8084 50120 8090
rect 50068 8026 50120 8032
rect 50632 8022 50660 8230
rect 50620 8016 50672 8022
rect 50620 7958 50672 7964
rect 50160 7404 50212 7410
rect 50160 7346 50212 7352
rect 50172 7206 50200 7346
rect 50620 7336 50672 7342
rect 50620 7278 50672 7284
rect 50160 7200 50212 7206
rect 50160 7142 50212 7148
rect 50300 7100 50596 7120
rect 50356 7098 50380 7100
rect 50436 7098 50460 7100
rect 50516 7098 50540 7100
rect 50378 7046 50380 7098
rect 50442 7046 50454 7098
rect 50516 7046 50518 7098
rect 50356 7044 50380 7046
rect 50436 7044 50460 7046
rect 50516 7044 50540 7046
rect 50300 7024 50596 7044
rect 49976 6656 50028 6662
rect 49976 6598 50028 6604
rect 50436 6656 50488 6662
rect 50436 6598 50488 6604
rect 50448 6254 50476 6598
rect 50436 6248 50488 6254
rect 50172 6208 50436 6236
rect 50068 6180 50120 6186
rect 50068 6122 50120 6128
rect 50080 5846 50108 6122
rect 49976 5840 50028 5846
rect 49976 5782 50028 5788
rect 50068 5840 50120 5846
rect 50068 5782 50120 5788
rect 49988 5545 50016 5782
rect 49974 5536 50030 5545
rect 49974 5471 50030 5480
rect 49976 5092 50028 5098
rect 49976 5034 50028 5040
rect 49988 4826 50016 5034
rect 49976 4820 50028 4826
rect 49976 4762 50028 4768
rect 50080 4690 50108 5782
rect 50172 5778 50200 6208
rect 50436 6190 50488 6196
rect 50632 6118 50660 7278
rect 50724 7206 50752 9114
rect 50908 9110 50936 11614
rect 51000 10062 51028 12922
rect 51276 12850 51304 13806
rect 51368 13394 51396 14350
rect 51460 14346 51488 14826
rect 51448 14340 51500 14346
rect 51448 14282 51500 14288
rect 51540 13864 51592 13870
rect 51540 13806 51592 13812
rect 51356 13388 51408 13394
rect 51356 13330 51408 13336
rect 51264 12844 51316 12850
rect 51264 12786 51316 12792
rect 51172 12640 51224 12646
rect 51172 12582 51224 12588
rect 51184 12306 51212 12582
rect 51172 12300 51224 12306
rect 51172 12242 51224 12248
rect 51080 12232 51132 12238
rect 51080 12174 51132 12180
rect 51092 11898 51120 12174
rect 51080 11892 51132 11898
rect 51080 11834 51132 11840
rect 51184 11694 51212 12242
rect 51172 11688 51224 11694
rect 51172 11630 51224 11636
rect 51264 10464 51316 10470
rect 51264 10406 51316 10412
rect 51276 10198 51304 10406
rect 51264 10192 51316 10198
rect 51264 10134 51316 10140
rect 51172 10124 51224 10130
rect 51172 10066 51224 10072
rect 50988 10056 51040 10062
rect 50988 9998 51040 10004
rect 51000 9450 51028 9998
rect 51184 9722 51212 10066
rect 51172 9716 51224 9722
rect 51172 9658 51224 9664
rect 51368 9518 51396 13330
rect 51448 13320 51500 13326
rect 51448 13262 51500 13268
rect 51460 12986 51488 13262
rect 51448 12980 51500 12986
rect 51448 12922 51500 12928
rect 51552 12594 51580 13806
rect 51644 13802 51672 15982
rect 51908 15632 51960 15638
rect 51908 15574 51960 15580
rect 51920 15162 51948 15574
rect 52012 15570 52040 15982
rect 52000 15564 52052 15570
rect 52000 15506 52052 15512
rect 51908 15156 51960 15162
rect 51908 15098 51960 15104
rect 52000 15088 52052 15094
rect 52000 15030 52052 15036
rect 52012 14074 52040 15030
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 52092 13864 52144 13870
rect 52092 13806 52144 13812
rect 51632 13796 51684 13802
rect 51632 13738 51684 13744
rect 51460 12566 51580 12594
rect 51460 11218 51488 12566
rect 51540 11620 51592 11626
rect 51540 11562 51592 11568
rect 51552 11354 51580 11562
rect 51540 11348 51592 11354
rect 51540 11290 51592 11296
rect 51448 11212 51500 11218
rect 51448 11154 51500 11160
rect 51356 9512 51408 9518
rect 51356 9454 51408 9460
rect 50988 9444 51040 9450
rect 50988 9386 51040 9392
rect 51644 9110 51672 13738
rect 52000 13320 52052 13326
rect 52000 13262 52052 13268
rect 52012 12986 52040 13262
rect 52000 12980 52052 12986
rect 52000 12922 52052 12928
rect 51724 12776 51776 12782
rect 51724 12718 51776 12724
rect 51816 12776 51868 12782
rect 51816 12718 51868 12724
rect 51736 12306 51764 12718
rect 51828 12646 51856 12718
rect 51816 12640 51868 12646
rect 51816 12582 51868 12588
rect 51724 12300 51776 12306
rect 51724 12242 51776 12248
rect 51736 11898 51764 12242
rect 51828 12238 51856 12582
rect 52012 12442 52040 12922
rect 52000 12436 52052 12442
rect 52000 12378 52052 12384
rect 52000 12300 52052 12306
rect 52000 12242 52052 12248
rect 51816 12232 51868 12238
rect 51816 12174 51868 12180
rect 52012 11898 52040 12242
rect 51724 11892 51776 11898
rect 51724 11834 51776 11840
rect 52000 11892 52052 11898
rect 52000 11834 52052 11840
rect 52012 11218 52040 11834
rect 52000 11212 52052 11218
rect 52000 11154 52052 11160
rect 52104 11082 52132 13806
rect 52092 11076 52144 11082
rect 52092 11018 52144 11024
rect 52104 10690 52132 11018
rect 51920 10662 52132 10690
rect 51920 10606 51948 10662
rect 51908 10600 51960 10606
rect 52092 10600 52144 10606
rect 51908 10542 51960 10548
rect 52012 10560 52092 10588
rect 51816 9512 51868 9518
rect 51816 9454 51868 9460
rect 50896 9104 50948 9110
rect 50896 9046 50948 9052
rect 51632 9104 51684 9110
rect 51632 9046 51684 9052
rect 50804 9036 50856 9042
rect 50804 8978 50856 8984
rect 50816 8294 50844 8978
rect 51448 8968 51500 8974
rect 51448 8910 51500 8916
rect 51460 8566 51488 8910
rect 51448 8560 51500 8566
rect 51448 8502 51500 8508
rect 50804 8288 50856 8294
rect 50804 8230 50856 8236
rect 51264 8288 51316 8294
rect 51264 8230 51316 8236
rect 50816 7954 50844 8230
rect 51276 8022 51304 8230
rect 51264 8016 51316 8022
rect 51264 7958 51316 7964
rect 51356 8016 51408 8022
rect 51356 7958 51408 7964
rect 50804 7948 50856 7954
rect 50804 7890 50856 7896
rect 50988 7948 51040 7954
rect 50988 7890 51040 7896
rect 50816 7410 50844 7890
rect 50804 7404 50856 7410
rect 50804 7346 50856 7352
rect 50712 7200 50764 7206
rect 50712 7142 50764 7148
rect 50896 7200 50948 7206
rect 50896 7142 50948 7148
rect 50908 6866 50936 7142
rect 50896 6860 50948 6866
rect 50896 6802 50948 6808
rect 50804 6792 50856 6798
rect 51000 6769 51028 7890
rect 51368 7750 51396 7958
rect 51356 7744 51408 7750
rect 51356 7686 51408 7692
rect 51460 7546 51488 8502
rect 51828 8498 51856 9454
rect 52012 9178 52040 10560
rect 52196 10588 52224 27798
rect 52656 27418 52684 29038
rect 52748 28014 52776 29158
rect 52920 28484 52972 28490
rect 52920 28426 52972 28432
rect 52828 28144 52880 28150
rect 52828 28086 52880 28092
rect 52736 28008 52788 28014
rect 52736 27950 52788 27956
rect 52748 27606 52776 27950
rect 52840 27606 52868 28086
rect 52736 27600 52788 27606
rect 52736 27542 52788 27548
rect 52828 27600 52880 27606
rect 52828 27542 52880 27548
rect 52736 27464 52788 27470
rect 52656 27412 52736 27418
rect 52656 27406 52788 27412
rect 52656 27390 52776 27406
rect 52368 27328 52420 27334
rect 52368 27270 52420 27276
rect 52644 27328 52696 27334
rect 52644 27270 52696 27276
rect 52380 26994 52408 27270
rect 52368 26988 52420 26994
rect 52368 26930 52420 26936
rect 52656 26858 52684 27270
rect 52748 27062 52776 27390
rect 52828 27328 52880 27334
rect 52828 27270 52880 27276
rect 52736 27056 52788 27062
rect 52736 26998 52788 27004
rect 52644 26852 52696 26858
rect 52644 26794 52696 26800
rect 52460 26240 52512 26246
rect 52460 26182 52512 26188
rect 52472 25702 52500 26182
rect 52460 25696 52512 25702
rect 52460 25638 52512 25644
rect 52368 24676 52420 24682
rect 52368 24618 52420 24624
rect 52380 23866 52408 24618
rect 52460 24064 52512 24070
rect 52460 24006 52512 24012
rect 52368 23860 52420 23866
rect 52368 23802 52420 23808
rect 52472 23662 52500 24006
rect 52460 23656 52512 23662
rect 52460 23598 52512 23604
rect 52552 23656 52604 23662
rect 52552 23598 52604 23604
rect 52564 23526 52592 23598
rect 52552 23520 52604 23526
rect 52552 23462 52604 23468
rect 52368 22568 52420 22574
rect 52368 22510 52420 22516
rect 52276 22500 52328 22506
rect 52276 22442 52328 22448
rect 52288 20262 52316 22442
rect 52380 22166 52408 22510
rect 52368 22160 52420 22166
rect 52368 22102 52420 22108
rect 52564 22098 52592 23462
rect 52656 22506 52684 26794
rect 52840 26314 52868 27270
rect 52932 26489 52960 28426
rect 53024 28014 53052 30518
rect 53300 29782 53328 32302
rect 53484 30394 53512 33390
rect 53576 33114 53604 34478
rect 53564 33108 53616 33114
rect 53564 33050 53616 33056
rect 53656 32972 53708 32978
rect 53656 32914 53708 32920
rect 53668 32434 53696 32914
rect 53760 32434 53788 36790
rect 53852 36242 53880 36858
rect 54036 36718 54064 37062
rect 54864 36718 54892 37742
rect 54944 37732 54996 37738
rect 54944 37674 54996 37680
rect 54956 37466 54984 37674
rect 54944 37460 54996 37466
rect 54944 37402 54996 37408
rect 55140 37330 55168 40530
rect 55232 40497 55260 40598
rect 55218 40488 55274 40497
rect 55218 40423 55274 40432
rect 55220 39024 55272 39030
rect 55218 38992 55220 39001
rect 55272 38992 55274 39001
rect 55218 38927 55274 38936
rect 55220 37664 55272 37670
rect 55220 37606 55272 37612
rect 55232 37369 55260 37606
rect 55218 37360 55274 37369
rect 55128 37324 55180 37330
rect 55218 37295 55274 37304
rect 55128 37266 55180 37272
rect 54024 36712 54076 36718
rect 54024 36654 54076 36660
rect 54300 36712 54352 36718
rect 54300 36654 54352 36660
rect 54852 36712 54904 36718
rect 54852 36654 54904 36660
rect 54036 36310 54064 36654
rect 54116 36576 54168 36582
rect 54116 36518 54168 36524
rect 54024 36304 54076 36310
rect 54024 36246 54076 36252
rect 54128 36242 54156 36518
rect 53840 36236 53892 36242
rect 53840 36178 53892 36184
rect 54116 36236 54168 36242
rect 54116 36178 54168 36184
rect 53932 35624 53984 35630
rect 53932 35566 53984 35572
rect 53944 35290 53972 35566
rect 53932 35284 53984 35290
rect 53932 35226 53984 35232
rect 54312 35086 54340 36654
rect 54668 36644 54720 36650
rect 54668 36586 54720 36592
rect 54680 36378 54708 36586
rect 54852 36576 54904 36582
rect 54852 36518 54904 36524
rect 54668 36372 54720 36378
rect 54668 36314 54720 36320
rect 54864 36038 54892 36518
rect 54852 36032 54904 36038
rect 54852 35974 54904 35980
rect 54944 36032 54996 36038
rect 54944 35974 54996 35980
rect 54392 35488 54444 35494
rect 54390 35456 54392 35465
rect 54444 35456 54446 35465
rect 54390 35391 54446 35400
rect 54956 35193 54984 35974
rect 55140 35494 55168 37266
rect 55218 35864 55274 35873
rect 55218 35799 55220 35808
rect 55272 35799 55274 35808
rect 55220 35770 55272 35776
rect 55128 35488 55180 35494
rect 55128 35430 55180 35436
rect 54942 35184 54998 35193
rect 54392 35148 54444 35154
rect 54444 35108 54616 35136
rect 54942 35119 54998 35128
rect 55036 35148 55088 35154
rect 54392 35090 54444 35096
rect 53840 35080 53892 35086
rect 53840 35022 53892 35028
rect 54300 35080 54352 35086
rect 54300 35022 54352 35028
rect 53852 33998 53880 35022
rect 54208 34944 54260 34950
rect 54208 34886 54260 34892
rect 54300 34944 54352 34950
rect 54300 34886 54352 34892
rect 54220 34542 54248 34886
rect 54312 34746 54340 34886
rect 54300 34740 54352 34746
rect 54300 34682 54352 34688
rect 54588 34542 54616 35108
rect 54956 34678 54984 35119
rect 55036 35090 55088 35096
rect 55048 34746 55076 35090
rect 55036 34740 55088 34746
rect 55036 34682 55088 34688
rect 55128 34740 55180 34746
rect 55128 34682 55180 34688
rect 54944 34672 54996 34678
rect 54944 34614 54996 34620
rect 54668 34604 54720 34610
rect 54668 34546 54720 34552
rect 54852 34604 54904 34610
rect 54852 34546 54904 34552
rect 54208 34536 54260 34542
rect 54208 34478 54260 34484
rect 54576 34536 54628 34542
rect 54576 34478 54628 34484
rect 54588 34377 54616 34478
rect 54574 34368 54630 34377
rect 54574 34303 54630 34312
rect 53840 33992 53892 33998
rect 53840 33934 53892 33940
rect 53656 32428 53708 32434
rect 53656 32370 53708 32376
rect 53748 32428 53800 32434
rect 53748 32370 53800 32376
rect 53852 31929 53880 33934
rect 54392 33584 54444 33590
rect 54444 33544 54616 33572
rect 54680 33561 54708 34546
rect 54864 34474 54892 34546
rect 54852 34468 54904 34474
rect 54852 34410 54904 34416
rect 55140 33862 55168 34682
rect 55218 34232 55274 34241
rect 55218 34167 55274 34176
rect 55232 34134 55260 34167
rect 55220 34128 55272 34134
rect 55220 34070 55272 34076
rect 55324 33946 55352 54674
rect 55508 54670 55536 55558
rect 55784 54874 55812 55762
rect 56140 55072 56192 55078
rect 56140 55014 56192 55020
rect 55772 54868 55824 54874
rect 55772 54810 55824 54816
rect 56152 54738 56180 55014
rect 56244 54806 56272 56374
rect 56520 55758 56548 57967
rect 56600 57044 56652 57050
rect 56600 56986 56652 56992
rect 56612 56506 56640 56986
rect 56876 56772 56928 56778
rect 56876 56714 56928 56720
rect 57060 56772 57112 56778
rect 57060 56714 57112 56720
rect 56600 56500 56652 56506
rect 56600 56442 56652 56448
rect 56888 56370 56916 56714
rect 57072 56545 57100 56714
rect 57058 56536 57114 56545
rect 57058 56471 57114 56480
rect 56876 56364 56928 56370
rect 56876 56306 56928 56312
rect 57164 56234 57192 59200
rect 57992 57474 58020 59200
rect 57992 57446 58296 57474
rect 57980 57316 58032 57322
rect 57980 57258 58032 57264
rect 58164 57316 58216 57322
rect 58164 57258 58216 57264
rect 57992 57050 58020 57258
rect 58072 57248 58124 57254
rect 58072 57190 58124 57196
rect 57980 57044 58032 57050
rect 57980 56986 58032 56992
rect 57980 56908 58032 56914
rect 57980 56850 58032 56856
rect 57612 56840 57664 56846
rect 57612 56782 57664 56788
rect 57152 56228 57204 56234
rect 57152 56170 57204 56176
rect 57624 55962 57652 56782
rect 57704 56704 57756 56710
rect 57704 56646 57756 56652
rect 57716 56370 57744 56646
rect 57704 56364 57756 56370
rect 57704 56306 57756 56312
rect 57612 55956 57664 55962
rect 57612 55898 57664 55904
rect 57336 55820 57388 55826
rect 57336 55762 57388 55768
rect 56508 55752 56560 55758
rect 56508 55694 56560 55700
rect 57244 55276 57296 55282
rect 57244 55218 57296 55224
rect 56324 55208 56376 55214
rect 56324 55150 56376 55156
rect 56600 55208 56652 55214
rect 56600 55150 56652 55156
rect 56336 54874 56364 55150
rect 56324 54868 56376 54874
rect 56324 54810 56376 54816
rect 56232 54800 56284 54806
rect 56232 54742 56284 54748
rect 56140 54732 56192 54738
rect 56140 54674 56192 54680
rect 55496 54664 55548 54670
rect 55496 54606 55548 54612
rect 56324 54596 56376 54602
rect 56324 54538 56376 54544
rect 55494 54496 55550 54505
rect 55494 54431 55550 54440
rect 55508 54126 55536 54431
rect 56336 54126 56364 54538
rect 56612 54330 56640 55150
rect 56876 55140 56928 55146
rect 56876 55082 56928 55088
rect 57060 55140 57112 55146
rect 57060 55082 57112 55088
rect 56888 54330 56916 55082
rect 57072 54913 57100 55082
rect 57058 54904 57114 54913
rect 57058 54839 57114 54848
rect 56600 54324 56652 54330
rect 56600 54266 56652 54272
rect 56876 54324 56928 54330
rect 56876 54266 56928 54272
rect 57256 54194 57284 55218
rect 57348 54874 57376 55762
rect 57992 55214 58020 56850
rect 58084 56506 58112 57190
rect 58176 57089 58204 57258
rect 58162 57080 58218 57089
rect 58162 57015 58218 57024
rect 58072 56500 58124 56506
rect 58072 56442 58124 56448
rect 58268 56438 58296 57446
rect 58256 56432 58308 56438
rect 58256 56374 58308 56380
rect 58256 55888 58308 55894
rect 58256 55830 58308 55836
rect 58164 55684 58216 55690
rect 58164 55626 58216 55632
rect 58176 55457 58204 55626
rect 58162 55448 58218 55457
rect 58162 55383 58218 55392
rect 57980 55208 58032 55214
rect 57980 55150 58032 55156
rect 57336 54868 57388 54874
rect 57336 54810 57388 54816
rect 57980 54732 58032 54738
rect 57980 54674 58032 54680
rect 57244 54188 57296 54194
rect 57244 54130 57296 54136
rect 55496 54120 55548 54126
rect 55496 54062 55548 54068
rect 56324 54120 56376 54126
rect 56324 54062 56376 54068
rect 55588 53644 55640 53650
rect 55588 53586 55640 53592
rect 55600 52873 55628 53586
rect 56336 53038 56364 54062
rect 57428 54052 57480 54058
rect 57428 53994 57480 54000
rect 56968 53984 57020 53990
rect 56968 53926 57020 53932
rect 56416 53576 56468 53582
rect 56416 53518 56468 53524
rect 56428 53242 56456 53518
rect 56980 53417 57008 53926
rect 57244 53576 57296 53582
rect 57244 53518 57296 53524
rect 56966 53408 57022 53417
rect 56966 53343 57022 53352
rect 57256 53242 57284 53518
rect 57440 53514 57468 53994
rect 57428 53508 57480 53514
rect 57428 53450 57480 53456
rect 57992 53242 58020 54674
rect 58164 54596 58216 54602
rect 58164 54538 58216 54544
rect 58176 53961 58204 54538
rect 58162 53952 58218 53961
rect 58162 53887 58218 53896
rect 56416 53236 56468 53242
rect 56416 53178 56468 53184
rect 57244 53236 57296 53242
rect 57244 53178 57296 53184
rect 57980 53236 58032 53242
rect 57980 53178 58032 53184
rect 56324 53032 56376 53038
rect 56324 52974 56376 52980
rect 57244 53032 57296 53038
rect 57244 52974 57296 52980
rect 55586 52864 55642 52873
rect 55586 52799 55642 52808
rect 55496 51944 55548 51950
rect 55496 51886 55548 51892
rect 55508 51377 55536 51886
rect 55494 51368 55550 51377
rect 55494 51303 55550 51312
rect 56336 50862 56364 52974
rect 57256 52698 57284 52974
rect 57244 52692 57296 52698
rect 57244 52634 57296 52640
rect 57428 52556 57480 52562
rect 57428 52498 57480 52504
rect 57980 52556 58032 52562
rect 57980 52498 58032 52504
rect 57058 51912 57114 51921
rect 56876 51876 56928 51882
rect 57440 51882 57468 52498
rect 57888 52488 57940 52494
rect 57888 52430 57940 52436
rect 57900 52329 57928 52430
rect 57886 52320 57942 52329
rect 57886 52255 57942 52264
rect 57992 52154 58020 52498
rect 57980 52148 58032 52154
rect 57980 52090 58032 52096
rect 57520 51944 57572 51950
rect 57520 51886 57572 51892
rect 57058 51847 57060 51856
rect 56876 51818 56928 51824
rect 57112 51847 57114 51856
rect 57428 51876 57480 51882
rect 57060 51818 57112 51824
rect 57428 51818 57480 51824
rect 56888 51610 56916 51818
rect 56876 51604 56928 51610
rect 56876 51546 56928 51552
rect 57244 51400 57296 51406
rect 57244 51342 57296 51348
rect 57256 51066 57284 51342
rect 57244 51060 57296 51066
rect 57244 51002 57296 51008
rect 57440 50862 57468 51818
rect 57532 51474 57560 51886
rect 57520 51468 57572 51474
rect 57520 51410 57572 51416
rect 56324 50856 56376 50862
rect 56324 50798 56376 50804
rect 57428 50856 57480 50862
rect 57428 50798 57480 50804
rect 58162 50824 58218 50833
rect 56336 49978 56364 50798
rect 56876 50380 56928 50386
rect 56876 50322 56928 50328
rect 56888 49978 56916 50322
rect 57058 50280 57114 50289
rect 57058 50215 57060 50224
rect 57112 50215 57114 50224
rect 57060 50186 57112 50192
rect 57152 50176 57204 50182
rect 57152 50118 57204 50124
rect 56324 49972 56376 49978
rect 56324 49914 56376 49920
rect 56876 49972 56928 49978
rect 56876 49914 56928 49920
rect 55956 49836 56008 49842
rect 55956 49778 56008 49784
rect 55772 49088 55824 49094
rect 55772 49030 55824 49036
rect 55784 48754 55812 49030
rect 55772 48748 55824 48754
rect 55772 48690 55824 48696
rect 55496 48680 55548 48686
rect 55496 48622 55548 48628
rect 55508 48249 55536 48622
rect 55494 48240 55550 48249
rect 55494 48175 55550 48184
rect 55496 48136 55548 48142
rect 55496 48078 55548 48084
rect 55508 47802 55536 48078
rect 55496 47796 55548 47802
rect 55496 47738 55548 47744
rect 55680 47592 55732 47598
rect 55680 47534 55732 47540
rect 55692 46918 55720 47534
rect 55968 47122 55996 49778
rect 56336 49774 56364 49914
rect 57164 49842 57192 50118
rect 57152 49836 57204 49842
rect 57152 49778 57204 49784
rect 56324 49768 56376 49774
rect 56324 49710 56376 49716
rect 57440 49298 57468 50798
rect 57520 50788 57572 50794
rect 57520 50730 57572 50736
rect 57980 50788 58032 50794
rect 58162 50759 58164 50768
rect 57980 50730 58032 50736
rect 58216 50759 58218 50768
rect 58164 50730 58216 50736
rect 57532 50386 57560 50730
rect 57704 50720 57756 50726
rect 57704 50662 57756 50668
rect 57716 50386 57744 50662
rect 57992 50522 58020 50730
rect 57980 50516 58032 50522
rect 57980 50458 58032 50464
rect 57520 50380 57572 50386
rect 57520 50322 57572 50328
rect 57704 50380 57756 50386
rect 57704 50322 57756 50328
rect 58162 49328 58218 49337
rect 57428 49292 57480 49298
rect 57428 49234 57480 49240
rect 57796 49292 57848 49298
rect 57796 49234 57848 49240
rect 57980 49292 58032 49298
rect 58162 49263 58164 49272
rect 57980 49234 58032 49240
rect 58216 49263 58218 49272
rect 58164 49234 58216 49240
rect 57704 49088 57756 49094
rect 57704 49030 57756 49036
rect 57060 48816 57112 48822
rect 57058 48784 57060 48793
rect 57112 48784 57114 48793
rect 57716 48754 57744 49030
rect 57058 48719 57114 48728
rect 57704 48748 57756 48754
rect 57704 48690 57756 48696
rect 57060 48680 57112 48686
rect 57060 48622 57112 48628
rect 57072 48210 57100 48622
rect 57428 48612 57480 48618
rect 57428 48554 57480 48560
rect 57060 48204 57112 48210
rect 57060 48146 57112 48152
rect 57440 48074 57468 48554
rect 57428 48068 57480 48074
rect 57428 48010 57480 48016
rect 57520 48000 57572 48006
rect 57520 47942 57572 47948
rect 57058 47696 57114 47705
rect 57532 47666 57560 47942
rect 57058 47631 57060 47640
rect 57112 47631 57114 47640
rect 57520 47660 57572 47666
rect 57060 47602 57112 47608
rect 57520 47602 57572 47608
rect 57808 47598 57836 49234
rect 57992 48890 58020 49234
rect 57980 48884 58032 48890
rect 57980 48826 58032 48832
rect 57796 47592 57848 47598
rect 57796 47534 57848 47540
rect 57426 47152 57482 47161
rect 55956 47116 56008 47122
rect 55956 47058 56008 47064
rect 57244 47116 57296 47122
rect 57426 47087 57428 47096
rect 57244 47058 57296 47064
rect 57480 47087 57482 47096
rect 57428 47058 57480 47064
rect 55680 46912 55732 46918
rect 55680 46854 55732 46860
rect 55692 46510 55720 46854
rect 55680 46504 55732 46510
rect 55680 46446 55732 46452
rect 55692 45422 55720 46446
rect 55968 46034 55996 47058
rect 57256 46714 57284 47058
rect 57520 46980 57572 46986
rect 57520 46922 57572 46928
rect 57244 46708 57296 46714
rect 57244 46650 57296 46656
rect 55772 46028 55824 46034
rect 55772 45970 55824 45976
rect 55956 46028 56008 46034
rect 55956 45970 56008 45976
rect 55784 45898 55812 45970
rect 55772 45892 55824 45898
rect 55772 45834 55824 45840
rect 55680 45416 55732 45422
rect 55680 45358 55732 45364
rect 55404 45280 55456 45286
rect 55404 45222 55456 45228
rect 55416 43858 55444 45222
rect 55588 44940 55640 44946
rect 55588 44882 55640 44888
rect 55600 44470 55628 44882
rect 55588 44464 55640 44470
rect 55588 44406 55640 44412
rect 55404 43852 55456 43858
rect 55404 43794 55456 43800
rect 55692 43722 55720 45358
rect 55680 43716 55732 43722
rect 55680 43658 55732 43664
rect 55404 42696 55456 42702
rect 55404 42638 55456 42644
rect 55416 42362 55444 42638
rect 55404 42356 55456 42362
rect 55404 42298 55456 42304
rect 55404 42084 55456 42090
rect 55404 42026 55456 42032
rect 55416 41818 55444 42026
rect 55404 41812 55456 41818
rect 55404 41754 55456 41760
rect 55496 40588 55548 40594
rect 55496 40530 55548 40536
rect 55404 40384 55456 40390
rect 55404 40326 55456 40332
rect 55416 39982 55444 40326
rect 55404 39976 55456 39982
rect 55404 39918 55456 39924
rect 55508 39846 55536 40530
rect 55588 40452 55640 40458
rect 55588 40394 55640 40400
rect 55496 39840 55548 39846
rect 55496 39782 55548 39788
rect 55508 39642 55536 39782
rect 55496 39636 55548 39642
rect 55496 39578 55548 39584
rect 55508 38894 55536 39578
rect 55600 39098 55628 40394
rect 55588 39092 55640 39098
rect 55588 39034 55640 39040
rect 55496 38888 55548 38894
rect 55496 38830 55548 38836
rect 55588 38344 55640 38350
rect 55588 38286 55640 38292
rect 55600 38214 55628 38286
rect 55588 38208 55640 38214
rect 55588 38150 55640 38156
rect 55496 37732 55548 37738
rect 55496 37674 55548 37680
rect 55508 37466 55536 37674
rect 55496 37460 55548 37466
rect 55496 37402 55548 37408
rect 55600 37330 55628 38150
rect 55588 37324 55640 37330
rect 55588 37266 55640 37272
rect 55404 36304 55456 36310
rect 55404 36246 55456 36252
rect 55416 35562 55444 36246
rect 55588 36236 55640 36242
rect 55588 36178 55640 36184
rect 55404 35556 55456 35562
rect 55404 35498 55456 35504
rect 55416 34474 55444 35498
rect 55600 34950 55628 36178
rect 55588 34944 55640 34950
rect 55588 34886 55640 34892
rect 55404 34468 55456 34474
rect 55404 34410 55456 34416
rect 55494 34368 55550 34377
rect 55494 34303 55550 34312
rect 55232 33918 55352 33946
rect 55404 33924 55456 33930
rect 55128 33856 55180 33862
rect 54758 33824 54814 33833
rect 55128 33798 55180 33804
rect 54758 33759 54814 33768
rect 54392 33526 54444 33532
rect 54392 33448 54444 33454
rect 54588 33436 54616 33544
rect 54666 33552 54722 33561
rect 54772 33522 54800 33759
rect 54666 33487 54722 33496
rect 54760 33516 54812 33522
rect 54760 33458 54812 33464
rect 54668 33448 54720 33454
rect 54588 33408 54668 33436
rect 54392 33390 54444 33396
rect 54668 33390 54720 33396
rect 54300 33108 54352 33114
rect 54300 33050 54352 33056
rect 54116 33040 54168 33046
rect 54116 32982 54168 32988
rect 54024 32836 54076 32842
rect 54024 32778 54076 32784
rect 53838 31920 53894 31929
rect 53838 31855 53894 31864
rect 53654 30832 53710 30841
rect 53654 30767 53656 30776
rect 53708 30767 53710 30776
rect 53838 30832 53894 30841
rect 53838 30767 53840 30776
rect 53656 30738 53708 30744
rect 53892 30767 53894 30776
rect 53840 30738 53892 30744
rect 53472 30388 53524 30394
rect 53472 30330 53524 30336
rect 54036 30258 54064 32778
rect 54128 32230 54156 32982
rect 54312 32978 54340 33050
rect 54300 32972 54352 32978
rect 54300 32914 54352 32920
rect 54300 32768 54352 32774
rect 54300 32710 54352 32716
rect 54312 32434 54340 32710
rect 54300 32428 54352 32434
rect 54300 32370 54352 32376
rect 54116 32224 54168 32230
rect 54116 32166 54168 32172
rect 54300 32224 54352 32230
rect 54300 32166 54352 32172
rect 54312 31958 54340 32166
rect 54300 31952 54352 31958
rect 54300 31894 54352 31900
rect 54404 31686 54432 33390
rect 55036 33312 55088 33318
rect 55036 33254 55088 33260
rect 54588 32966 54800 32994
rect 54484 32836 54536 32842
rect 54588 32824 54616 32966
rect 54772 32842 54800 32966
rect 54536 32796 54616 32824
rect 54760 32836 54812 32842
rect 54484 32778 54536 32784
rect 54760 32778 54812 32784
rect 54852 32768 54904 32774
rect 54904 32716 54984 32722
rect 54852 32710 54984 32716
rect 54864 32694 54984 32710
rect 54956 32502 54984 32694
rect 54944 32496 54996 32502
rect 54944 32438 54996 32444
rect 54484 32020 54536 32026
rect 54484 31962 54536 31968
rect 54392 31680 54444 31686
rect 54392 31622 54444 31628
rect 54404 31482 54432 31622
rect 54392 31476 54444 31482
rect 54392 31418 54444 31424
rect 54496 30802 54524 31962
rect 54956 31906 54984 32438
rect 55048 32434 55076 33254
rect 55128 33108 55180 33114
rect 55128 33050 55180 33056
rect 55036 32428 55088 32434
rect 55036 32370 55088 32376
rect 55140 31958 55168 33050
rect 54772 31890 54984 31906
rect 55128 31952 55180 31958
rect 55128 31894 55180 31900
rect 54576 31884 54628 31890
rect 54576 31826 54628 31832
rect 54772 31884 54996 31890
rect 54772 31878 54944 31884
rect 54588 31754 54616 31826
rect 54576 31748 54628 31754
rect 54576 31690 54628 31696
rect 54588 30802 54616 31690
rect 54668 31680 54720 31686
rect 54668 31622 54720 31628
rect 54680 31278 54708 31622
rect 54772 31482 54800 31878
rect 54944 31826 54996 31832
rect 55140 31754 55168 31894
rect 54864 31726 55168 31754
rect 54760 31476 54812 31482
rect 54760 31418 54812 31424
rect 54864 31278 54892 31726
rect 55232 31634 55260 33918
rect 55404 33866 55456 33872
rect 55416 33833 55444 33866
rect 55402 33824 55458 33833
rect 55402 33759 55458 33768
rect 55508 33454 55536 34303
rect 55600 33658 55628 34886
rect 55588 33652 55640 33658
rect 55588 33594 55640 33600
rect 55600 33561 55628 33594
rect 55586 33552 55642 33561
rect 55586 33487 55642 33496
rect 55496 33448 55548 33454
rect 55496 33390 55548 33396
rect 55496 32836 55548 32842
rect 55496 32778 55548 32784
rect 55404 32292 55456 32298
rect 55404 32234 55456 32240
rect 55140 31606 55260 31634
rect 54668 31272 54720 31278
rect 54668 31214 54720 31220
rect 54852 31272 54904 31278
rect 54852 31214 54904 31220
rect 54944 31272 54996 31278
rect 54944 31214 54996 31220
rect 54758 30832 54814 30841
rect 54484 30796 54536 30802
rect 54484 30738 54536 30744
rect 54576 30796 54628 30802
rect 54758 30767 54760 30776
rect 54576 30738 54628 30744
rect 54812 30767 54814 30776
rect 54760 30738 54812 30744
rect 54208 30660 54260 30666
rect 54208 30602 54260 30608
rect 54024 30252 54076 30258
rect 54024 30194 54076 30200
rect 54220 30190 54248 30602
rect 54496 30274 54524 30738
rect 54772 30394 54800 30738
rect 54760 30388 54812 30394
rect 54760 30330 54812 30336
rect 54496 30246 54708 30274
rect 54680 30190 54708 30246
rect 54208 30184 54260 30190
rect 54208 30126 54260 30132
rect 54668 30184 54720 30190
rect 54668 30126 54720 30132
rect 54116 30048 54168 30054
rect 54116 29990 54168 29996
rect 53288 29776 53340 29782
rect 53288 29718 53340 29724
rect 54024 29708 54076 29714
rect 54024 29650 54076 29656
rect 53748 29572 53800 29578
rect 53748 29514 53800 29520
rect 53760 29170 53788 29514
rect 54036 29306 54064 29650
rect 54024 29300 54076 29306
rect 54024 29242 54076 29248
rect 53748 29164 53800 29170
rect 53748 29106 53800 29112
rect 53472 29096 53524 29102
rect 53472 29038 53524 29044
rect 53196 28552 53248 28558
rect 53196 28494 53248 28500
rect 53012 28008 53064 28014
rect 53012 27950 53064 27956
rect 53024 27402 53052 27950
rect 53208 27402 53236 28494
rect 53484 27878 53512 29038
rect 53472 27872 53524 27878
rect 53472 27814 53524 27820
rect 53484 27674 53512 27814
rect 53472 27668 53524 27674
rect 53472 27610 53524 27616
rect 53012 27396 53064 27402
rect 53012 27338 53064 27344
rect 53196 27396 53248 27402
rect 53196 27338 53248 27344
rect 53208 26926 53236 27338
rect 53012 26920 53064 26926
rect 53012 26862 53064 26868
rect 53196 26920 53248 26926
rect 53196 26862 53248 26868
rect 53024 26790 53052 26862
rect 53012 26784 53064 26790
rect 53012 26726 53064 26732
rect 52918 26480 52974 26489
rect 52918 26415 52920 26424
rect 52972 26415 52974 26424
rect 52920 26386 52972 26392
rect 52828 26308 52880 26314
rect 52828 26250 52880 26256
rect 52736 25900 52788 25906
rect 52736 25842 52788 25848
rect 52748 25158 52776 25842
rect 53656 25220 53708 25226
rect 53656 25162 53708 25168
rect 52736 25152 52788 25158
rect 52736 25094 52788 25100
rect 53668 24954 53696 25162
rect 53656 24948 53708 24954
rect 53656 24890 53708 24896
rect 53760 24834 53788 29106
rect 54128 29102 54156 29990
rect 54864 29714 54892 31214
rect 54956 29782 54984 31214
rect 55140 31090 55168 31606
rect 55218 31240 55274 31249
rect 55218 31175 55220 31184
rect 55272 31175 55274 31184
rect 55220 31146 55272 31152
rect 55140 31062 55260 31090
rect 55128 30388 55180 30394
rect 55128 30330 55180 30336
rect 55140 30258 55168 30330
rect 55128 30252 55180 30258
rect 55128 30194 55180 30200
rect 54944 29776 54996 29782
rect 54944 29718 54996 29724
rect 54852 29708 54904 29714
rect 54852 29650 54904 29656
rect 54208 29640 54260 29646
rect 54208 29582 54260 29588
rect 54116 29096 54168 29102
rect 54116 29038 54168 29044
rect 54220 28422 54248 29582
rect 54956 29186 54984 29718
rect 54956 29158 55076 29186
rect 54944 29096 54996 29102
rect 54944 29038 54996 29044
rect 54208 28416 54260 28422
rect 54208 28358 54260 28364
rect 54300 28416 54352 28422
rect 54300 28358 54352 28364
rect 54208 28144 54260 28150
rect 54208 28086 54260 28092
rect 54024 27872 54076 27878
rect 54024 27814 54076 27820
rect 53932 26852 53984 26858
rect 53932 26794 53984 26800
rect 53668 24818 53880 24834
rect 53668 24812 53892 24818
rect 53668 24806 53840 24812
rect 53012 24336 53064 24342
rect 53012 24278 53064 24284
rect 52828 24200 52880 24206
rect 52828 24142 52880 24148
rect 52736 23656 52788 23662
rect 52736 23598 52788 23604
rect 52748 22817 52776 23598
rect 52734 22808 52790 22817
rect 52734 22743 52790 22752
rect 52748 22574 52776 22743
rect 52736 22568 52788 22574
rect 52736 22510 52788 22516
rect 52644 22500 52696 22506
rect 52644 22442 52696 22448
rect 52840 22098 52868 24142
rect 53024 23866 53052 24278
rect 53012 23860 53064 23866
rect 53012 23802 53064 23808
rect 53668 23526 53696 24806
rect 53840 24754 53892 24760
rect 53944 24750 53972 26794
rect 54036 26790 54064 27814
rect 54220 27577 54248 28086
rect 54206 27568 54262 27577
rect 54312 27538 54340 28358
rect 54668 28076 54720 28082
rect 54668 28018 54720 28024
rect 54680 27538 54708 28018
rect 54206 27503 54262 27512
rect 54300 27532 54352 27538
rect 54220 27470 54248 27503
rect 54300 27474 54352 27480
rect 54668 27532 54720 27538
rect 54668 27474 54720 27480
rect 54116 27464 54168 27470
rect 54116 27406 54168 27412
rect 54208 27464 54260 27470
rect 54208 27406 54260 27412
rect 54128 27130 54156 27406
rect 54116 27124 54168 27130
rect 54116 27066 54168 27072
rect 54208 26988 54260 26994
rect 54208 26930 54260 26936
rect 54024 26784 54076 26790
rect 54024 26726 54076 26732
rect 54116 26444 54168 26450
rect 54116 26386 54168 26392
rect 54128 24818 54156 26386
rect 54220 26382 54248 26930
rect 54312 26858 54340 27474
rect 54576 27464 54628 27470
rect 54576 27406 54628 27412
rect 54300 26852 54352 26858
rect 54300 26794 54352 26800
rect 54588 26790 54616 27406
rect 54576 26784 54628 26790
rect 54576 26726 54628 26732
rect 54300 26580 54352 26586
rect 54300 26522 54352 26528
rect 54208 26376 54260 26382
rect 54208 26318 54260 26324
rect 54312 25838 54340 26522
rect 54392 26444 54444 26450
rect 54392 26386 54444 26392
rect 54300 25832 54352 25838
rect 54300 25774 54352 25780
rect 54404 25702 54432 26386
rect 54852 26376 54904 26382
rect 54852 26318 54904 26324
rect 54760 25832 54812 25838
rect 54760 25774 54812 25780
rect 54392 25696 54444 25702
rect 54392 25638 54444 25644
rect 54404 25430 54432 25638
rect 54392 25424 54444 25430
rect 54392 25366 54444 25372
rect 54772 24818 54800 25774
rect 54864 25770 54892 26318
rect 54852 25764 54904 25770
rect 54852 25706 54904 25712
rect 54956 25362 54984 29038
rect 55048 28014 55076 29158
rect 55232 29152 55260 31062
rect 55416 30938 55444 32234
rect 55404 30932 55456 30938
rect 55404 30874 55456 30880
rect 55508 30802 55536 32778
rect 55680 31204 55732 31210
rect 55680 31146 55732 31152
rect 55312 30796 55364 30802
rect 55312 30738 55364 30744
rect 55496 30796 55548 30802
rect 55496 30738 55548 30744
rect 55324 30190 55352 30738
rect 55692 30394 55720 31146
rect 55680 30388 55732 30394
rect 55680 30330 55732 30336
rect 55312 30184 55364 30190
rect 55312 30126 55364 30132
rect 55494 29608 55550 29617
rect 55494 29543 55550 29552
rect 55508 29238 55536 29543
rect 55496 29232 55548 29238
rect 55496 29174 55548 29180
rect 55232 29124 55444 29152
rect 55128 29096 55180 29102
rect 55128 29038 55180 29044
rect 55140 28762 55168 29038
rect 55220 29028 55272 29034
rect 55220 28970 55272 28976
rect 55128 28756 55180 28762
rect 55128 28698 55180 28704
rect 55140 28150 55168 28698
rect 55128 28144 55180 28150
rect 55128 28086 55180 28092
rect 55232 28014 55260 28970
rect 55312 28688 55364 28694
rect 55312 28630 55364 28636
rect 55324 28121 55352 28630
rect 55310 28112 55366 28121
rect 55310 28047 55366 28056
rect 55036 28008 55088 28014
rect 55220 28008 55272 28014
rect 55088 27968 55168 27996
rect 55036 27950 55088 27956
rect 55036 26852 55088 26858
rect 55036 26794 55088 26800
rect 55048 26586 55076 26794
rect 55036 26580 55088 26586
rect 55036 26522 55088 26528
rect 55140 25888 55168 27968
rect 55220 27950 55272 27956
rect 55220 27600 55272 27606
rect 55220 27542 55272 27548
rect 55232 26994 55260 27542
rect 55312 27532 55364 27538
rect 55312 27474 55364 27480
rect 55220 26988 55272 26994
rect 55220 26930 55272 26936
rect 55324 26926 55352 27474
rect 55312 26920 55364 26926
rect 55312 26862 55364 26868
rect 55220 26852 55272 26858
rect 55220 26794 55272 26800
rect 55232 26518 55260 26794
rect 55220 26512 55272 26518
rect 55220 26454 55272 26460
rect 55324 26246 55352 26862
rect 55312 26240 55364 26246
rect 55312 26182 55364 26188
rect 55048 25860 55168 25888
rect 55048 25770 55076 25860
rect 55036 25764 55088 25770
rect 55036 25706 55088 25712
rect 55128 25764 55180 25770
rect 55128 25706 55180 25712
rect 55312 25764 55364 25770
rect 55312 25706 55364 25712
rect 55140 25498 55168 25706
rect 55128 25492 55180 25498
rect 55128 25434 55180 25440
rect 54944 25356 54996 25362
rect 54944 25298 54996 25304
rect 54116 24812 54168 24818
rect 54116 24754 54168 24760
rect 54760 24812 54812 24818
rect 54760 24754 54812 24760
rect 53932 24744 53984 24750
rect 53932 24686 53984 24692
rect 54852 24676 54904 24682
rect 54956 24664 54984 25298
rect 55324 25294 55352 25706
rect 55312 25288 55364 25294
rect 55312 25230 55364 25236
rect 55218 24984 55274 24993
rect 55218 24919 55220 24928
rect 55272 24919 55274 24928
rect 55220 24890 55272 24896
rect 54904 24636 54984 24664
rect 54852 24618 54904 24624
rect 53748 24608 53800 24614
rect 53748 24550 53800 24556
rect 54208 24608 54260 24614
rect 54208 24550 54260 24556
rect 53760 24274 53788 24550
rect 53748 24268 53800 24274
rect 53748 24210 53800 24216
rect 54220 24206 54248 24550
rect 54576 24404 54628 24410
rect 54576 24346 54628 24352
rect 54588 24274 54616 24346
rect 54668 24336 54720 24342
rect 54668 24278 54720 24284
rect 54576 24268 54628 24274
rect 54576 24210 54628 24216
rect 54208 24200 54260 24206
rect 54208 24142 54260 24148
rect 54392 23656 54444 23662
rect 54392 23598 54444 23604
rect 54484 23656 54536 23662
rect 54484 23598 54536 23604
rect 53656 23520 53708 23526
rect 53656 23462 53708 23468
rect 54208 23180 54260 23186
rect 54208 23122 54260 23128
rect 53840 23044 53892 23050
rect 53840 22986 53892 22992
rect 53748 22772 53800 22778
rect 53748 22714 53800 22720
rect 53760 22642 53788 22714
rect 53748 22636 53800 22642
rect 53748 22578 53800 22584
rect 53380 22432 53432 22438
rect 53380 22374 53432 22380
rect 52552 22092 52604 22098
rect 52552 22034 52604 22040
rect 52828 22092 52880 22098
rect 52828 22034 52880 22040
rect 52564 21078 52592 22034
rect 52644 21888 52696 21894
rect 52644 21830 52696 21836
rect 52552 21072 52604 21078
rect 52656 21049 52684 21830
rect 53392 21690 53420 22374
rect 53196 21684 53248 21690
rect 53196 21626 53248 21632
rect 53380 21684 53432 21690
rect 53380 21626 53432 21632
rect 52736 21616 52788 21622
rect 52920 21616 52972 21622
rect 52788 21564 52920 21570
rect 52736 21558 52972 21564
rect 52748 21542 52960 21558
rect 52736 21480 52788 21486
rect 52736 21422 52788 21428
rect 52552 21014 52604 21020
rect 52642 21040 52698 21049
rect 52642 20975 52644 20984
rect 52696 20975 52698 20984
rect 52644 20946 52696 20952
rect 52552 20936 52604 20942
rect 52656 20915 52684 20946
rect 52748 20942 52776 21422
rect 52920 21004 52972 21010
rect 52840 20964 52920 20992
rect 52736 20936 52788 20942
rect 52552 20878 52604 20884
rect 52736 20878 52788 20884
rect 52564 20346 52592 20878
rect 52840 20466 52868 20964
rect 52920 20946 52972 20952
rect 53104 20936 53156 20942
rect 53104 20878 53156 20884
rect 52920 20800 52972 20806
rect 52920 20742 52972 20748
rect 52828 20460 52880 20466
rect 52748 20420 52828 20448
rect 52564 20318 52684 20346
rect 52276 20256 52328 20262
rect 52276 20198 52328 20204
rect 52276 20052 52328 20058
rect 52276 19994 52328 20000
rect 52288 19854 52316 19994
rect 52368 19916 52420 19922
rect 52368 19858 52420 19864
rect 52276 19848 52328 19854
rect 52276 19790 52328 19796
rect 52380 19514 52408 19858
rect 52368 19508 52420 19514
rect 52368 19450 52420 19456
rect 52550 19272 52606 19281
rect 52550 19207 52552 19216
rect 52604 19207 52606 19216
rect 52552 19178 52604 19184
rect 52274 18864 52330 18873
rect 52656 18834 52684 20318
rect 52748 19174 52776 20420
rect 52828 20402 52880 20408
rect 52828 20324 52880 20330
rect 52828 20266 52880 20272
rect 52736 19168 52788 19174
rect 52736 19110 52788 19116
rect 52274 18799 52330 18808
rect 52644 18828 52696 18834
rect 52288 18766 52316 18799
rect 52644 18770 52696 18776
rect 52276 18760 52328 18766
rect 52276 18702 52328 18708
rect 52288 16658 52316 18702
rect 52460 18216 52512 18222
rect 52460 18158 52512 18164
rect 52368 18148 52420 18154
rect 52368 18090 52420 18096
rect 52380 16998 52408 18090
rect 52472 17746 52500 18158
rect 52460 17740 52512 17746
rect 52460 17682 52512 17688
rect 52552 17740 52604 17746
rect 52552 17682 52604 17688
rect 52368 16992 52420 16998
rect 52368 16934 52420 16940
rect 52564 16794 52592 17682
rect 52552 16788 52604 16794
rect 52552 16730 52604 16736
rect 52276 16652 52328 16658
rect 52276 16594 52328 16600
rect 52460 16448 52512 16454
rect 52460 16390 52512 16396
rect 52472 15162 52500 16390
rect 52564 16114 52592 16730
rect 52552 16108 52604 16114
rect 52552 16050 52604 16056
rect 52656 15994 52684 18770
rect 52840 18630 52868 20266
rect 52932 18834 52960 20742
rect 53116 20398 53144 20878
rect 53104 20392 53156 20398
rect 53104 20334 53156 20340
rect 53102 19952 53158 19961
rect 53012 19916 53064 19922
rect 53102 19887 53104 19896
rect 53012 19858 53064 19864
rect 53156 19887 53158 19896
rect 53104 19858 53156 19864
rect 53024 19825 53052 19858
rect 53010 19816 53066 19825
rect 53010 19751 53066 19760
rect 53104 19508 53156 19514
rect 53104 19450 53156 19456
rect 53116 19310 53144 19450
rect 53104 19304 53156 19310
rect 53104 19246 53156 19252
rect 52920 18828 52972 18834
rect 52920 18770 52972 18776
rect 52828 18624 52880 18630
rect 52828 18566 52880 18572
rect 53116 18358 53144 19246
rect 53208 18873 53236 21626
rect 53288 21344 53340 21350
rect 53288 21286 53340 21292
rect 53300 21078 53328 21286
rect 53288 21072 53340 21078
rect 53852 21026 53880 22986
rect 54116 22976 54168 22982
rect 54116 22918 54168 22924
rect 54128 22574 54156 22918
rect 54116 22568 54168 22574
rect 54116 22510 54168 22516
rect 54024 22094 54076 22098
rect 54128 22094 54156 22510
rect 54220 22438 54248 23122
rect 54404 23050 54432 23598
rect 54496 23186 54524 23598
rect 54484 23180 54536 23186
rect 54484 23122 54536 23128
rect 54680 23118 54708 24278
rect 54956 23662 54984 24636
rect 55036 24676 55088 24682
rect 55036 24618 55088 24624
rect 55048 23866 55076 24618
rect 55128 24064 55180 24070
rect 55128 24006 55180 24012
rect 55036 23860 55088 23866
rect 55036 23802 55088 23808
rect 55140 23662 55168 24006
rect 54944 23656 54996 23662
rect 54944 23598 54996 23604
rect 55128 23656 55180 23662
rect 55128 23598 55180 23604
rect 55140 23186 55168 23598
rect 55220 23588 55272 23594
rect 55220 23530 55272 23536
rect 55232 23497 55260 23530
rect 55218 23488 55274 23497
rect 55218 23423 55274 23432
rect 55128 23180 55180 23186
rect 55128 23122 55180 23128
rect 54668 23112 54720 23118
rect 54668 23054 54720 23060
rect 54392 23044 54444 23050
rect 54312 23004 54392 23032
rect 54208 22432 54260 22438
rect 54208 22374 54260 22380
rect 54220 22166 54248 22374
rect 54312 22234 54340 23004
rect 54392 22986 54444 22992
rect 54852 22568 54904 22574
rect 54852 22510 54904 22516
rect 54300 22228 54352 22234
rect 54300 22170 54352 22176
rect 54208 22160 54260 22166
rect 54208 22102 54260 22108
rect 54024 22092 54156 22094
rect 54076 22066 54156 22092
rect 54024 22034 54076 22040
rect 54312 21962 54340 22170
rect 54760 22092 54812 22098
rect 54760 22034 54812 22040
rect 54116 21956 54168 21962
rect 54116 21898 54168 21904
rect 54300 21956 54352 21962
rect 54300 21898 54352 21904
rect 54392 21956 54444 21962
rect 54392 21898 54444 21904
rect 54128 21842 54156 21898
rect 54404 21842 54432 21898
rect 54128 21814 54432 21842
rect 54484 21548 54536 21554
rect 54484 21490 54536 21496
rect 54116 21480 54168 21486
rect 54116 21422 54168 21428
rect 54024 21344 54076 21350
rect 54024 21286 54076 21292
rect 53288 21014 53340 21020
rect 53760 21010 53880 21026
rect 53748 21004 53880 21010
rect 53800 20998 53880 21004
rect 53748 20946 53800 20952
rect 53656 20936 53708 20942
rect 54036 20890 54064 21286
rect 54128 21146 54156 21422
rect 54116 21140 54168 21146
rect 54116 21082 54168 21088
rect 54298 21040 54354 21049
rect 54298 20975 54300 20984
rect 54352 20975 54354 20984
rect 54300 20946 54352 20952
rect 54116 20936 54168 20942
rect 53656 20878 53708 20884
rect 53944 20884 54116 20890
rect 53944 20878 54168 20884
rect 53668 20754 53696 20878
rect 53840 20868 53892 20874
rect 53944 20862 54156 20878
rect 54300 20868 54352 20874
rect 53944 20856 53972 20862
rect 53892 20828 53972 20856
rect 53840 20810 53892 20816
rect 54300 20810 54352 20816
rect 54024 20800 54076 20806
rect 53668 20748 54024 20754
rect 53668 20742 54076 20748
rect 53668 20726 54064 20742
rect 54312 20602 54340 20810
rect 54496 20602 54524 21490
rect 54576 21412 54628 21418
rect 54576 21354 54628 21360
rect 54588 21010 54616 21354
rect 54576 21004 54628 21010
rect 54576 20946 54628 20952
rect 54300 20596 54352 20602
rect 54300 20538 54352 20544
rect 54484 20596 54536 20602
rect 54484 20538 54536 20544
rect 53286 20496 53342 20505
rect 53286 20431 53288 20440
rect 53340 20431 53342 20440
rect 53288 20402 53340 20408
rect 54588 20398 54616 20946
rect 54300 20392 54352 20398
rect 54300 20334 54352 20340
rect 54576 20392 54628 20398
rect 54576 20334 54628 20340
rect 54312 20262 54340 20334
rect 54484 20324 54536 20330
rect 54484 20266 54536 20272
rect 54300 20256 54352 20262
rect 54300 20198 54352 20204
rect 53380 19916 53432 19922
rect 53380 19858 53432 19864
rect 53288 19372 53340 19378
rect 53288 19314 53340 19320
rect 53194 18864 53250 18873
rect 53194 18799 53250 18808
rect 53300 18630 53328 19314
rect 53392 19281 53420 19858
rect 54208 19712 54260 19718
rect 54208 19654 54260 19660
rect 54116 19304 54168 19310
rect 53378 19272 53434 19281
rect 54116 19246 54168 19252
rect 53378 19207 53434 19216
rect 53840 19236 53892 19242
rect 53840 19178 53892 19184
rect 53380 18828 53432 18834
rect 53380 18770 53432 18776
rect 53288 18624 53340 18630
rect 53288 18566 53340 18572
rect 53104 18352 53156 18358
rect 53104 18294 53156 18300
rect 53300 18222 53328 18566
rect 53012 18216 53064 18222
rect 53288 18216 53340 18222
rect 53064 18176 53144 18204
rect 53012 18158 53064 18164
rect 52920 18148 52972 18154
rect 52920 18090 52972 18096
rect 52828 18080 52880 18086
rect 52828 18022 52880 18028
rect 52736 17808 52788 17814
rect 52736 17750 52788 17756
rect 52748 16794 52776 17750
rect 52840 17746 52868 18022
rect 52932 17746 52960 18090
rect 53116 17785 53144 18176
rect 53288 18158 53340 18164
rect 53196 18148 53248 18154
rect 53196 18090 53248 18096
rect 53102 17776 53158 17785
rect 52828 17740 52880 17746
rect 52828 17682 52880 17688
rect 52920 17740 52972 17746
rect 53102 17711 53158 17720
rect 52920 17682 52972 17688
rect 52828 17604 52880 17610
rect 52828 17546 52880 17552
rect 52840 17134 52868 17546
rect 53116 17202 53144 17711
rect 53104 17196 53156 17202
rect 53104 17138 53156 17144
rect 52828 17128 52880 17134
rect 53012 17128 53064 17134
rect 52828 17070 52880 17076
rect 52932 17088 53012 17116
rect 52736 16788 52788 16794
rect 52736 16730 52788 16736
rect 52828 16652 52880 16658
rect 52828 16594 52880 16600
rect 52840 16561 52868 16594
rect 52932 16590 52960 17088
rect 53208 17082 53236 18090
rect 53392 17746 53420 18770
rect 53380 17740 53432 17746
rect 53380 17682 53432 17688
rect 53852 17678 53880 19178
rect 53932 19168 53984 19174
rect 53932 19110 53984 19116
rect 53944 18630 53972 19110
rect 54128 18834 54156 19246
rect 54220 19242 54248 19654
rect 54312 19514 54340 20198
rect 54392 19848 54444 19854
rect 54392 19790 54444 19796
rect 54300 19508 54352 19514
rect 54300 19450 54352 19456
rect 54208 19236 54260 19242
rect 54208 19178 54260 19184
rect 54312 18834 54340 19450
rect 54404 19446 54432 19790
rect 54496 19718 54524 20266
rect 54666 19952 54722 19961
rect 54772 19922 54800 22034
rect 54864 21468 54892 22510
rect 54944 22500 54996 22506
rect 54944 22442 54996 22448
rect 54956 22234 54984 22442
rect 54944 22228 54996 22234
rect 54944 22170 54996 22176
rect 54944 22092 54996 22098
rect 55128 22092 55180 22098
rect 55416 22094 55444 29124
rect 55496 27532 55548 27538
rect 55496 27474 55548 27480
rect 55680 27532 55732 27538
rect 55680 27474 55732 27480
rect 55508 26586 55536 27474
rect 55692 27130 55720 27474
rect 55680 27124 55732 27130
rect 55680 27066 55732 27072
rect 55496 26580 55548 26586
rect 55496 26522 55548 26528
rect 55494 26480 55550 26489
rect 55494 26415 55550 26424
rect 55508 26314 55536 26415
rect 55496 26308 55548 26314
rect 55496 26250 55548 26256
rect 55588 23180 55640 23186
rect 55588 23122 55640 23128
rect 55600 22778 55628 23122
rect 55588 22772 55640 22778
rect 55588 22714 55640 22720
rect 54996 22052 55128 22080
rect 54944 22034 54996 22040
rect 55128 22034 55180 22040
rect 55324 22066 55444 22094
rect 55680 22092 55732 22098
rect 55220 21888 55272 21894
rect 55218 21856 55220 21865
rect 55272 21856 55274 21865
rect 55218 21791 55274 21800
rect 55036 21480 55088 21486
rect 54864 21440 55036 21468
rect 55036 21422 55088 21428
rect 54666 19887 54722 19896
rect 54760 19916 54812 19922
rect 54574 19816 54630 19825
rect 54574 19751 54630 19760
rect 54484 19712 54536 19718
rect 54484 19654 54536 19660
rect 54392 19440 54444 19446
rect 54392 19382 54444 19388
rect 54496 19310 54524 19654
rect 54588 19378 54616 19751
rect 54576 19372 54628 19378
rect 54576 19314 54628 19320
rect 54680 19310 54708 19887
rect 54760 19858 54812 19864
rect 54772 19417 54800 19858
rect 54758 19408 54814 19417
rect 54758 19343 54814 19352
rect 54484 19304 54536 19310
rect 54484 19246 54536 19252
rect 54668 19304 54720 19310
rect 54668 19246 54720 19252
rect 54392 19236 54444 19242
rect 54392 19178 54444 19184
rect 54576 19236 54628 19242
rect 54576 19178 54628 19184
rect 54404 18834 54432 19178
rect 54116 18828 54168 18834
rect 54116 18770 54168 18776
rect 54300 18828 54352 18834
rect 54300 18770 54352 18776
rect 54392 18828 54444 18834
rect 54392 18770 54444 18776
rect 54588 18714 54616 19178
rect 54404 18686 54616 18714
rect 54404 18630 54432 18686
rect 53932 18624 53984 18630
rect 53932 18566 53984 18572
rect 54208 18624 54260 18630
rect 54208 18566 54260 18572
rect 54392 18624 54444 18630
rect 54392 18566 54444 18572
rect 54220 18222 54248 18566
rect 54680 18290 54708 19246
rect 54668 18284 54720 18290
rect 54668 18226 54720 18232
rect 54208 18216 54260 18222
rect 54208 18158 54260 18164
rect 54772 17746 54800 19343
rect 55048 19310 55076 21422
rect 55324 20482 55352 22066
rect 55680 22034 55732 22040
rect 55496 21888 55548 21894
rect 55496 21830 55548 21836
rect 55508 21418 55536 21830
rect 55496 21412 55548 21418
rect 55496 21354 55548 21360
rect 55692 21010 55720 22034
rect 55784 21298 55812 45834
rect 55864 43172 55916 43178
rect 55864 43114 55916 43120
rect 55876 42362 55904 43114
rect 55864 42356 55916 42362
rect 55864 42298 55916 42304
rect 55968 41414 55996 45970
rect 56508 45824 56560 45830
rect 56508 45766 56560 45772
rect 56048 45280 56100 45286
rect 56048 45222 56100 45228
rect 56060 44946 56088 45222
rect 56048 44940 56100 44946
rect 56048 44882 56100 44888
rect 56520 44402 56548 45766
rect 57058 45656 57114 45665
rect 57058 45591 57114 45600
rect 57072 45558 57100 45591
rect 57060 45552 57112 45558
rect 57060 45494 57112 45500
rect 57532 45490 57560 46922
rect 57612 46436 57664 46442
rect 57612 46378 57664 46384
rect 57624 46170 57652 46378
rect 57808 46170 57836 47534
rect 57980 47116 58032 47122
rect 57980 47058 58032 47064
rect 57888 46980 57940 46986
rect 57888 46922 57940 46928
rect 57900 46209 57928 46922
rect 57886 46200 57942 46209
rect 57612 46164 57664 46170
rect 57612 46106 57664 46112
rect 57796 46164 57848 46170
rect 57886 46135 57942 46144
rect 57796 46106 57848 46112
rect 57992 45558 58020 47058
rect 58268 46578 58296 55830
rect 58728 55758 58756 59200
rect 59556 57594 59584 59200
rect 59544 57588 59596 57594
rect 59544 57530 59596 57536
rect 58716 55752 58768 55758
rect 58716 55694 58768 55700
rect 58256 46572 58308 46578
rect 58256 46514 58308 46520
rect 58256 46028 58308 46034
rect 58256 45970 58308 45976
rect 57980 45552 58032 45558
rect 57980 45494 58032 45500
rect 57520 45484 57572 45490
rect 57520 45426 57572 45432
rect 57612 45416 57664 45422
rect 57612 45358 57664 45364
rect 58072 45416 58124 45422
rect 58072 45358 58124 45364
rect 57336 45348 57388 45354
rect 57336 45290 57388 45296
rect 57348 45082 57376 45290
rect 57336 45076 57388 45082
rect 57336 45018 57388 45024
rect 56692 44872 56744 44878
rect 56692 44814 56744 44820
rect 56704 44538 56732 44814
rect 56692 44532 56744 44538
rect 56692 44474 56744 44480
rect 56508 44396 56560 44402
rect 56508 44338 56560 44344
rect 56876 44260 56928 44266
rect 56876 44202 56928 44208
rect 57060 44260 57112 44266
rect 57060 44202 57112 44208
rect 56888 43994 56916 44202
rect 57072 44169 57100 44202
rect 57058 44160 57114 44169
rect 57058 44095 57114 44104
rect 56876 43988 56928 43994
rect 56876 43930 56928 43936
rect 57624 43858 57652 45358
rect 57704 45280 57756 45286
rect 57704 45222 57756 45228
rect 57716 44402 57744 45222
rect 57980 44940 58032 44946
rect 57980 44882 58032 44888
rect 57992 44538 58020 44882
rect 57980 44532 58032 44538
rect 57980 44474 58032 44480
rect 57704 44396 57756 44402
rect 57704 44338 57756 44344
rect 58084 43994 58112 45358
rect 58164 44804 58216 44810
rect 58164 44746 58216 44752
rect 58176 44577 58204 44746
rect 58162 44568 58218 44577
rect 58162 44503 58218 44512
rect 58072 43988 58124 43994
rect 58072 43930 58124 43936
rect 57612 43852 57664 43858
rect 57612 43794 57664 43800
rect 56416 43104 56468 43110
rect 56416 43046 56468 43052
rect 56428 42838 56456 43046
rect 56416 42832 56468 42838
rect 56416 42774 56468 42780
rect 57152 42764 57204 42770
rect 57152 42706 57204 42712
rect 56968 42560 57020 42566
rect 56966 42528 56968 42537
rect 57020 42528 57022 42537
rect 56966 42463 57022 42472
rect 57164 42362 57192 42706
rect 57152 42356 57204 42362
rect 57152 42298 57204 42304
rect 56140 42152 56192 42158
rect 56140 42094 56192 42100
rect 56152 41546 56180 42094
rect 57520 41608 57572 41614
rect 57520 41550 57572 41556
rect 56140 41540 56192 41546
rect 56140 41482 56192 41488
rect 56416 41540 56468 41546
rect 56416 41482 56468 41488
rect 55876 41386 55996 41414
rect 55876 39574 55904 41386
rect 56428 40730 56456 41482
rect 57060 41472 57112 41478
rect 57060 41414 57112 41420
rect 56416 40724 56468 40730
rect 56416 40666 56468 40672
rect 56600 40588 56652 40594
rect 56600 40530 56652 40536
rect 56612 39846 56640 40530
rect 57072 40526 57100 41414
rect 57532 41070 57560 41550
rect 57624 41478 57652 43794
rect 57980 43172 58032 43178
rect 57980 43114 58032 43120
rect 58164 43172 58216 43178
rect 58164 43114 58216 43120
rect 57992 42906 58020 43114
rect 58176 43081 58204 43114
rect 58162 43072 58218 43081
rect 58162 43007 58218 43016
rect 57980 42900 58032 42906
rect 57980 42842 58032 42848
rect 57704 42696 57756 42702
rect 57704 42638 57756 42644
rect 57716 41818 57744 42638
rect 57980 42084 58032 42090
rect 57980 42026 58032 42032
rect 58164 42084 58216 42090
rect 58164 42026 58216 42032
rect 57992 41818 58020 42026
rect 57704 41812 57756 41818
rect 57704 41754 57756 41760
rect 57980 41812 58032 41818
rect 57980 41754 58032 41760
rect 58176 41585 58204 42026
rect 58268 41682 58296 45970
rect 58256 41676 58308 41682
rect 58256 41618 58308 41624
rect 58162 41576 58218 41585
rect 58162 41511 58218 41520
rect 57612 41472 57664 41478
rect 57612 41414 57664 41420
rect 58268 41414 58296 41618
rect 58084 41386 58296 41414
rect 57520 41064 57572 41070
rect 57426 41032 57482 41041
rect 57244 40996 57296 41002
rect 57520 41006 57572 41012
rect 57426 40967 57428 40976
rect 57244 40938 57296 40944
rect 57480 40967 57482 40976
rect 57980 40996 58032 41002
rect 57428 40938 57480 40944
rect 57980 40938 58032 40944
rect 57060 40520 57112 40526
rect 57060 40462 57112 40468
rect 57152 40520 57204 40526
rect 57152 40462 57204 40468
rect 56600 39840 56652 39846
rect 56600 39782 56652 39788
rect 55864 39568 55916 39574
rect 55864 39510 55916 39516
rect 55876 22094 55904 39510
rect 56232 38888 56284 38894
rect 56232 38830 56284 38836
rect 56244 35562 56272 38830
rect 56612 38826 56640 39782
rect 56692 39432 56744 39438
rect 56692 39374 56744 39380
rect 56966 39400 57022 39409
rect 56600 38820 56652 38826
rect 56600 38762 56652 38768
rect 56704 38554 56732 39374
rect 56966 39335 56968 39344
rect 57020 39335 57022 39344
rect 56968 39306 57020 39312
rect 56692 38548 56744 38554
rect 56692 38490 56744 38496
rect 57072 38418 57100 40462
rect 57164 39302 57192 40462
rect 57256 40186 57284 40938
rect 57888 40928 57940 40934
rect 57888 40870 57940 40876
rect 57612 40520 57664 40526
rect 57612 40462 57664 40468
rect 57244 40180 57296 40186
rect 57244 40122 57296 40128
rect 57520 39432 57572 39438
rect 57520 39374 57572 39380
rect 57152 39296 57204 39302
rect 57152 39238 57204 39244
rect 57532 38758 57560 39374
rect 57520 38752 57572 38758
rect 57520 38694 57572 38700
rect 57624 38554 57652 40462
rect 57900 39953 57928 40870
rect 57992 40730 58020 40938
rect 57980 40724 58032 40730
rect 57980 40666 58032 40672
rect 57886 39944 57942 39953
rect 57886 39879 57942 39888
rect 57704 38820 57756 38826
rect 57704 38762 57756 38768
rect 57612 38548 57664 38554
rect 57612 38490 57664 38496
rect 57060 38412 57112 38418
rect 57060 38354 57112 38360
rect 56968 38276 57020 38282
rect 56968 38218 57020 38224
rect 56980 37942 57008 38218
rect 56968 37936 57020 37942
rect 56968 37878 57020 37884
rect 57612 37800 57664 37806
rect 57612 37742 57664 37748
rect 57060 37256 57112 37262
rect 57058 37224 57060 37233
rect 57112 37224 57114 37233
rect 57058 37159 57114 37168
rect 57624 36922 57652 37742
rect 57716 37466 57744 38762
rect 57888 38752 57940 38758
rect 57888 38694 57940 38700
rect 57900 37913 57928 38694
rect 57980 38412 58032 38418
rect 57980 38354 58032 38360
rect 57992 38010 58020 38354
rect 57980 38004 58032 38010
rect 57980 37946 58032 37952
rect 57886 37904 57942 37913
rect 57886 37839 57942 37848
rect 57704 37460 57756 37466
rect 57704 37402 57756 37408
rect 57612 36916 57664 36922
rect 57612 36858 57664 36864
rect 57428 36712 57480 36718
rect 57428 36654 57480 36660
rect 56966 36408 57022 36417
rect 56966 36343 56968 36352
rect 57020 36343 57022 36352
rect 56968 36314 57020 36320
rect 56876 36236 56928 36242
rect 56876 36178 56928 36184
rect 56968 36236 57020 36242
rect 56968 36178 57020 36184
rect 56888 35834 56916 36178
rect 56876 35828 56928 35834
rect 56876 35770 56928 35776
rect 56980 35698 57008 36178
rect 56968 35692 57020 35698
rect 56968 35634 57020 35640
rect 56232 35556 56284 35562
rect 56232 35498 56284 35504
rect 56692 35556 56744 35562
rect 56692 35498 56744 35504
rect 56324 35488 56376 35494
rect 56600 35488 56652 35494
rect 56324 35430 56376 35436
rect 56598 35456 56600 35465
rect 56652 35456 56654 35465
rect 56336 35222 56364 35430
rect 56598 35391 56654 35400
rect 56324 35216 56376 35222
rect 56324 35158 56376 35164
rect 56414 34776 56470 34785
rect 56414 34711 56470 34720
rect 56428 34678 56456 34711
rect 56416 34672 56468 34678
rect 56416 34614 56468 34620
rect 55956 34468 56008 34474
rect 55956 34410 56008 34416
rect 55968 33436 55996 34410
rect 56704 34202 56732 35498
rect 57440 35494 57468 36654
rect 57980 36644 58032 36650
rect 57980 36586 58032 36592
rect 57992 36378 58020 36586
rect 57980 36372 58032 36378
rect 57980 36314 58032 36320
rect 58084 35630 58112 41386
rect 58162 38448 58218 38457
rect 58162 38383 58164 38392
rect 58216 38383 58218 38392
rect 58164 38354 58216 38360
rect 58162 36816 58218 36825
rect 58162 36751 58164 36760
rect 58216 36751 58218 36760
rect 58164 36722 58216 36728
rect 58072 35624 58124 35630
rect 58072 35566 58124 35572
rect 58348 35624 58400 35630
rect 58348 35566 58400 35572
rect 57428 35488 57480 35494
rect 57428 35430 57480 35436
rect 57888 35488 57940 35494
rect 57888 35430 57940 35436
rect 56966 35320 57022 35329
rect 56966 35255 56968 35264
rect 57020 35255 57022 35264
rect 56968 35226 57020 35232
rect 57058 34640 57114 34649
rect 57058 34575 57060 34584
rect 57112 34575 57114 34584
rect 57060 34546 57112 34552
rect 56876 34536 56928 34542
rect 56874 34504 56876 34513
rect 56928 34504 56930 34513
rect 56874 34439 56930 34448
rect 57152 34400 57204 34406
rect 57152 34342 57204 34348
rect 56692 34196 56744 34202
rect 56692 34138 56744 34144
rect 56048 34060 56100 34066
rect 56048 34002 56100 34008
rect 56060 33658 56088 34002
rect 56048 33652 56100 33658
rect 56048 33594 56100 33600
rect 56048 33448 56100 33454
rect 55968 33408 56048 33436
rect 56048 33390 56100 33396
rect 55956 32360 56008 32366
rect 55956 32302 56008 32308
rect 55968 31278 55996 32302
rect 55956 31272 56008 31278
rect 55956 31214 56008 31220
rect 56060 30734 56088 33390
rect 56600 32768 56652 32774
rect 56600 32710 56652 32716
rect 56612 32502 56640 32710
rect 56600 32496 56652 32502
rect 56600 32438 56652 32444
rect 56704 31754 56732 34138
rect 56784 34128 56836 34134
rect 56782 34096 56784 34105
rect 56836 34096 56838 34105
rect 56782 34031 56838 34040
rect 57164 32978 57192 34342
rect 57612 33992 57664 33998
rect 57612 33934 57664 33940
rect 57520 33380 57572 33386
rect 57520 33322 57572 33328
rect 57336 33312 57388 33318
rect 57334 33280 57336 33289
rect 57388 33280 57390 33289
rect 57334 33215 57390 33224
rect 57152 32972 57204 32978
rect 57152 32914 57204 32920
rect 57336 32904 57388 32910
rect 57336 32846 57388 32852
rect 56416 31748 56468 31754
rect 56704 31726 56824 31754
rect 56416 31690 56468 31696
rect 56428 31142 56456 31690
rect 56416 31136 56468 31142
rect 56416 31078 56468 31084
rect 56048 30728 56100 30734
rect 56048 30670 56100 30676
rect 55956 29640 56008 29646
rect 55956 29582 56008 29588
rect 55968 29209 55996 29582
rect 55954 29200 56010 29209
rect 55954 29135 56010 29144
rect 56428 29102 56456 31078
rect 56508 30660 56560 30666
rect 56508 30602 56560 30608
rect 56520 29238 56548 30602
rect 56796 30122 56824 31726
rect 57348 31482 57376 32846
rect 57532 32842 57560 33322
rect 57520 32836 57572 32842
rect 57520 32778 57572 32784
rect 57428 31816 57480 31822
rect 57428 31758 57480 31764
rect 57440 31657 57468 31758
rect 57426 31648 57482 31657
rect 57426 31583 57482 31592
rect 57336 31476 57388 31482
rect 57336 31418 57388 31424
rect 57428 31272 57480 31278
rect 57428 31214 57480 31220
rect 57440 30977 57468 31214
rect 57426 30968 57482 30977
rect 57426 30903 57482 30912
rect 57244 30796 57296 30802
rect 57244 30738 57296 30744
rect 56784 30116 56836 30122
rect 56784 30058 56836 30064
rect 56876 30116 56928 30122
rect 56876 30058 56928 30064
rect 56508 29232 56560 29238
rect 56508 29174 56560 29180
rect 56232 29096 56284 29102
rect 56232 29038 56284 29044
rect 56416 29096 56468 29102
rect 56416 29038 56468 29044
rect 56244 24682 56272 29038
rect 56600 28552 56652 28558
rect 56600 28494 56652 28500
rect 56508 27872 56560 27878
rect 56508 27814 56560 27820
rect 56520 26926 56548 27814
rect 56508 26920 56560 26926
rect 56508 26862 56560 26868
rect 56324 26240 56376 26246
rect 56324 26182 56376 26188
rect 56336 25974 56364 26182
rect 56324 25968 56376 25974
rect 56324 25910 56376 25916
rect 56612 25906 56640 28494
rect 56600 25900 56652 25906
rect 56600 25842 56652 25848
rect 56690 25392 56746 25401
rect 56690 25327 56692 25336
rect 56744 25327 56746 25336
rect 56692 25298 56744 25304
rect 56232 24676 56284 24682
rect 56232 24618 56284 24624
rect 55956 24608 56008 24614
rect 55956 24550 56008 24556
rect 55968 23662 55996 24550
rect 56244 23730 56272 24618
rect 56232 23724 56284 23730
rect 56232 23666 56284 23672
rect 55956 23656 56008 23662
rect 55956 23598 56008 23604
rect 56048 23520 56100 23526
rect 56048 23462 56100 23468
rect 56060 23254 56088 23462
rect 56048 23248 56100 23254
rect 56048 23190 56100 23196
rect 56232 22772 56284 22778
rect 56232 22714 56284 22720
rect 55876 22066 55996 22094
rect 55784 21270 55904 21298
rect 55680 21004 55732 21010
rect 55680 20946 55732 20952
rect 55494 20904 55550 20913
rect 55494 20839 55550 20848
rect 55508 20806 55536 20839
rect 55496 20800 55548 20806
rect 55496 20742 55548 20748
rect 55324 20454 55444 20482
rect 55508 20466 55536 20742
rect 55692 20602 55720 20946
rect 55680 20596 55732 20602
rect 55680 20538 55732 20544
rect 55310 20360 55366 20369
rect 55310 20295 55366 20304
rect 55128 20256 55180 20262
rect 55128 20198 55180 20204
rect 55140 20074 55168 20198
rect 55140 20046 55260 20074
rect 55324 20058 55352 20295
rect 55232 19922 55260 20046
rect 55312 20052 55364 20058
rect 55312 19994 55364 20000
rect 55128 19916 55180 19922
rect 55128 19858 55180 19864
rect 55220 19916 55272 19922
rect 55220 19858 55272 19864
rect 55140 19786 55168 19858
rect 55128 19780 55180 19786
rect 55128 19722 55180 19728
rect 55220 19712 55272 19718
rect 55220 19654 55272 19660
rect 55312 19712 55364 19718
rect 55312 19654 55364 19660
rect 55232 19310 55260 19654
rect 55036 19304 55088 19310
rect 55036 19246 55088 19252
rect 55220 19304 55272 19310
rect 55220 19246 55272 19252
rect 55324 19242 55352 19654
rect 55312 19236 55364 19242
rect 55312 19178 55364 19184
rect 55220 18896 55272 18902
rect 55220 18838 55272 18844
rect 55232 18737 55260 18838
rect 55218 18728 55274 18737
rect 55218 18663 55274 18672
rect 54852 18148 54904 18154
rect 54852 18090 54904 18096
rect 54864 17882 54892 18090
rect 54852 17876 54904 17882
rect 54852 17818 54904 17824
rect 54942 17776 54998 17785
rect 53932 17740 53984 17746
rect 54760 17740 54812 17746
rect 53984 17700 54064 17728
rect 53932 17682 53984 17688
rect 53472 17672 53524 17678
rect 53472 17614 53524 17620
rect 53840 17672 53892 17678
rect 53840 17614 53892 17620
rect 53064 17076 53236 17082
rect 53012 17070 53236 17076
rect 53024 17054 53236 17070
rect 53484 17066 53512 17614
rect 53472 17060 53524 17066
rect 53472 17002 53524 17008
rect 53012 16720 53064 16726
rect 53012 16662 53064 16668
rect 53194 16688 53250 16697
rect 52920 16584 52972 16590
rect 52826 16552 52882 16561
rect 52920 16526 52972 16532
rect 52826 16487 52882 16496
rect 52564 15966 52684 15994
rect 52564 15910 52592 15966
rect 52552 15904 52604 15910
rect 52552 15846 52604 15852
rect 52644 15904 52696 15910
rect 52644 15846 52696 15852
rect 52656 15706 52684 15846
rect 52644 15700 52696 15706
rect 52644 15642 52696 15648
rect 52460 15156 52512 15162
rect 52460 15098 52512 15104
rect 52472 14958 52500 15098
rect 52460 14952 52512 14958
rect 52460 14894 52512 14900
rect 52552 14952 52604 14958
rect 52552 14894 52604 14900
rect 52736 14952 52788 14958
rect 52736 14894 52788 14900
rect 52564 14521 52592 14894
rect 52550 14512 52606 14521
rect 52368 14476 52420 14482
rect 52550 14447 52606 14456
rect 52644 14476 52696 14482
rect 52368 14418 52420 14424
rect 52644 14418 52696 14424
rect 52380 13977 52408 14418
rect 52656 14074 52684 14418
rect 52644 14068 52696 14074
rect 52644 14010 52696 14016
rect 52366 13968 52422 13977
rect 52366 13903 52422 13912
rect 52748 13870 52776 14894
rect 52552 13864 52604 13870
rect 52550 13832 52552 13841
rect 52736 13864 52788 13870
rect 52604 13832 52606 13841
rect 52736 13806 52788 13812
rect 52550 13767 52606 13776
rect 52564 13734 52592 13767
rect 52552 13728 52604 13734
rect 52840 13716 52868 16487
rect 53024 16454 53052 16662
rect 53104 16652 53156 16658
rect 53194 16623 53250 16632
rect 53104 16594 53156 16600
rect 53012 16448 53064 16454
rect 53012 16390 53064 16396
rect 53024 16114 53052 16390
rect 53012 16108 53064 16114
rect 53012 16050 53064 16056
rect 53012 15972 53064 15978
rect 53012 15914 53064 15920
rect 53024 15706 53052 15914
rect 53012 15700 53064 15706
rect 53012 15642 53064 15648
rect 53012 15564 53064 15570
rect 53116 15552 53144 16594
rect 53208 16590 53236 16623
rect 53196 16584 53248 16590
rect 53196 16526 53248 16532
rect 53288 16584 53340 16590
rect 53288 16526 53340 16532
rect 53064 15524 53144 15552
rect 53012 15506 53064 15512
rect 53208 15366 53236 16526
rect 53300 16046 53328 16526
rect 53288 16040 53340 16046
rect 53288 15982 53340 15988
rect 53300 15706 53328 15982
rect 53288 15700 53340 15706
rect 53288 15642 53340 15648
rect 53852 15638 53880 17614
rect 53930 17504 53986 17513
rect 53930 17439 53986 17448
rect 53944 17134 53972 17439
rect 54036 17377 54064 17700
rect 54942 17711 54944 17720
rect 54760 17682 54812 17688
rect 54996 17711 54998 17720
rect 54944 17682 54996 17688
rect 54758 17640 54814 17649
rect 54128 17598 54340 17626
rect 54022 17368 54078 17377
rect 54022 17303 54078 17312
rect 54128 17270 54156 17598
rect 54312 17542 54340 17598
rect 54758 17575 54814 17584
rect 54208 17536 54260 17542
rect 54208 17478 54260 17484
rect 54300 17536 54352 17542
rect 54300 17478 54352 17484
rect 54116 17264 54168 17270
rect 54116 17206 54168 17212
rect 54220 17134 54248 17478
rect 53932 17128 53984 17134
rect 53932 17070 53984 17076
rect 54208 17128 54260 17134
rect 54208 17070 54260 17076
rect 53944 16114 53972 17070
rect 54576 17060 54628 17066
rect 54576 17002 54628 17008
rect 54206 16688 54262 16697
rect 54206 16623 54208 16632
rect 54260 16623 54262 16632
rect 54484 16652 54536 16658
rect 54208 16594 54260 16600
rect 54484 16594 54536 16600
rect 53932 16108 53984 16114
rect 53932 16050 53984 16056
rect 53840 15632 53892 15638
rect 53840 15574 53892 15580
rect 53288 15564 53340 15570
rect 53288 15506 53340 15512
rect 53472 15564 53524 15570
rect 53472 15506 53524 15512
rect 53196 15360 53248 15366
rect 53196 15302 53248 15308
rect 52920 13932 52972 13938
rect 52920 13874 52972 13880
rect 52552 13670 52604 13676
rect 52748 13688 52868 13716
rect 52460 12640 52512 12646
rect 52460 12582 52512 12588
rect 52644 12640 52696 12646
rect 52644 12582 52696 12588
rect 52368 12436 52420 12442
rect 52368 12378 52420 12384
rect 52274 12336 52330 12345
rect 52274 12271 52276 12280
rect 52328 12271 52330 12280
rect 52276 12242 52328 12248
rect 52380 11286 52408 12378
rect 52472 11558 52500 12582
rect 52460 11552 52512 11558
rect 52460 11494 52512 11500
rect 52552 11552 52604 11558
rect 52552 11494 52604 11500
rect 52564 11286 52592 11494
rect 52368 11280 52420 11286
rect 52368 11222 52420 11228
rect 52552 11280 52604 11286
rect 52552 11222 52604 11228
rect 52656 11150 52684 12582
rect 52748 11354 52776 13688
rect 52932 13190 52960 13874
rect 53300 13814 53328 15506
rect 53484 15162 53512 15506
rect 54024 15360 54076 15366
rect 54024 15302 54076 15308
rect 53472 15156 53524 15162
rect 53472 15098 53524 15104
rect 54036 14958 54064 15302
rect 54024 14952 54076 14958
rect 54024 14894 54076 14900
rect 54116 14816 54168 14822
rect 54116 14758 54168 14764
rect 54024 14612 54076 14618
rect 54024 14554 54076 14560
rect 53930 14512 53986 14521
rect 53930 14447 53986 14456
rect 53944 14074 53972 14447
rect 54036 14278 54064 14554
rect 54024 14272 54076 14278
rect 54024 14214 54076 14220
rect 53932 14068 53984 14074
rect 53932 14010 53984 14016
rect 53024 13786 53328 13814
rect 52920 13184 52972 13190
rect 52920 13126 52972 13132
rect 52828 12776 52880 12782
rect 52828 12718 52880 12724
rect 52840 11898 52868 12718
rect 53024 12306 53052 13786
rect 53944 13462 53972 14010
rect 54036 13462 54064 14214
rect 54128 13802 54156 14758
rect 54220 14618 54248 16594
rect 54496 16561 54524 16594
rect 54482 16552 54538 16561
rect 54482 16487 54538 16496
rect 54484 15904 54536 15910
rect 54484 15846 54536 15852
rect 54496 15570 54524 15846
rect 54484 15564 54536 15570
rect 54404 15524 54484 15552
rect 54300 14952 54352 14958
rect 54300 14894 54352 14900
rect 54312 14618 54340 14894
rect 54208 14612 54260 14618
rect 54208 14554 54260 14560
rect 54300 14612 54352 14618
rect 54300 14554 54352 14560
rect 54404 14482 54432 15524
rect 54484 15506 54536 15512
rect 54588 15162 54616 17002
rect 54772 16794 54800 17575
rect 55220 17332 55272 17338
rect 55220 17274 55272 17280
rect 55232 17241 55260 17274
rect 55218 17232 55274 17241
rect 55218 17167 55274 17176
rect 55220 17060 55272 17066
rect 55220 17002 55272 17008
rect 54760 16788 54812 16794
rect 54760 16730 54812 16736
rect 55232 16658 55260 17002
rect 55220 16652 55272 16658
rect 55220 16594 55272 16600
rect 54852 16040 54904 16046
rect 54852 15982 54904 15988
rect 55416 15994 55444 20454
rect 55496 20460 55548 20466
rect 55496 20402 55548 20408
rect 55588 18624 55640 18630
rect 55588 18566 55640 18572
rect 55600 18222 55628 18566
rect 55588 18216 55640 18222
rect 55588 18158 55640 18164
rect 55496 17740 55548 17746
rect 55496 17682 55548 17688
rect 55508 17338 55536 17682
rect 55496 17332 55548 17338
rect 55496 17274 55548 17280
rect 55600 17270 55628 18158
rect 55678 17368 55734 17377
rect 55678 17303 55680 17312
rect 55732 17303 55734 17312
rect 55680 17274 55732 17280
rect 55588 17264 55640 17270
rect 55588 17206 55640 17212
rect 55680 16040 55732 16046
rect 54668 15360 54720 15366
rect 54668 15302 54720 15308
rect 54576 15156 54628 15162
rect 54576 15098 54628 15104
rect 54576 14612 54628 14618
rect 54576 14554 54628 14560
rect 54392 14476 54444 14482
rect 54312 14436 54392 14464
rect 54312 13954 54340 14436
rect 54392 14418 54444 14424
rect 54484 14476 54536 14482
rect 54484 14418 54536 14424
rect 54496 14346 54524 14418
rect 54484 14340 54536 14346
rect 54484 14282 54536 14288
rect 54312 13926 54432 13954
rect 54404 13870 54432 13926
rect 54300 13864 54352 13870
rect 54300 13806 54352 13812
rect 54392 13864 54444 13870
rect 54392 13806 54444 13812
rect 54116 13796 54168 13802
rect 54116 13738 54168 13744
rect 54312 13682 54340 13806
rect 54496 13682 54524 14282
rect 54588 13734 54616 14554
rect 54680 14482 54708 15302
rect 54864 15042 54892 15982
rect 55416 15966 55536 15994
rect 55680 15982 55732 15988
rect 55128 15700 55180 15706
rect 55128 15642 55180 15648
rect 54864 15014 54984 15042
rect 54956 14958 54984 15014
rect 54944 14952 54996 14958
rect 54944 14894 54996 14900
rect 54760 14884 54812 14890
rect 54760 14826 54812 14832
rect 54668 14476 54720 14482
rect 54668 14418 54720 14424
rect 54668 14272 54720 14278
rect 54668 14214 54720 14220
rect 54680 14074 54708 14214
rect 54668 14068 54720 14074
rect 54668 14010 54720 14016
rect 54772 14006 54800 14826
rect 54760 14000 54812 14006
rect 54760 13942 54812 13948
rect 54312 13654 54524 13682
rect 54576 13728 54628 13734
rect 54576 13670 54628 13676
rect 53932 13456 53984 13462
rect 53932 13398 53984 13404
rect 54024 13456 54076 13462
rect 54024 13398 54076 13404
rect 54404 13394 54432 13654
rect 54588 13394 54616 13670
rect 53196 13388 53248 13394
rect 53196 13330 53248 13336
rect 54392 13388 54444 13394
rect 54392 13330 54444 13336
rect 54576 13388 54628 13394
rect 54576 13330 54628 13336
rect 53104 13184 53156 13190
rect 53104 13126 53156 13132
rect 53116 12782 53144 13126
rect 53104 12776 53156 12782
rect 53104 12718 53156 12724
rect 53116 12646 53144 12718
rect 53104 12640 53156 12646
rect 53104 12582 53156 12588
rect 53208 12306 53236 13330
rect 54300 13320 54352 13326
rect 54300 13262 54352 13268
rect 54208 12980 54260 12986
rect 54208 12922 54260 12928
rect 54220 12782 54248 12922
rect 54312 12850 54340 13262
rect 54956 12850 54984 14894
rect 55140 14278 55168 15642
rect 55220 15564 55272 15570
rect 55220 15506 55272 15512
rect 55232 14822 55260 15506
rect 55312 14884 55364 14890
rect 55312 14826 55364 14832
rect 55220 14816 55272 14822
rect 55220 14758 55272 14764
rect 55232 14482 55260 14758
rect 55220 14476 55272 14482
rect 55220 14418 55272 14424
rect 55128 14272 55180 14278
rect 55128 14214 55180 14220
rect 55218 13832 55274 13841
rect 55218 13767 55274 13776
rect 55232 13394 55260 13767
rect 55324 13530 55352 14826
rect 55312 13524 55364 13530
rect 55312 13466 55364 13472
rect 55220 13388 55272 13394
rect 55220 13330 55272 13336
rect 55220 12980 55272 12986
rect 55220 12922 55272 12928
rect 54300 12844 54352 12850
rect 54300 12786 54352 12792
rect 54944 12844 54996 12850
rect 54944 12786 54996 12792
rect 53932 12776 53984 12782
rect 53932 12718 53984 12724
rect 54208 12776 54260 12782
rect 54208 12718 54260 12724
rect 53564 12640 53616 12646
rect 53564 12582 53616 12588
rect 53656 12640 53708 12646
rect 53656 12582 53708 12588
rect 52920 12300 52972 12306
rect 52920 12242 52972 12248
rect 53012 12300 53064 12306
rect 53196 12300 53248 12306
rect 53064 12260 53144 12288
rect 53012 12242 53064 12248
rect 52932 12102 52960 12242
rect 52920 12096 52972 12102
rect 52920 12038 52972 12044
rect 52828 11892 52880 11898
rect 52828 11834 52880 11840
rect 52840 11694 52868 11834
rect 52828 11688 52880 11694
rect 52828 11630 52880 11636
rect 53012 11552 53064 11558
rect 52840 11500 53012 11506
rect 52840 11494 53064 11500
rect 52840 11478 53052 11494
rect 52736 11348 52788 11354
rect 52736 11290 52788 11296
rect 52840 11218 52868 11478
rect 53012 11348 53064 11354
rect 53012 11290 53064 11296
rect 53024 11218 53052 11290
rect 52828 11212 52880 11218
rect 52828 11154 52880 11160
rect 53012 11212 53064 11218
rect 53012 11154 53064 11160
rect 52644 11144 52696 11150
rect 52644 11086 52696 11092
rect 52144 10560 52224 10588
rect 52092 10542 52144 10548
rect 52920 10464 52972 10470
rect 52920 10406 52972 10412
rect 52460 10124 52512 10130
rect 52380 10084 52460 10112
rect 52000 9172 52052 9178
rect 52000 9114 52052 9120
rect 51816 8492 51868 8498
rect 51816 8434 51868 8440
rect 51908 8424 51960 8430
rect 51908 8366 51960 8372
rect 51540 7880 51592 7886
rect 51540 7822 51592 7828
rect 51552 7546 51580 7822
rect 51448 7540 51500 7546
rect 51448 7482 51500 7488
rect 51540 7540 51592 7546
rect 51540 7482 51592 7488
rect 51724 7472 51776 7478
rect 51724 7414 51776 7420
rect 51632 7404 51684 7410
rect 51632 7346 51684 7352
rect 51644 6934 51672 7346
rect 51632 6928 51684 6934
rect 51632 6870 51684 6876
rect 50804 6734 50856 6740
rect 50986 6760 51042 6769
rect 50712 6248 50764 6254
rect 50712 6190 50764 6196
rect 50620 6112 50672 6118
rect 50620 6054 50672 6060
rect 50300 6012 50596 6032
rect 50356 6010 50380 6012
rect 50436 6010 50460 6012
rect 50516 6010 50540 6012
rect 50378 5958 50380 6010
rect 50442 5958 50454 6010
rect 50516 5958 50518 6010
rect 50356 5956 50380 5958
rect 50436 5956 50460 5958
rect 50516 5956 50540 5958
rect 50300 5936 50596 5956
rect 50160 5772 50212 5778
rect 50160 5714 50212 5720
rect 50724 5370 50752 6190
rect 50712 5364 50764 5370
rect 50712 5306 50764 5312
rect 50724 5166 50752 5306
rect 50160 5160 50212 5166
rect 50160 5102 50212 5108
rect 50712 5160 50764 5166
rect 50712 5102 50764 5108
rect 50172 4826 50200 5102
rect 50300 4924 50596 4944
rect 50356 4922 50380 4924
rect 50436 4922 50460 4924
rect 50516 4922 50540 4924
rect 50378 4870 50380 4922
rect 50442 4870 50454 4922
rect 50516 4870 50518 4922
rect 50356 4868 50380 4870
rect 50436 4868 50460 4870
rect 50516 4868 50540 4870
rect 50300 4848 50596 4868
rect 50160 4820 50212 4826
rect 50160 4762 50212 4768
rect 50252 4752 50304 4758
rect 50252 4694 50304 4700
rect 49884 4684 49936 4690
rect 49884 4626 49936 4632
rect 50068 4684 50120 4690
rect 50068 4626 50120 4632
rect 49792 4480 49844 4486
rect 49792 4422 49844 4428
rect 50264 4214 50292 4694
rect 50712 4616 50764 4622
rect 50710 4584 50712 4593
rect 50764 4584 50766 4593
rect 50710 4519 50766 4528
rect 50252 4208 50304 4214
rect 50066 4176 50122 4185
rect 50252 4150 50304 4156
rect 50066 4111 50122 4120
rect 50080 3942 50108 4111
rect 50068 3936 50120 3942
rect 50264 3924 50292 4150
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50356 4010 50384 4082
rect 50344 4004 50396 4010
rect 50344 3946 50396 3952
rect 50068 3878 50120 3884
rect 50172 3896 50292 3924
rect 50172 3602 50200 3896
rect 50300 3836 50596 3856
rect 50356 3834 50380 3836
rect 50436 3834 50460 3836
rect 50516 3834 50540 3836
rect 50378 3782 50380 3834
rect 50442 3782 50454 3834
rect 50516 3782 50518 3834
rect 50356 3780 50380 3782
rect 50436 3780 50460 3782
rect 50516 3780 50540 3782
rect 50300 3760 50596 3780
rect 50160 3596 50212 3602
rect 50160 3538 50212 3544
rect 50712 2916 50764 2922
rect 50712 2858 50764 2864
rect 50160 2848 50212 2854
rect 50080 2808 50160 2836
rect 49700 2508 49752 2514
rect 49700 2450 49752 2456
rect 49516 2372 49568 2378
rect 49516 2314 49568 2320
rect 49424 1896 49476 1902
rect 49424 1838 49476 1844
rect 50080 800 50108 2808
rect 50160 2790 50212 2796
rect 50300 2748 50596 2768
rect 50356 2746 50380 2748
rect 50436 2746 50460 2748
rect 50516 2746 50540 2748
rect 50378 2694 50380 2746
rect 50442 2694 50454 2746
rect 50516 2694 50518 2746
rect 50356 2692 50380 2694
rect 50436 2692 50460 2694
rect 50516 2692 50540 2694
rect 50300 2672 50596 2692
rect 50724 2650 50752 2858
rect 50712 2644 50764 2650
rect 50712 2586 50764 2592
rect 50816 2446 50844 6734
rect 50986 6695 51042 6704
rect 51540 6724 51592 6730
rect 51540 6666 51592 6672
rect 51172 6656 51224 6662
rect 51172 6598 51224 6604
rect 50896 6316 50948 6322
rect 50896 6258 50948 6264
rect 50908 6118 50936 6258
rect 50896 6112 50948 6118
rect 50896 6054 50948 6060
rect 50986 5808 51042 5817
rect 50986 5743 51042 5752
rect 51000 5710 51028 5743
rect 50896 5704 50948 5710
rect 50894 5672 50896 5681
rect 50988 5704 51040 5710
rect 50948 5672 50950 5681
rect 50988 5646 51040 5652
rect 50894 5607 50950 5616
rect 51184 5574 51212 6598
rect 51552 6322 51580 6666
rect 51540 6316 51592 6322
rect 51540 6258 51592 6264
rect 51264 6248 51316 6254
rect 51264 6190 51316 6196
rect 51172 5568 51224 5574
rect 51172 5510 51224 5516
rect 51172 5364 51224 5370
rect 51276 5352 51304 6190
rect 51736 6186 51764 7414
rect 51920 6730 51948 8366
rect 51908 6724 51960 6730
rect 51908 6666 51960 6672
rect 51816 6452 51868 6458
rect 51816 6394 51868 6400
rect 51724 6180 51776 6186
rect 51724 6122 51776 6128
rect 51356 5840 51408 5846
rect 51356 5782 51408 5788
rect 51224 5324 51304 5352
rect 51172 5306 51224 5312
rect 51184 5273 51212 5306
rect 51170 5264 51226 5273
rect 51170 5199 51226 5208
rect 50894 5128 50950 5137
rect 50894 5063 50950 5072
rect 51078 5128 51134 5137
rect 51078 5063 51134 5072
rect 50908 4622 50936 5063
rect 51092 5030 51120 5063
rect 51080 5024 51132 5030
rect 51080 4966 51132 4972
rect 51172 5024 51224 5030
rect 51172 4966 51224 4972
rect 50896 4616 50948 4622
rect 50896 4558 50948 4564
rect 50896 4480 50948 4486
rect 50894 4448 50896 4457
rect 51080 4480 51132 4486
rect 50948 4448 50950 4457
rect 50894 4383 50950 4392
rect 51078 4448 51080 4457
rect 51132 4448 51134 4457
rect 51078 4383 51134 4392
rect 50908 4078 50936 4383
rect 50896 4072 50948 4078
rect 50896 4014 50948 4020
rect 50988 3936 51040 3942
rect 51184 3924 51212 4966
rect 51040 3896 51212 3924
rect 50988 3878 51040 3884
rect 51080 2848 51132 2854
rect 51080 2790 51132 2796
rect 50804 2440 50856 2446
rect 50804 2382 50856 2388
rect 51092 800 51120 2790
rect 51368 2514 51396 5782
rect 51632 5704 51684 5710
rect 51632 5646 51684 5652
rect 51540 5568 51592 5574
rect 51540 5510 51592 5516
rect 51552 4758 51580 5510
rect 51540 4752 51592 4758
rect 51540 4694 51592 4700
rect 51448 4548 51500 4554
rect 51448 4490 51500 4496
rect 51460 3670 51488 4490
rect 51644 4060 51672 5646
rect 51724 4072 51776 4078
rect 51644 4032 51724 4060
rect 51724 4014 51776 4020
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 51540 3188 51592 3194
rect 51540 3130 51592 3136
rect 51448 2916 51500 2922
rect 51552 2904 51580 3130
rect 51632 2916 51684 2922
rect 51552 2876 51632 2904
rect 51448 2858 51500 2864
rect 51632 2858 51684 2864
rect 51460 2650 51488 2858
rect 51448 2644 51500 2650
rect 51448 2586 51500 2592
rect 51356 2508 51408 2514
rect 51356 2450 51408 2456
rect 51828 2446 51856 6394
rect 52012 5914 52040 9114
rect 52380 9042 52408 10084
rect 52460 10066 52512 10072
rect 52460 9512 52512 9518
rect 52460 9454 52512 9460
rect 52472 9382 52500 9454
rect 52460 9376 52512 9382
rect 52460 9318 52512 9324
rect 52368 9036 52420 9042
rect 52368 8978 52420 8984
rect 52092 8288 52144 8294
rect 52092 8230 52144 8236
rect 52104 8022 52132 8230
rect 52092 8016 52144 8022
rect 52092 7958 52144 7964
rect 52184 7336 52236 7342
rect 52184 7278 52236 7284
rect 52092 7200 52144 7206
rect 52092 7142 52144 7148
rect 52104 7002 52132 7142
rect 52092 6996 52144 7002
rect 52092 6938 52144 6944
rect 52104 6866 52132 6938
rect 52092 6860 52144 6866
rect 52092 6802 52144 6808
rect 52092 6248 52144 6254
rect 52092 6190 52144 6196
rect 51908 5908 51960 5914
rect 51908 5850 51960 5856
rect 52000 5908 52052 5914
rect 52000 5850 52052 5856
rect 51920 5574 51948 5850
rect 52104 5710 52132 6190
rect 52196 5778 52224 7278
rect 52380 6458 52408 8978
rect 52472 8566 52500 9318
rect 52932 9110 52960 10406
rect 53024 9110 53052 11154
rect 53116 10742 53144 12260
rect 53196 12242 53248 12248
rect 53472 12164 53524 12170
rect 53472 12106 53524 12112
rect 53484 11762 53512 12106
rect 53576 11898 53604 12582
rect 53564 11892 53616 11898
rect 53564 11834 53616 11840
rect 53472 11756 53524 11762
rect 53472 11698 53524 11704
rect 53668 11286 53696 12582
rect 53944 12345 53972 12718
rect 54312 12442 54340 12786
rect 54852 12640 54904 12646
rect 54852 12582 54904 12588
rect 54300 12436 54352 12442
rect 54300 12378 54352 12384
rect 53930 12336 53986 12345
rect 54208 12300 54260 12306
rect 53930 12271 53986 12280
rect 53944 11830 53972 12271
rect 54036 12260 54208 12288
rect 53932 11824 53984 11830
rect 53932 11766 53984 11772
rect 53656 11280 53708 11286
rect 53656 11222 53708 11228
rect 53196 11144 53248 11150
rect 53196 11086 53248 11092
rect 53104 10736 53156 10742
rect 53104 10678 53156 10684
rect 53208 10470 53236 11086
rect 54036 10810 54064 12260
rect 54208 12242 54260 12248
rect 54760 12164 54812 12170
rect 54760 12106 54812 12112
rect 54576 12096 54628 12102
rect 54576 12038 54628 12044
rect 54208 11280 54260 11286
rect 54208 11222 54260 11228
rect 54024 10804 54076 10810
rect 54024 10746 54076 10752
rect 53840 10736 53892 10742
rect 53840 10678 53892 10684
rect 53196 10464 53248 10470
rect 53196 10406 53248 10412
rect 53852 10130 53880 10678
rect 53840 10124 53892 10130
rect 53840 10066 53892 10072
rect 53932 10124 53984 10130
rect 53932 10066 53984 10072
rect 53840 9512 53892 9518
rect 53840 9454 53892 9460
rect 52920 9104 52972 9110
rect 52920 9046 52972 9052
rect 53012 9104 53064 9110
rect 53012 9046 53064 9052
rect 52828 8968 52880 8974
rect 52828 8910 52880 8916
rect 52460 8560 52512 8566
rect 52460 8502 52512 8508
rect 52840 8430 52868 8910
rect 53852 8430 53880 9454
rect 53944 9178 53972 10066
rect 54036 9518 54064 10746
rect 54220 9926 54248 11222
rect 54588 11218 54616 12038
rect 54772 11694 54800 12106
rect 54864 11694 54892 12582
rect 54956 12306 54984 12786
rect 55232 12617 55260 12922
rect 55218 12608 55274 12617
rect 55218 12543 55274 12552
rect 55128 12436 55180 12442
rect 55416 12434 55444 15966
rect 55508 15910 55536 15966
rect 55496 15904 55548 15910
rect 55496 15846 55548 15852
rect 55692 15570 55720 15982
rect 55680 15564 55732 15570
rect 55680 15506 55732 15512
rect 55588 14816 55640 14822
rect 55588 14758 55640 14764
rect 55494 14648 55550 14657
rect 55600 14618 55628 14758
rect 55494 14583 55550 14592
rect 55588 14612 55640 14618
rect 55508 14006 55536 14583
rect 55588 14554 55640 14560
rect 55600 14482 55628 14554
rect 55588 14476 55640 14482
rect 55588 14418 55640 14424
rect 55496 14000 55548 14006
rect 55496 13942 55548 13948
rect 55692 13938 55720 15506
rect 55772 15360 55824 15366
rect 55772 15302 55824 15308
rect 55784 14482 55812 15302
rect 55772 14476 55824 14482
rect 55772 14418 55824 14424
rect 55772 14272 55824 14278
rect 55772 14214 55824 14220
rect 55680 13932 55732 13938
rect 55680 13874 55732 13880
rect 55784 13870 55812 14214
rect 55772 13864 55824 13870
rect 55772 13806 55824 13812
rect 55772 13320 55824 13326
rect 55772 13262 55824 13268
rect 55588 12708 55640 12714
rect 55588 12650 55640 12656
rect 55128 12378 55180 12384
rect 55232 12406 55444 12434
rect 54944 12300 54996 12306
rect 54944 12242 54996 12248
rect 55140 11694 55168 12378
rect 54760 11688 54812 11694
rect 54760 11630 54812 11636
rect 54852 11688 54904 11694
rect 54852 11630 54904 11636
rect 55128 11688 55180 11694
rect 55128 11630 55180 11636
rect 54668 11620 54720 11626
rect 54668 11562 54720 11568
rect 54680 11286 54708 11562
rect 54668 11280 54720 11286
rect 54668 11222 54720 11228
rect 54576 11212 54628 11218
rect 54576 11154 54628 11160
rect 54680 11082 54708 11222
rect 55232 11098 55260 12406
rect 55404 12096 55456 12102
rect 55404 12038 55456 12044
rect 55416 11898 55444 12038
rect 55600 11898 55628 12650
rect 55404 11892 55456 11898
rect 55404 11834 55456 11840
rect 55588 11892 55640 11898
rect 55588 11834 55640 11840
rect 55784 11778 55812 13262
rect 55600 11750 55812 11778
rect 55600 11694 55628 11750
rect 55588 11688 55640 11694
rect 55588 11630 55640 11636
rect 55600 11286 55628 11630
rect 55588 11280 55640 11286
rect 55588 11222 55640 11228
rect 55496 11212 55548 11218
rect 55496 11154 55548 11160
rect 55680 11212 55732 11218
rect 55680 11154 55732 11160
rect 54668 11076 54720 11082
rect 55232 11070 55352 11098
rect 54668 11018 54720 11024
rect 55220 11008 55272 11014
rect 55218 10976 55220 10985
rect 55272 10976 55274 10985
rect 55218 10911 55274 10920
rect 54944 10804 54996 10810
rect 54944 10746 54996 10752
rect 54300 10736 54352 10742
rect 54300 10678 54352 10684
rect 54312 10266 54340 10678
rect 54392 10668 54444 10674
rect 54392 10610 54444 10616
rect 54760 10668 54812 10674
rect 54760 10610 54812 10616
rect 54404 10266 54432 10610
rect 54668 10532 54720 10538
rect 54668 10474 54720 10480
rect 54484 10464 54536 10470
rect 54484 10406 54536 10412
rect 54576 10464 54628 10470
rect 54576 10406 54628 10412
rect 54300 10260 54352 10266
rect 54300 10202 54352 10208
rect 54392 10260 54444 10266
rect 54392 10202 54444 10208
rect 54496 10062 54524 10406
rect 54588 10130 54616 10406
rect 54576 10124 54628 10130
rect 54576 10066 54628 10072
rect 54484 10056 54536 10062
rect 54484 9998 54536 10004
rect 54116 9920 54168 9926
rect 54116 9862 54168 9868
rect 54208 9920 54260 9926
rect 54208 9862 54260 9868
rect 54128 9518 54156 9862
rect 54024 9512 54076 9518
rect 54024 9454 54076 9460
rect 54116 9512 54168 9518
rect 54116 9454 54168 9460
rect 54220 9382 54248 9862
rect 54208 9376 54260 9382
rect 54208 9318 54260 9324
rect 54496 9178 54524 9998
rect 54680 9382 54708 10474
rect 54668 9376 54720 9382
rect 54668 9318 54720 9324
rect 53932 9172 53984 9178
rect 53932 9114 53984 9120
rect 54484 9172 54536 9178
rect 54484 9114 54536 9120
rect 53944 8498 53972 9114
rect 54392 9104 54444 9110
rect 54392 9046 54444 9052
rect 54116 8832 54168 8838
rect 54116 8774 54168 8780
rect 53932 8492 53984 8498
rect 53932 8434 53984 8440
rect 54128 8430 54156 8774
rect 52828 8424 52880 8430
rect 52828 8366 52880 8372
rect 52920 8424 52972 8430
rect 52920 8366 52972 8372
rect 53840 8424 53892 8430
rect 53840 8366 53892 8372
rect 54116 8424 54168 8430
rect 54116 8366 54168 8372
rect 52932 7954 52960 8366
rect 52920 7948 52972 7954
rect 52920 7890 52972 7896
rect 53196 7948 53248 7954
rect 53196 7890 53248 7896
rect 52828 7472 52880 7478
rect 52828 7414 52880 7420
rect 52736 6996 52788 7002
rect 52736 6938 52788 6944
rect 52748 6798 52776 6938
rect 52736 6792 52788 6798
rect 52736 6734 52788 6740
rect 52368 6452 52420 6458
rect 52368 6394 52420 6400
rect 52748 6322 52776 6734
rect 52460 6316 52512 6322
rect 52460 6258 52512 6264
rect 52736 6316 52788 6322
rect 52736 6258 52788 6264
rect 52472 6118 52500 6258
rect 52644 6248 52696 6254
rect 52644 6190 52696 6196
rect 52460 6112 52512 6118
rect 52460 6054 52512 6060
rect 52656 5914 52684 6190
rect 52644 5908 52696 5914
rect 52644 5850 52696 5856
rect 52184 5772 52236 5778
rect 52184 5714 52236 5720
rect 52092 5704 52144 5710
rect 52092 5646 52144 5652
rect 51908 5568 51960 5574
rect 51908 5510 51960 5516
rect 51920 5166 51948 5510
rect 52104 5166 52132 5646
rect 52196 5370 52224 5714
rect 52656 5574 52684 5850
rect 52840 5681 52868 7414
rect 53208 6866 53236 7890
rect 53472 7744 53524 7750
rect 53472 7686 53524 7692
rect 53564 7744 53616 7750
rect 53564 7686 53616 7692
rect 53484 7342 53512 7686
rect 53288 7336 53340 7342
rect 53288 7278 53340 7284
rect 53472 7336 53524 7342
rect 53472 7278 53524 7284
rect 53196 6860 53248 6866
rect 53196 6802 53248 6808
rect 53208 6662 53236 6802
rect 53196 6656 53248 6662
rect 53196 6598 53248 6604
rect 53300 6458 53328 7278
rect 53380 6860 53432 6866
rect 53484 6848 53512 7278
rect 53432 6820 53512 6848
rect 53380 6802 53432 6808
rect 53576 6798 53604 7686
rect 53656 7404 53708 7410
rect 53656 7346 53708 7352
rect 53564 6792 53616 6798
rect 53564 6734 53616 6740
rect 53288 6452 53340 6458
rect 53288 6394 53340 6400
rect 53196 6112 53248 6118
rect 53196 6054 53248 6060
rect 53208 5914 53236 6054
rect 53196 5908 53248 5914
rect 53196 5850 53248 5856
rect 53300 5778 53328 6394
rect 53576 6322 53604 6734
rect 53564 6316 53616 6322
rect 53564 6258 53616 6264
rect 52920 5772 52972 5778
rect 52920 5714 52972 5720
rect 53288 5772 53340 5778
rect 53288 5714 53340 5720
rect 52826 5672 52882 5681
rect 52826 5607 52882 5616
rect 52840 5574 52868 5607
rect 52644 5568 52696 5574
rect 52644 5510 52696 5516
rect 52828 5568 52880 5574
rect 52828 5510 52880 5516
rect 52184 5364 52236 5370
rect 52184 5306 52236 5312
rect 52932 5166 52960 5714
rect 53300 5370 53328 5714
rect 53288 5364 53340 5370
rect 53288 5306 53340 5312
rect 53380 5364 53432 5370
rect 53380 5306 53432 5312
rect 51908 5160 51960 5166
rect 51908 5102 51960 5108
rect 52092 5160 52144 5166
rect 52092 5102 52144 5108
rect 52920 5160 52972 5166
rect 52920 5102 52972 5108
rect 52932 4554 52960 5102
rect 53392 5030 53420 5306
rect 53380 5024 53432 5030
rect 53380 4966 53432 4972
rect 53472 5024 53524 5030
rect 53472 4966 53524 4972
rect 53380 4616 53432 4622
rect 53484 4604 53512 4966
rect 53432 4576 53512 4604
rect 53380 4558 53432 4564
rect 52920 4548 52972 4554
rect 52920 4490 52972 4496
rect 52736 4072 52788 4078
rect 52458 4040 52514 4049
rect 52458 3975 52514 3984
rect 52734 4040 52736 4049
rect 52788 4040 52790 4049
rect 52734 3975 52790 3984
rect 53104 4004 53156 4010
rect 52472 3670 52500 3975
rect 53104 3946 53156 3952
rect 52368 3664 52420 3670
rect 52368 3606 52420 3612
rect 52460 3664 52512 3670
rect 52460 3606 52512 3612
rect 52000 3392 52052 3398
rect 52000 3334 52052 3340
rect 51816 2440 51868 2446
rect 51816 2382 51868 2388
rect 51172 2372 51224 2378
rect 51172 2314 51224 2320
rect 51184 2038 51212 2314
rect 51172 2032 51224 2038
rect 51172 1974 51224 1980
rect 52012 800 52040 3334
rect 52380 2990 52408 3606
rect 52644 3596 52696 3602
rect 52644 3538 52696 3544
rect 53012 3596 53064 3602
rect 53012 3538 53064 3544
rect 52368 2984 52420 2990
rect 52368 2926 52420 2932
rect 52656 2378 52684 3538
rect 52920 3392 52972 3398
rect 52920 3334 52972 3340
rect 52644 2372 52696 2378
rect 52644 2314 52696 2320
rect 52932 800 52960 3334
rect 53024 3194 53052 3538
rect 53116 3194 53144 3946
rect 53668 3534 53696 7346
rect 53852 6798 53880 8366
rect 54404 7342 54432 9046
rect 54680 9042 54708 9318
rect 54772 9042 54800 10610
rect 54956 10606 54984 10746
rect 54944 10600 54996 10606
rect 54944 10542 54996 10548
rect 55220 10124 55272 10130
rect 55220 10066 55272 10072
rect 55232 9602 55260 10066
rect 55324 9738 55352 11070
rect 55508 10130 55536 11154
rect 55588 11144 55640 11150
rect 55588 11086 55640 11092
rect 55600 10452 55628 11086
rect 55692 10810 55720 11154
rect 55772 11144 55824 11150
rect 55772 11086 55824 11092
rect 55680 10804 55732 10810
rect 55680 10746 55732 10752
rect 55680 10464 55732 10470
rect 55600 10424 55680 10452
rect 55680 10406 55732 10412
rect 55692 10130 55720 10406
rect 55496 10124 55548 10130
rect 55496 10066 55548 10072
rect 55680 10124 55732 10130
rect 55680 10066 55732 10072
rect 55508 9994 55536 10066
rect 55496 9988 55548 9994
rect 55496 9930 55548 9936
rect 55324 9710 55444 9738
rect 55232 9574 55352 9602
rect 55218 9480 55274 9489
rect 55324 9450 55352 9574
rect 55218 9415 55220 9424
rect 55272 9415 55274 9424
rect 55312 9444 55364 9450
rect 55220 9386 55272 9392
rect 55312 9386 55364 9392
rect 54668 9036 54720 9042
rect 54668 8978 54720 8984
rect 54760 9036 54812 9042
rect 54760 8978 54812 8984
rect 54772 8430 54800 8978
rect 54944 8832 54996 8838
rect 54944 8774 54996 8780
rect 54760 8424 54812 8430
rect 54760 8366 54812 8372
rect 54956 8022 54984 8774
rect 55128 8424 55180 8430
rect 55128 8366 55180 8372
rect 54944 8016 54996 8022
rect 54944 7958 54996 7964
rect 55140 7954 55168 8366
rect 55220 8084 55272 8090
rect 55220 8026 55272 8032
rect 55232 7993 55260 8026
rect 55218 7984 55274 7993
rect 54760 7948 54812 7954
rect 54760 7890 54812 7896
rect 55128 7948 55180 7954
rect 55218 7919 55274 7928
rect 55128 7890 55180 7896
rect 54772 7750 54800 7890
rect 54760 7744 54812 7750
rect 55416 7721 55444 9710
rect 55692 9674 55720 10066
rect 55784 10062 55812 11086
rect 55772 10056 55824 10062
rect 55772 9998 55824 10004
rect 55600 9646 55720 9674
rect 55600 9518 55628 9646
rect 55588 9512 55640 9518
rect 55588 9454 55640 9460
rect 55876 7750 55904 21270
rect 55968 15706 55996 22066
rect 56244 22030 56272 22714
rect 56232 22024 56284 22030
rect 56232 21966 56284 21972
rect 56508 21888 56560 21894
rect 56508 21830 56560 21836
rect 56048 21344 56100 21350
rect 56520 21321 56548 21830
rect 56600 21480 56652 21486
rect 56600 21422 56652 21428
rect 56048 21286 56100 21292
rect 56506 21312 56562 21321
rect 56060 20942 56088 21286
rect 56506 21247 56562 21256
rect 56048 20936 56100 20942
rect 56048 20878 56100 20884
rect 56060 20398 56088 20878
rect 56612 20874 56640 21422
rect 56600 20868 56652 20874
rect 56600 20810 56652 20816
rect 56048 20392 56100 20398
rect 56048 20334 56100 20340
rect 56692 18896 56744 18902
rect 56692 18838 56744 18844
rect 56140 18828 56192 18834
rect 56140 18770 56192 18776
rect 56152 18426 56180 18770
rect 56140 18420 56192 18426
rect 56140 18362 56192 18368
rect 56152 18034 56180 18362
rect 56152 18006 56272 18034
rect 56244 17134 56272 18006
rect 56508 17672 56560 17678
rect 56508 17614 56560 17620
rect 56520 17134 56548 17614
rect 56232 17128 56284 17134
rect 56232 17070 56284 17076
rect 56508 17128 56560 17134
rect 56508 17070 56560 17076
rect 56600 16652 56652 16658
rect 56600 16594 56652 16600
rect 55956 15700 56008 15706
rect 55956 15642 56008 15648
rect 56324 15700 56376 15706
rect 56324 15642 56376 15648
rect 55956 14476 56008 14482
rect 55956 14418 56008 14424
rect 55968 13394 55996 14418
rect 56046 14240 56102 14249
rect 56046 14175 56102 14184
rect 56060 13870 56088 14175
rect 56048 13864 56100 13870
rect 56048 13806 56100 13812
rect 56140 13728 56192 13734
rect 56138 13696 56140 13705
rect 56192 13696 56194 13705
rect 56138 13631 56194 13640
rect 55956 13388 56008 13394
rect 55956 13330 56008 13336
rect 56336 11694 56364 15642
rect 56612 15570 56640 16594
rect 56704 16454 56732 18838
rect 56796 18834 56824 30058
rect 56888 29306 56916 30058
rect 57256 29578 57284 30738
rect 57428 30660 57480 30666
rect 57428 30602 57480 30608
rect 57440 30161 57468 30602
rect 57520 30592 57572 30598
rect 57520 30534 57572 30540
rect 57532 30258 57560 30534
rect 57520 30252 57572 30258
rect 57520 30194 57572 30200
rect 57426 30152 57482 30161
rect 57426 30087 57482 30096
rect 57520 30048 57572 30054
rect 57520 29990 57572 29996
rect 57244 29572 57296 29578
rect 57244 29514 57296 29520
rect 56876 29300 56928 29306
rect 56876 29242 56928 29248
rect 57058 28656 57114 28665
rect 56876 28620 56928 28626
rect 57532 28626 57560 29990
rect 57624 29306 57652 33934
rect 57900 29714 57928 35430
rect 58256 35080 58308 35086
rect 58256 35022 58308 35028
rect 57980 34536 58032 34542
rect 57980 34478 58032 34484
rect 57992 33998 58020 34478
rect 57980 33992 58032 33998
rect 57980 33934 58032 33940
rect 57980 33856 58032 33862
rect 57980 33798 58032 33804
rect 58162 33824 58218 33833
rect 57992 33454 58020 33798
rect 58162 33759 58218 33768
rect 58176 33590 58204 33759
rect 58164 33584 58216 33590
rect 58164 33526 58216 33532
rect 57980 33448 58032 33454
rect 57980 33390 58032 33396
rect 57980 32224 58032 32230
rect 57980 32166 58032 32172
rect 58162 32192 58218 32201
rect 57992 31958 58020 32166
rect 58162 32127 58218 32136
rect 58176 31958 58204 32127
rect 57980 31952 58032 31958
rect 57980 31894 58032 31900
rect 58164 31952 58216 31958
rect 58164 31894 58216 31900
rect 58072 31884 58124 31890
rect 58072 31826 58124 31832
rect 58084 31482 58112 31826
rect 58072 31476 58124 31482
rect 58072 31418 58124 31424
rect 57980 30796 58032 30802
rect 57980 30738 58032 30744
rect 57992 30394 58020 30738
rect 58162 30696 58218 30705
rect 58162 30631 58164 30640
rect 58216 30631 58218 30640
rect 58164 30602 58216 30608
rect 57980 30388 58032 30394
rect 57980 30330 58032 30336
rect 58268 29850 58296 35022
rect 58256 29844 58308 29850
rect 58256 29786 58308 29792
rect 57888 29708 57940 29714
rect 57888 29650 57940 29656
rect 57612 29300 57664 29306
rect 57612 29242 57664 29248
rect 57900 29102 57928 29650
rect 57888 29096 57940 29102
rect 57888 29038 57940 29044
rect 58162 29064 58218 29073
rect 57980 29028 58032 29034
rect 58162 28999 58164 29008
rect 57980 28970 58032 28976
rect 58216 28999 58218 29008
rect 58164 28970 58216 28976
rect 57992 28762 58020 28970
rect 57980 28756 58032 28762
rect 57980 28698 58032 28704
rect 57058 28591 57060 28600
rect 56876 28562 56928 28568
rect 57112 28591 57114 28600
rect 57520 28620 57572 28626
rect 57060 28562 57112 28568
rect 57520 28562 57572 28568
rect 56888 28218 56916 28562
rect 56876 28212 56928 28218
rect 56876 28154 56928 28160
rect 57244 28008 57296 28014
rect 57244 27950 57296 27956
rect 57060 27600 57112 27606
rect 57058 27568 57060 27577
rect 57112 27568 57114 27577
rect 57058 27503 57114 27512
rect 57256 27062 57284 27950
rect 57704 27464 57756 27470
rect 57704 27406 57756 27412
rect 57244 27056 57296 27062
rect 57244 26998 57296 27004
rect 57334 27024 57390 27033
rect 57334 26959 57390 26968
rect 57152 26920 57204 26926
rect 57152 26862 57204 26868
rect 57164 26042 57192 26862
rect 57244 26784 57296 26790
rect 57244 26726 57296 26732
rect 57256 26518 57284 26726
rect 57348 26586 57376 26959
rect 57336 26580 57388 26586
rect 57336 26522 57388 26528
rect 57244 26512 57296 26518
rect 57244 26454 57296 26460
rect 57152 26036 57204 26042
rect 57152 25978 57204 25984
rect 57716 25945 57744 27406
rect 57980 26444 58032 26450
rect 57980 26386 58032 26392
rect 57888 26308 57940 26314
rect 57888 26250 57940 26256
rect 57900 26081 57928 26250
rect 57886 26072 57942 26081
rect 57992 26042 58020 26386
rect 57886 26007 57942 26016
rect 57980 26036 58032 26042
rect 57980 25978 58032 25984
rect 57702 25936 57758 25945
rect 57702 25871 57758 25880
rect 57704 25832 57756 25838
rect 57704 25774 57756 25780
rect 57716 25158 57744 25774
rect 58162 25528 58218 25537
rect 58162 25463 58218 25472
rect 58176 25430 58204 25463
rect 58164 25424 58216 25430
rect 58164 25366 58216 25372
rect 57704 25152 57756 25158
rect 57704 25094 57756 25100
rect 58360 24750 58388 35566
rect 57336 24744 57388 24750
rect 57336 24686 57388 24692
rect 58348 24744 58400 24750
rect 58348 24686 58400 24692
rect 56876 24268 56928 24274
rect 56876 24210 56928 24216
rect 56888 23050 56916 24210
rect 56968 24064 57020 24070
rect 56968 24006 57020 24012
rect 56980 23905 57008 24006
rect 56966 23896 57022 23905
rect 56966 23831 57022 23840
rect 57244 23588 57296 23594
rect 57244 23530 57296 23536
rect 57150 23216 57206 23225
rect 57150 23151 57152 23160
rect 57204 23151 57206 23160
rect 57152 23122 57204 23128
rect 56876 23044 56928 23050
rect 56876 22986 56928 22992
rect 57256 22778 57284 23530
rect 57244 22772 57296 22778
rect 57244 22714 57296 22720
rect 57244 20936 57296 20942
rect 57244 20878 57296 20884
rect 57256 20534 57284 20878
rect 57244 20528 57296 20534
rect 57244 20470 57296 20476
rect 56876 19916 56928 19922
rect 56876 19858 56928 19864
rect 56888 19514 56916 19858
rect 57060 19780 57112 19786
rect 57060 19722 57112 19728
rect 56876 19508 56928 19514
rect 56876 19450 56928 19456
rect 56968 19304 57020 19310
rect 57072 19281 57100 19722
rect 57152 19304 57204 19310
rect 56968 19246 57020 19252
rect 57058 19272 57114 19281
rect 56980 19009 57008 19246
rect 57152 19246 57204 19252
rect 57058 19207 57114 19216
rect 56966 19000 57022 19009
rect 57164 18970 57192 19246
rect 56966 18935 57022 18944
rect 57152 18964 57204 18970
rect 57152 18906 57204 18912
rect 57348 18902 57376 24686
rect 57980 24676 58032 24682
rect 57980 24618 58032 24624
rect 58164 24676 58216 24682
rect 58164 24618 58216 24624
rect 57992 24410 58020 24618
rect 58176 24449 58204 24618
rect 58162 24440 58218 24449
rect 57980 24404 58032 24410
rect 58162 24375 58218 24384
rect 57980 24346 58032 24352
rect 57704 24200 57756 24206
rect 57704 24142 57756 24148
rect 57716 23798 57744 24142
rect 57704 23792 57756 23798
rect 57704 23734 57756 23740
rect 57428 23588 57480 23594
rect 57428 23530 57480 23536
rect 57980 23588 58032 23594
rect 57980 23530 58032 23536
rect 57440 22409 57468 23530
rect 57888 23520 57940 23526
rect 57888 23462 57940 23468
rect 57900 22953 57928 23462
rect 57886 22944 57942 22953
rect 57886 22879 57942 22888
rect 57426 22400 57482 22409
rect 57426 22335 57482 22344
rect 57704 22024 57756 22030
rect 57704 21966 57756 21972
rect 57716 21690 57744 21966
rect 57992 21962 58020 23530
rect 58072 22160 58124 22166
rect 58072 22102 58124 22108
rect 57980 21956 58032 21962
rect 57980 21898 58032 21904
rect 58084 21690 58112 22102
rect 57704 21684 57756 21690
rect 57704 21626 57756 21632
rect 58072 21684 58124 21690
rect 58072 21626 58124 21632
rect 57518 20904 57574 20913
rect 57518 20839 57574 20848
rect 57428 20800 57480 20806
rect 57428 20742 57480 20748
rect 57440 20398 57468 20742
rect 57532 20534 57560 20839
rect 57520 20528 57572 20534
rect 57520 20470 57572 20476
rect 57428 20392 57480 20398
rect 57428 20334 57480 20340
rect 57980 20324 58032 20330
rect 57980 20266 58032 20272
rect 58164 20324 58216 20330
rect 58164 20266 58216 20272
rect 57992 20058 58020 20266
rect 57980 20052 58032 20058
rect 57980 19994 58032 20000
rect 58176 19825 58204 20266
rect 58162 19816 58218 19825
rect 58162 19751 58218 19760
rect 57336 18896 57388 18902
rect 57336 18838 57388 18844
rect 56784 18828 56836 18834
rect 56784 18770 56836 18776
rect 57980 18828 58032 18834
rect 57980 18770 58032 18776
rect 56796 18465 56824 18770
rect 56782 18456 56838 18465
rect 57992 18426 58020 18770
rect 58164 18692 58216 18698
rect 58164 18634 58216 18640
rect 56782 18391 56838 18400
rect 57980 18420 58032 18426
rect 57980 18362 58032 18368
rect 58176 18329 58204 18634
rect 58162 18320 58218 18329
rect 58162 18255 58218 18264
rect 57520 18216 57572 18222
rect 57520 18158 57572 18164
rect 56876 18148 56928 18154
rect 56876 18090 56928 18096
rect 57060 18148 57112 18154
rect 57060 18090 57112 18096
rect 56888 17610 56916 18090
rect 57072 17785 57100 18090
rect 57058 17776 57114 17785
rect 57058 17711 57114 17720
rect 56968 17672 57020 17678
rect 56968 17614 57020 17620
rect 57152 17672 57204 17678
rect 57152 17614 57204 17620
rect 56876 17604 56928 17610
rect 56876 17546 56928 17552
rect 56980 16998 57008 17614
rect 57164 17105 57192 17614
rect 57532 17542 57560 18158
rect 57520 17536 57572 17542
rect 57520 17478 57572 17484
rect 57150 17096 57206 17105
rect 57150 17031 57206 17040
rect 57244 17060 57296 17066
rect 57244 17002 57296 17008
rect 57428 17060 57480 17066
rect 57428 17002 57480 17008
rect 57980 17060 58032 17066
rect 57980 17002 58032 17008
rect 58164 17060 58216 17066
rect 58164 17002 58216 17008
rect 56968 16992 57020 16998
rect 56968 16934 57020 16940
rect 56692 16448 56744 16454
rect 56692 16390 56744 16396
rect 57256 16250 57284 17002
rect 57244 16244 57296 16250
rect 57244 16186 57296 16192
rect 57440 16153 57468 17002
rect 57992 16794 58020 17002
rect 57980 16788 58032 16794
rect 57980 16730 58032 16736
rect 58176 16697 58204 17002
rect 58162 16688 58218 16697
rect 58162 16623 58218 16632
rect 57426 16144 57482 16153
rect 57426 16079 57482 16088
rect 56600 15564 56652 15570
rect 56600 15506 56652 15512
rect 57980 15564 58032 15570
rect 57980 15506 58032 15512
rect 57888 15360 57940 15366
rect 57888 15302 57940 15308
rect 57900 15201 57928 15302
rect 57886 15192 57942 15201
rect 57992 15162 58020 15506
rect 57886 15127 57942 15136
rect 57980 15156 58032 15162
rect 57980 15098 58032 15104
rect 57060 13864 57112 13870
rect 57060 13806 57112 13812
rect 57520 13864 57572 13870
rect 57520 13806 57572 13812
rect 57704 13864 57756 13870
rect 57704 13806 57756 13812
rect 57072 13569 57100 13806
rect 57058 13560 57114 13569
rect 57058 13495 57114 13504
rect 57244 13184 57296 13190
rect 57244 13126 57296 13132
rect 57334 13152 57390 13161
rect 57256 12782 57284 13126
rect 57334 13087 57390 13096
rect 57348 12986 57376 13087
rect 57336 12980 57388 12986
rect 57336 12922 57388 12928
rect 57532 12850 57560 13806
rect 57520 12844 57572 12850
rect 57520 12786 57572 12792
rect 57244 12776 57296 12782
rect 57244 12718 57296 12724
rect 56692 12640 56744 12646
rect 56692 12582 56744 12588
rect 56704 12306 56732 12582
rect 56692 12300 56744 12306
rect 56692 12242 56744 12248
rect 57612 12232 57664 12238
rect 57612 12174 57664 12180
rect 56692 11824 56744 11830
rect 56692 11766 56744 11772
rect 56324 11688 56376 11694
rect 56324 11630 56376 11636
rect 56704 11354 56732 11766
rect 57152 11688 57204 11694
rect 57150 11656 57152 11665
rect 57204 11656 57206 11665
rect 57150 11591 57206 11600
rect 56692 11348 56744 11354
rect 56692 11290 56744 11296
rect 56704 11098 56732 11290
rect 56704 11070 56824 11098
rect 56692 11008 56744 11014
rect 56692 10950 56744 10956
rect 56704 10606 56732 10950
rect 56692 10600 56744 10606
rect 56692 10542 56744 10548
rect 55956 9376 56008 9382
rect 55956 9318 56008 9324
rect 55968 8362 55996 9318
rect 56796 9042 56824 11070
rect 57520 10532 57572 10538
rect 57520 10474 57572 10480
rect 56876 10124 56928 10130
rect 56876 10066 56928 10072
rect 56888 9722 56916 10066
rect 57058 10024 57114 10033
rect 57058 9959 57060 9968
rect 57112 9959 57114 9968
rect 57060 9930 57112 9936
rect 56876 9716 56928 9722
rect 56876 9658 56928 9664
rect 56968 9512 57020 9518
rect 56968 9454 57020 9460
rect 56784 9036 56836 9042
rect 56784 8978 56836 8984
rect 56600 8424 56652 8430
rect 56600 8366 56652 8372
rect 55956 8356 56008 8362
rect 55956 8298 56008 8304
rect 56612 8129 56640 8366
rect 56598 8120 56654 8129
rect 56598 8055 56654 8064
rect 56796 7954 56824 8978
rect 56980 8906 57008 9454
rect 57532 9042 57560 10474
rect 57520 9036 57572 9042
rect 57520 8978 57572 8984
rect 56968 8900 57020 8906
rect 56968 8842 57020 8848
rect 57428 8288 57480 8294
rect 57428 8230 57480 8236
rect 56784 7948 56836 7954
rect 56784 7890 56836 7896
rect 55496 7744 55548 7750
rect 54760 7686 54812 7692
rect 55402 7712 55458 7721
rect 55496 7686 55548 7692
rect 55864 7744 55916 7750
rect 55864 7686 55916 7692
rect 55402 7647 55458 7656
rect 54576 7404 54628 7410
rect 54576 7346 54628 7352
rect 54392 7336 54444 7342
rect 54128 7296 54392 7324
rect 53840 6792 53892 6798
rect 53840 6734 53892 6740
rect 53748 6112 53800 6118
rect 53748 6054 53800 6060
rect 53760 5778 53788 6054
rect 53748 5772 53800 5778
rect 53748 5714 53800 5720
rect 53852 5030 53880 6734
rect 54024 6248 54076 6254
rect 54024 6190 54076 6196
rect 54036 5778 54064 6190
rect 54024 5772 54076 5778
rect 54024 5714 54076 5720
rect 54024 5160 54076 5166
rect 54128 5148 54156 7296
rect 54392 7278 54444 7284
rect 54208 6452 54260 6458
rect 54208 6394 54260 6400
rect 54220 6254 54248 6394
rect 54588 6254 54616 7346
rect 54760 7200 54812 7206
rect 54760 7142 54812 7148
rect 54772 6934 54800 7142
rect 54760 6928 54812 6934
rect 54760 6870 54812 6876
rect 55312 6860 55364 6866
rect 55312 6802 55364 6808
rect 55220 6656 55272 6662
rect 55220 6598 55272 6604
rect 55232 6254 55260 6598
rect 55324 6361 55352 6802
rect 55310 6352 55366 6361
rect 55310 6287 55366 6296
rect 54208 6248 54260 6254
rect 54208 6190 54260 6196
rect 54300 6248 54352 6254
rect 54300 6190 54352 6196
rect 54576 6248 54628 6254
rect 54576 6190 54628 6196
rect 55220 6248 55272 6254
rect 55220 6190 55272 6196
rect 54220 5166 54248 6190
rect 54312 5574 54340 6190
rect 55508 6066 55536 7686
rect 56796 7410 56824 7890
rect 56968 7880 57020 7886
rect 57336 7880 57388 7886
rect 56968 7822 57020 7828
rect 57334 7848 57336 7857
rect 57388 7848 57390 7857
rect 56876 7744 56928 7750
rect 56876 7686 56928 7692
rect 56784 7404 56836 7410
rect 56784 7346 56836 7352
rect 56508 6248 56560 6254
rect 56508 6190 56560 6196
rect 55232 6038 55536 6066
rect 54760 5772 54812 5778
rect 54760 5714 54812 5720
rect 54300 5568 54352 5574
rect 54300 5510 54352 5516
rect 54076 5120 54156 5148
rect 54208 5160 54260 5166
rect 54024 5102 54076 5108
rect 54392 5160 54444 5166
rect 54208 5102 54260 5108
rect 54390 5128 54392 5137
rect 54444 5128 54446 5137
rect 54390 5063 54446 5072
rect 53840 5024 53892 5030
rect 53840 4966 53892 4972
rect 54116 5024 54168 5030
rect 54116 4966 54168 4972
rect 54128 4758 54156 4966
rect 54116 4752 54168 4758
rect 54116 4694 54168 4700
rect 54772 4486 54800 5714
rect 55232 4978 55260 6038
rect 55404 5908 55456 5914
rect 55404 5850 55456 5856
rect 55312 5228 55364 5234
rect 55312 5170 55364 5176
rect 55140 4950 55260 4978
rect 55140 4706 55168 4950
rect 55218 4856 55274 4865
rect 55218 4791 55220 4800
rect 55272 4791 55274 4800
rect 55220 4762 55272 4768
rect 55140 4678 55260 4706
rect 54760 4480 54812 4486
rect 54760 4422 54812 4428
rect 55232 4049 55260 4678
rect 55218 4040 55274 4049
rect 55036 4004 55088 4010
rect 55218 3975 55274 3984
rect 55036 3946 55088 3952
rect 54208 3936 54260 3942
rect 54206 3904 54208 3913
rect 54484 3936 54536 3942
rect 54260 3904 54262 3913
rect 54484 3878 54536 3884
rect 54206 3839 54262 3848
rect 53656 3528 53708 3534
rect 53656 3470 53708 3476
rect 54392 3392 54444 3398
rect 54392 3334 54444 3340
rect 53012 3188 53064 3194
rect 53012 3130 53064 3136
rect 53104 3188 53156 3194
rect 53104 3130 53156 3136
rect 54404 2990 54432 3334
rect 54392 2984 54444 2990
rect 54392 2926 54444 2932
rect 54116 2916 54168 2922
rect 54116 2858 54168 2864
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 53852 800 53880 2790
rect 54128 2650 54156 2858
rect 54116 2644 54168 2650
rect 54116 2586 54168 2592
rect 54496 1698 54524 3878
rect 55048 3194 55076 3946
rect 55232 3602 55260 3975
rect 55220 3596 55272 3602
rect 55220 3538 55272 3544
rect 55220 3460 55272 3466
rect 55220 3402 55272 3408
rect 55232 3233 55260 3402
rect 55324 3398 55352 5170
rect 55312 3392 55364 3398
rect 55312 3334 55364 3340
rect 55218 3224 55274 3233
rect 54852 3188 54904 3194
rect 54852 3130 54904 3136
rect 55036 3188 55088 3194
rect 55218 3159 55274 3168
rect 55036 3130 55088 3136
rect 54864 2961 54892 3130
rect 54850 2952 54906 2961
rect 54850 2887 54906 2896
rect 54760 2848 54812 2854
rect 54760 2790 54812 2796
rect 54668 2304 54720 2310
rect 54668 2246 54720 2252
rect 54680 2106 54708 2246
rect 54668 2100 54720 2106
rect 54668 2042 54720 2048
rect 54484 1692 54536 1698
rect 54484 1634 54536 1640
rect 54772 800 54800 2790
rect 55416 2774 55444 5850
rect 56324 5772 56376 5778
rect 56324 5714 56376 5720
rect 55496 5364 55548 5370
rect 55496 5306 55548 5312
rect 55508 5166 55536 5306
rect 55772 5296 55824 5302
rect 55772 5238 55824 5244
rect 55496 5160 55548 5166
rect 55496 5102 55548 5108
rect 55588 4548 55640 4554
rect 55588 4490 55640 4496
rect 55600 4282 55628 4490
rect 55588 4276 55640 4282
rect 55588 4218 55640 4224
rect 55588 4004 55640 4010
rect 55588 3946 55640 3952
rect 55494 3360 55550 3369
rect 55494 3295 55550 3304
rect 55508 3058 55536 3295
rect 55496 3052 55548 3058
rect 55496 2994 55548 3000
rect 55324 2746 55444 2774
rect 55220 2576 55272 2582
rect 55220 2518 55272 2524
rect 55128 2440 55180 2446
rect 55128 2382 55180 2388
rect 55140 1970 55168 2382
rect 55128 1964 55180 1970
rect 55128 1906 55180 1912
rect 55232 1737 55260 2518
rect 55324 2514 55352 2746
rect 55600 2650 55628 3946
rect 55680 3936 55732 3942
rect 55680 3878 55732 3884
rect 55588 2644 55640 2650
rect 55588 2586 55640 2592
rect 55312 2508 55364 2514
rect 55312 2450 55364 2456
rect 55218 1728 55274 1737
rect 55218 1663 55274 1672
rect 55220 1352 55272 1358
rect 55220 1294 55272 1300
rect 2962 504 3018 513
rect 2962 439 3018 448
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9770 0 9826 800
rect 10782 0 10838 800
rect 11702 0 11758 800
rect 12622 0 12678 800
rect 13542 0 13598 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17314 0 17370 800
rect 18234 0 18290 800
rect 19154 0 19210 800
rect 20074 0 20130 800
rect 21086 0 21142 800
rect 22006 0 22062 800
rect 22926 0 22982 800
rect 23846 0 23902 800
rect 24766 0 24822 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32310 0 32366 800
rect 33230 0 33286 800
rect 34150 0 34206 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38842 0 38898 800
rect 39762 0 39818 800
rect 40774 0 40830 800
rect 41694 0 41750 800
rect 42614 0 42670 800
rect 43534 0 43590 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46386 0 46442 800
rect 47306 0 47362 800
rect 48226 0 48282 800
rect 49146 0 49202 800
rect 50066 0 50122 800
rect 51078 0 51134 800
rect 51998 0 52054 800
rect 52918 0 52974 800
rect 53838 0 53894 800
rect 54758 0 54814 800
rect 55232 241 55260 1294
rect 55692 898 55720 3878
rect 55784 3670 55812 5238
rect 56232 5024 56284 5030
rect 56232 4966 56284 4972
rect 55954 4040 56010 4049
rect 55954 3975 56010 3984
rect 56048 4004 56100 4010
rect 55772 3664 55824 3670
rect 55772 3606 55824 3612
rect 55772 3460 55824 3466
rect 55772 3402 55824 3408
rect 55784 2281 55812 3402
rect 55968 2990 55996 3975
rect 56048 3946 56100 3952
rect 56060 3777 56088 3946
rect 56046 3768 56102 3777
rect 56046 3703 56102 3712
rect 56244 3194 56272 4966
rect 56232 3188 56284 3194
rect 56232 3130 56284 3136
rect 55956 2984 56008 2990
rect 55862 2952 55918 2961
rect 55956 2926 56008 2932
rect 55862 2887 55864 2896
rect 55916 2887 55918 2896
rect 55864 2858 55916 2864
rect 56336 2650 56364 5714
rect 56520 5642 56548 6190
rect 56692 5704 56744 5710
rect 56692 5646 56744 5652
rect 56784 5704 56836 5710
rect 56784 5646 56836 5652
rect 56508 5636 56560 5642
rect 56508 5578 56560 5584
rect 56416 5568 56468 5574
rect 56416 5510 56468 5516
rect 56600 5568 56652 5574
rect 56704 5545 56732 5646
rect 56600 5510 56652 5516
rect 56690 5536 56746 5545
rect 56428 3602 56456 5510
rect 56508 5092 56560 5098
rect 56508 5034 56560 5040
rect 56520 4282 56548 5034
rect 56508 4276 56560 4282
rect 56508 4218 56560 4224
rect 56612 4010 56640 5510
rect 56690 5471 56746 5480
rect 56690 4176 56746 4185
rect 56690 4111 56692 4120
rect 56744 4111 56746 4120
rect 56692 4082 56744 4088
rect 56600 4004 56652 4010
rect 56600 3946 56652 3952
rect 56796 3913 56824 5646
rect 56782 3904 56838 3913
rect 56782 3839 56838 3848
rect 56888 3670 56916 7686
rect 56980 6866 57008 7822
rect 57334 7783 57390 7792
rect 57060 7200 57112 7206
rect 57060 7142 57112 7148
rect 57072 6934 57100 7142
rect 57060 6928 57112 6934
rect 57060 6870 57112 6876
rect 57150 6896 57206 6905
rect 56968 6860 57020 6866
rect 57150 6831 57206 6840
rect 56968 6802 57020 6808
rect 57164 6798 57192 6831
rect 57440 6798 57468 8230
rect 57624 8090 57652 12174
rect 57716 9178 57744 13806
rect 57980 12708 58032 12714
rect 57980 12650 58032 12656
rect 57888 12640 57940 12646
rect 57888 12582 57940 12588
rect 57900 12073 57928 12582
rect 57992 12442 58020 12650
rect 57980 12436 58032 12442
rect 57980 12378 58032 12384
rect 57886 12064 57942 12073
rect 57886 11999 57942 12008
rect 57980 11552 58032 11558
rect 57980 11494 58032 11500
rect 58162 11520 58218 11529
rect 57992 11286 58020 11494
rect 58162 11455 58218 11464
rect 58176 11286 58204 11455
rect 57980 11280 58032 11286
rect 57980 11222 58032 11228
rect 58164 11280 58216 11286
rect 58164 11222 58216 11228
rect 58162 10568 58218 10577
rect 57980 10532 58032 10538
rect 58162 10503 58164 10512
rect 57980 10474 58032 10480
rect 58216 10503 58218 10512
rect 58164 10474 58216 10480
rect 57992 10266 58020 10474
rect 57980 10260 58032 10266
rect 57980 10202 58032 10208
rect 57980 9444 58032 9450
rect 57980 9386 58032 9392
rect 58164 9444 58216 9450
rect 58164 9386 58216 9392
rect 57992 9178 58020 9386
rect 57704 9172 57756 9178
rect 57704 9114 57756 9120
rect 57980 9172 58032 9178
rect 57980 9114 58032 9120
rect 57704 8968 57756 8974
rect 58176 8945 58204 9386
rect 57704 8910 57756 8916
rect 58162 8936 58218 8945
rect 57612 8084 57664 8090
rect 57612 8026 57664 8032
rect 57716 7546 57744 8910
rect 58162 8871 58218 8880
rect 58162 8392 58218 8401
rect 58162 8327 58164 8336
rect 58216 8327 58218 8336
rect 58164 8298 58216 8304
rect 57704 7540 57756 7546
rect 57704 7482 57756 7488
rect 58162 7440 58218 7449
rect 58162 7375 58164 7384
rect 58216 7375 58218 7384
rect 58164 7346 58216 7352
rect 57980 7268 58032 7274
rect 57980 7210 58032 7216
rect 57992 7002 58020 7210
rect 57520 6996 57572 7002
rect 57520 6938 57572 6944
rect 57980 6996 58032 7002
rect 57980 6938 58032 6944
rect 57152 6792 57204 6798
rect 57152 6734 57204 6740
rect 57428 6792 57480 6798
rect 57428 6734 57480 6740
rect 57532 6322 57560 6938
rect 57520 6316 57572 6322
rect 57520 6258 57572 6264
rect 58072 6248 58124 6254
rect 58072 6190 58124 6196
rect 57060 6112 57112 6118
rect 57060 6054 57112 6060
rect 57980 6112 58032 6118
rect 57980 6054 58032 6060
rect 56966 5400 57022 5409
rect 56966 5335 56968 5344
rect 57020 5335 57022 5344
rect 56968 5306 57020 5312
rect 57072 5166 57100 6054
rect 57992 5846 58020 6054
rect 57980 5840 58032 5846
rect 57980 5782 58032 5788
rect 57152 5296 57204 5302
rect 57152 5238 57204 5244
rect 57060 5160 57112 5166
rect 57060 5102 57112 5108
rect 57164 4758 57192 5238
rect 57336 5024 57388 5030
rect 57336 4966 57388 4972
rect 57152 4752 57204 4758
rect 57152 4694 57204 4700
rect 57244 4616 57296 4622
rect 57242 4584 57244 4593
rect 57296 4584 57298 4593
rect 57242 4519 57298 4528
rect 56968 4480 57020 4486
rect 56968 4422 57020 4428
rect 56980 4321 57008 4422
rect 56966 4312 57022 4321
rect 56966 4247 57022 4256
rect 57348 4214 57376 4966
rect 57980 4480 58032 4486
rect 57980 4422 58032 4428
rect 57336 4208 57388 4214
rect 57336 4150 57388 4156
rect 57992 4078 58020 4422
rect 57980 4072 58032 4078
rect 57980 4014 58032 4020
rect 57244 3936 57296 3942
rect 57244 3878 57296 3884
rect 56876 3664 56928 3670
rect 56876 3606 56928 3612
rect 56416 3596 56468 3602
rect 56416 3538 56468 3544
rect 56416 3392 56468 3398
rect 56416 3334 56468 3340
rect 56324 2644 56376 2650
rect 56324 2586 56376 2592
rect 56232 2440 56284 2446
rect 56232 2382 56284 2388
rect 55770 2272 55826 2281
rect 55770 2207 55826 2216
rect 56244 1902 56272 2382
rect 56232 1896 56284 1902
rect 56232 1838 56284 1844
rect 55692 870 55812 898
rect 55784 800 55812 870
rect 55218 232 55274 241
rect 55218 167 55274 176
rect 55770 0 55826 800
rect 56428 649 56456 3334
rect 57256 3126 57284 3878
rect 57612 3596 57664 3602
rect 57612 3538 57664 3544
rect 57244 3120 57296 3126
rect 57058 3088 57114 3097
rect 57244 3062 57296 3068
rect 57058 3023 57060 3032
rect 57112 3023 57114 3032
rect 57060 2994 57112 3000
rect 56692 1692 56744 1698
rect 56692 1634 56744 1640
rect 56704 800 56732 1634
rect 57624 800 57652 3538
rect 57980 3392 58032 3398
rect 57980 3334 58032 3340
rect 57992 2582 58020 3334
rect 58084 3194 58112 6190
rect 58162 5808 58218 5817
rect 58162 5743 58164 5752
rect 58216 5743 58218 5752
rect 58164 5714 58216 5720
rect 58164 4004 58216 4010
rect 58164 3946 58216 3952
rect 58072 3188 58124 3194
rect 58072 3130 58124 3136
rect 58176 2825 58204 3946
rect 58532 3120 58584 3126
rect 58532 3062 58584 3068
rect 58162 2816 58218 2825
rect 58162 2751 58218 2760
rect 57980 2576 58032 2582
rect 57980 2518 58032 2524
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 57900 1193 57928 2246
rect 57886 1184 57942 1193
rect 57886 1119 57942 1128
rect 58544 800 58572 3062
rect 59452 2916 59504 2922
rect 59452 2858 59504 2864
rect 59464 800 59492 2858
rect 56414 640 56470 649
rect 56414 575 56470 584
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58530 0 58586 800
rect 59450 0 59506 800
<< via2 >>
rect 2778 59472 2834 59528
rect 1398 57568 1454 57624
rect 1398 56616 1454 56672
rect 2042 58520 2098 58576
rect 56506 59608 56562 59664
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 1398 55664 1454 55720
rect 1398 54732 1454 54768
rect 1398 54712 1400 54732
rect 1400 54712 1452 54732
rect 1452 54712 1454 54732
rect 1398 53760 1454 53816
rect 1398 52808 1454 52864
rect 1398 51892 1400 51912
rect 1400 51892 1452 51912
rect 1452 51892 1454 51912
rect 1398 51856 1454 51892
rect 1398 51040 1454 51096
rect 1398 50088 1454 50144
rect 1398 49136 1454 49192
rect 1398 48204 1454 48240
rect 1398 48184 1400 48204
rect 1400 48184 1452 48204
rect 1452 48184 1454 48204
rect 1398 47232 1454 47288
rect 1398 46280 1454 46336
rect 1398 45364 1400 45384
rect 1400 45364 1452 45384
rect 1452 45364 1454 45384
rect 1398 45328 1454 45364
rect 1398 44376 1454 44432
rect 1398 43424 1454 43480
rect 1398 42608 1454 42664
rect 1398 41676 1454 41712
rect 1398 41656 1400 41676
rect 1400 41656 1452 41676
rect 1452 41656 1454 41676
rect 1398 40704 1454 40760
rect 1398 39752 1454 39808
rect 1398 38836 1400 38856
rect 1400 38836 1452 38856
rect 1452 38836 1454 38856
rect 1398 38800 1454 38836
rect 1398 37848 1454 37904
rect 1398 36896 1454 36952
rect 1398 35944 1454 36000
rect 1398 34992 1454 35048
rect 1398 34176 1454 34232
rect 1398 33224 1454 33280
rect 1398 32308 1400 32328
rect 1400 32308 1452 32328
rect 1452 32308 1454 32328
rect 1398 32272 1454 32308
rect 1398 31320 1454 31376
rect 1398 30368 1454 30424
rect 1950 29416 2006 29472
rect 1398 28464 1454 28520
rect 1950 27512 2006 27568
rect 1950 26560 2006 26616
rect 2042 25764 2098 25800
rect 2042 25744 2044 25764
rect 2044 25744 2096 25764
rect 2096 25744 2098 25764
rect 2778 24812 2834 24848
rect 2778 24792 2780 24812
rect 2780 24792 2832 24812
rect 2832 24792 2834 24812
rect 1950 23840 2006 23896
rect 1950 22924 1952 22944
rect 1952 22924 2004 22944
rect 2004 22924 2006 22944
rect 1950 22888 2006 22924
rect 2042 21956 2098 21992
rect 2042 21936 2044 21956
rect 2044 21936 2096 21956
rect 2096 21936 2098 21956
rect 2778 21004 2834 21040
rect 2778 20984 2780 21004
rect 2780 20984 2832 21004
rect 2832 20984 2834 21004
rect 1950 20032 2006 20088
rect 2778 19080 2834 19136
rect 1950 18128 2006 18184
rect 1950 17312 2006 17368
rect 1950 16396 1952 16416
rect 1952 16396 2004 16416
rect 2004 16396 2006 16416
rect 1950 16360 2006 16396
rect 2778 15428 2834 15464
rect 2778 15408 2780 15428
rect 2780 15408 2832 15428
rect 2832 15408 2834 15428
rect 1950 14456 2006 14512
rect 1950 13504 2006 13560
rect 1950 12588 1952 12608
rect 1952 12588 2004 12608
rect 2004 12588 2006 12608
rect 1950 12552 2006 12588
rect 2778 11620 2834 11656
rect 2778 11600 2780 11620
rect 2780 11600 2832 11620
rect 2832 11600 2834 11620
rect 1950 10648 2006 10704
rect 1950 9696 2006 9752
rect 2778 8880 2834 8936
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 50300 57146 50356 57148
rect 50380 57146 50436 57148
rect 50460 57146 50516 57148
rect 50540 57146 50596 57148
rect 50300 57094 50326 57146
rect 50326 57094 50356 57146
rect 50380 57094 50390 57146
rect 50390 57094 50436 57146
rect 50460 57094 50506 57146
rect 50506 57094 50516 57146
rect 50540 57094 50570 57146
rect 50570 57094 50596 57146
rect 50300 57092 50356 57094
rect 50380 57092 50436 57094
rect 50460 57092 50516 57094
rect 50540 57092 50596 57094
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 50300 56058 50356 56060
rect 50380 56058 50436 56060
rect 50460 56058 50516 56060
rect 50540 56058 50596 56060
rect 50300 56006 50326 56058
rect 50326 56006 50356 56058
rect 50380 56006 50390 56058
rect 50390 56006 50436 56058
rect 50460 56006 50506 56058
rect 50506 56006 50516 56058
rect 50540 56006 50570 56058
rect 50570 56006 50596 56058
rect 50300 56004 50356 56006
rect 50380 56004 50436 56006
rect 50460 56004 50516 56006
rect 50540 56004 50596 56006
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 55034 58384 55090 58440
rect 54942 58112 54998 58168
rect 56322 59064 56378 59120
rect 55494 58520 55550 58576
rect 56322 58384 56378 58440
rect 56506 58112 56562 58168
rect 56506 57976 56562 58032
rect 55586 57432 55642 57488
rect 55678 55936 55734 55992
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 50300 54970 50356 54972
rect 50380 54970 50436 54972
rect 50460 54970 50516 54972
rect 50540 54970 50596 54972
rect 50300 54918 50326 54970
rect 50326 54918 50356 54970
rect 50380 54918 50390 54970
rect 50390 54918 50436 54970
rect 50460 54918 50506 54970
rect 50506 54918 50516 54970
rect 50540 54918 50570 54970
rect 50570 54918 50596 54970
rect 50300 54916 50356 54918
rect 50380 54916 50436 54918
rect 50460 54916 50516 54918
rect 50540 54916 50596 54918
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 50300 53882 50356 53884
rect 50380 53882 50436 53884
rect 50460 53882 50516 53884
rect 50540 53882 50596 53884
rect 50300 53830 50326 53882
rect 50326 53830 50356 53882
rect 50380 53830 50390 53882
rect 50390 53830 50436 53882
rect 50460 53830 50506 53882
rect 50506 53830 50516 53882
rect 50540 53830 50570 53882
rect 50570 53830 50596 53882
rect 50300 53828 50356 53830
rect 50380 53828 50436 53830
rect 50460 53828 50516 53830
rect 50540 53828 50596 53830
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 50300 52794 50356 52796
rect 50380 52794 50436 52796
rect 50460 52794 50516 52796
rect 50540 52794 50596 52796
rect 50300 52742 50326 52794
rect 50326 52742 50356 52794
rect 50380 52742 50390 52794
rect 50390 52742 50436 52794
rect 50460 52742 50506 52794
rect 50506 52742 50516 52794
rect 50540 52742 50570 52794
rect 50570 52742 50596 52794
rect 50300 52740 50356 52742
rect 50380 52740 50436 52742
rect 50460 52740 50516 52742
rect 50540 52740 50596 52742
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 50300 51706 50356 51708
rect 50380 51706 50436 51708
rect 50460 51706 50516 51708
rect 50540 51706 50596 51708
rect 50300 51654 50326 51706
rect 50326 51654 50356 51706
rect 50380 51654 50390 51706
rect 50390 51654 50436 51706
rect 50460 51654 50506 51706
rect 50506 51654 50516 51706
rect 50540 51654 50570 51706
rect 50570 51654 50596 51706
rect 50300 51652 50356 51654
rect 50380 51652 50436 51654
rect 50460 51652 50516 51654
rect 50540 51652 50596 51654
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 50300 50618 50356 50620
rect 50380 50618 50436 50620
rect 50460 50618 50516 50620
rect 50540 50618 50596 50620
rect 50300 50566 50326 50618
rect 50326 50566 50356 50618
rect 50380 50566 50390 50618
rect 50390 50566 50436 50618
rect 50460 50566 50506 50618
rect 50506 50566 50516 50618
rect 50540 50566 50570 50618
rect 50570 50566 50596 50618
rect 50300 50564 50356 50566
rect 50380 50564 50436 50566
rect 50460 50564 50516 50566
rect 50540 50564 50596 50566
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 55218 49716 55220 49736
rect 55220 49716 55272 49736
rect 55272 49716 55274 49736
rect 55218 49680 55274 49716
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 50300 49530 50356 49532
rect 50380 49530 50436 49532
rect 50460 49530 50516 49532
rect 50540 49530 50596 49532
rect 50300 49478 50326 49530
rect 50326 49478 50356 49530
rect 50380 49478 50390 49530
rect 50390 49478 50436 49530
rect 50460 49478 50506 49530
rect 50506 49478 50516 49530
rect 50540 49478 50570 49530
rect 50570 49478 50596 49530
rect 50300 49476 50356 49478
rect 50380 49476 50436 49478
rect 50460 49476 50516 49478
rect 50540 49476 50596 49478
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 50300 48442 50356 48444
rect 50380 48442 50436 48444
rect 50460 48442 50516 48444
rect 50540 48442 50596 48444
rect 50300 48390 50326 48442
rect 50326 48390 50356 48442
rect 50380 48390 50390 48442
rect 50390 48390 50436 48442
rect 50460 48390 50506 48442
rect 50506 48390 50516 48442
rect 50540 48390 50570 48442
rect 50570 48390 50596 48442
rect 50300 48388 50356 48390
rect 50380 48388 50436 48390
rect 50460 48388 50516 48390
rect 50540 48388 50596 48390
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 50300 47354 50356 47356
rect 50380 47354 50436 47356
rect 50460 47354 50516 47356
rect 50540 47354 50596 47356
rect 50300 47302 50326 47354
rect 50326 47302 50356 47354
rect 50380 47302 50390 47354
rect 50390 47302 50436 47354
rect 50460 47302 50506 47354
rect 50506 47302 50516 47354
rect 50540 47302 50570 47354
rect 50570 47302 50596 47354
rect 50300 47300 50356 47302
rect 50380 47300 50436 47302
rect 50460 47300 50516 47302
rect 50540 47300 50596 47302
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 55218 46688 55274 46744
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 50300 46266 50356 46268
rect 50380 46266 50436 46268
rect 50460 46266 50516 46268
rect 50540 46266 50596 46268
rect 50300 46214 50326 46266
rect 50326 46214 50356 46266
rect 50380 46214 50390 46266
rect 50390 46214 50436 46266
rect 50460 46214 50506 46266
rect 50506 46214 50516 46266
rect 50540 46214 50570 46266
rect 50570 46214 50596 46266
rect 50300 46212 50356 46214
rect 50380 46212 50436 46214
rect 50460 46212 50516 46214
rect 50540 46212 50596 46214
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 50300 45178 50356 45180
rect 50380 45178 50436 45180
rect 50460 45178 50516 45180
rect 50540 45178 50596 45180
rect 50300 45126 50326 45178
rect 50326 45126 50356 45178
rect 50380 45126 50390 45178
rect 50390 45126 50436 45178
rect 50460 45126 50506 45178
rect 50506 45126 50516 45178
rect 50540 45126 50570 45178
rect 50570 45126 50596 45178
rect 50300 45124 50356 45126
rect 50380 45124 50436 45126
rect 50460 45124 50516 45126
rect 50540 45124 50596 45126
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 50434 42236 50436 42256
rect 50436 42236 50488 42256
rect 50488 42236 50490 42256
rect 50434 42200 50490 42236
rect 49422 42100 49424 42120
rect 49424 42100 49476 42120
rect 49476 42100 49478 42120
rect 49422 42064 49478 42100
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 49790 37204 49792 37224
rect 49792 37204 49844 37224
rect 49844 37204 49846 37224
rect 49790 37168 49846 37204
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 52182 42236 52184 42256
rect 52184 42236 52236 42256
rect 52236 42236 52238 42256
rect 52182 42200 52238 42236
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50710 38548 50766 38584
rect 50710 38528 50712 38548
rect 50712 38528 50764 38548
rect 50764 38528 50766 38548
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 52550 38956 52606 38992
rect 52550 38936 52552 38956
rect 52552 38936 52604 38956
rect 52604 38936 52606 38956
rect 52458 38392 52514 38448
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 49882 35148 49938 35184
rect 49882 35128 49884 35148
rect 49884 35128 49936 35148
rect 49936 35128 49938 35148
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 49698 32680 49754 32736
rect 50342 34584 50398 34640
rect 50618 34448 50674 34504
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 51906 37032 51962 37088
rect 50802 34040 50858 34096
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 49514 29164 49570 29200
rect 49514 29144 49516 29164
rect 49516 29144 49568 29164
rect 49568 29144 49570 29164
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 48410 26424 48466 26480
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 49606 25336 49662 25392
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 50710 30932 50766 30968
rect 50710 30912 50712 30932
rect 50712 30912 50764 30932
rect 50764 30912 50766 30932
rect 50526 30796 50582 30832
rect 50526 30776 50528 30796
rect 50528 30776 50580 30796
rect 50580 30776 50582 30796
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 50300 28858 50356 28860
rect 50380 28858 50436 28860
rect 50460 28858 50516 28860
rect 50540 28858 50596 28860
rect 50300 28806 50326 28858
rect 50326 28806 50356 28858
rect 50380 28806 50390 28858
rect 50390 28806 50436 28858
rect 50460 28806 50506 28858
rect 50506 28806 50516 28858
rect 50540 28806 50570 28858
rect 50570 28806 50596 28858
rect 50300 28804 50356 28806
rect 50380 28804 50436 28806
rect 50460 28804 50516 28806
rect 50540 28804 50596 28806
rect 50710 28600 50766 28656
rect 50300 27770 50356 27772
rect 50380 27770 50436 27772
rect 50460 27770 50516 27772
rect 50540 27770 50596 27772
rect 50300 27718 50326 27770
rect 50326 27718 50356 27770
rect 50380 27718 50390 27770
rect 50390 27718 50436 27770
rect 50460 27718 50506 27770
rect 50506 27718 50516 27770
rect 50540 27718 50570 27770
rect 50570 27718 50596 27770
rect 50300 27716 50356 27718
rect 50380 27716 50436 27718
rect 50460 27716 50516 27718
rect 50540 27716 50596 27718
rect 50250 27548 50252 27568
rect 50252 27548 50304 27568
rect 50304 27548 50306 27568
rect 50250 27512 50306 27548
rect 52642 37032 52698 37088
rect 55034 45056 55090 45112
rect 54758 43560 54814 43616
rect 53286 38956 53342 38992
rect 53286 38936 53288 38956
rect 53288 38936 53340 38956
rect 53340 38936 53342 38956
rect 53378 38392 53434 38448
rect 54206 38548 54262 38584
rect 54206 38528 54208 38548
rect 54208 38528 54260 38548
rect 54260 38528 54262 38548
rect 50300 26682 50356 26684
rect 50380 26682 50436 26684
rect 50460 26682 50516 26684
rect 50540 26682 50596 26684
rect 50300 26630 50326 26682
rect 50326 26630 50356 26682
rect 50380 26630 50390 26682
rect 50390 26630 50436 26682
rect 50460 26630 50506 26682
rect 50506 26630 50516 26682
rect 50540 26630 50570 26682
rect 50570 26630 50596 26682
rect 50300 26628 50356 26630
rect 50380 26628 50436 26630
rect 50460 26628 50516 26630
rect 50540 26628 50596 26630
rect 50300 25594 50356 25596
rect 50380 25594 50436 25596
rect 50460 25594 50516 25596
rect 50540 25594 50596 25596
rect 50300 25542 50326 25594
rect 50326 25542 50356 25594
rect 50380 25542 50390 25594
rect 50390 25542 50436 25594
rect 50460 25542 50506 25594
rect 50506 25542 50516 25594
rect 50540 25542 50570 25594
rect 50570 25542 50596 25594
rect 50300 25540 50356 25542
rect 50380 25540 50436 25542
rect 50460 25540 50516 25542
rect 50540 25540 50596 25542
rect 50300 24506 50356 24508
rect 50380 24506 50436 24508
rect 50460 24506 50516 24508
rect 50540 24506 50596 24508
rect 50300 24454 50326 24506
rect 50326 24454 50356 24506
rect 50380 24454 50390 24506
rect 50390 24454 50436 24506
rect 50460 24454 50506 24506
rect 50506 24454 50516 24506
rect 50540 24454 50570 24506
rect 50570 24454 50596 24506
rect 50300 24452 50356 24454
rect 50380 24452 50436 24454
rect 50460 24452 50516 24454
rect 50540 24452 50596 24454
rect 50300 23418 50356 23420
rect 50380 23418 50436 23420
rect 50460 23418 50516 23420
rect 50540 23418 50596 23420
rect 50300 23366 50326 23418
rect 50326 23366 50356 23418
rect 50380 23366 50390 23418
rect 50390 23366 50436 23418
rect 50460 23366 50506 23418
rect 50506 23366 50516 23418
rect 50540 23366 50570 23418
rect 50570 23366 50596 23418
rect 50300 23364 50356 23366
rect 50380 23364 50436 23366
rect 50460 23364 50516 23366
rect 50540 23364 50596 23366
rect 50434 23196 50436 23216
rect 50436 23196 50488 23216
rect 50488 23196 50490 23216
rect 50434 23160 50490 23196
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 2042 7928 2098 7984
rect 1950 6976 2006 7032
rect 1950 6060 1952 6080
rect 1952 6060 2004 6080
rect 2004 6060 2006 6080
rect 1950 6024 2006 6060
rect 2778 5108 2780 5128
rect 2780 5108 2832 5128
rect 2832 5108 2834 5128
rect 2778 5072 2834 5108
rect 2870 4120 2926 4176
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 2778 3168 2834 3224
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 50300 22330 50356 22332
rect 50380 22330 50436 22332
rect 50460 22330 50516 22332
rect 50540 22330 50596 22332
rect 50300 22278 50326 22330
rect 50326 22278 50356 22330
rect 50380 22278 50390 22330
rect 50390 22278 50436 22330
rect 50460 22278 50506 22330
rect 50506 22278 50516 22330
rect 50540 22278 50570 22330
rect 50570 22278 50596 22330
rect 50300 22276 50356 22278
rect 50380 22276 50436 22278
rect 50460 22276 50516 22278
rect 50540 22276 50596 22278
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 48410 19896 48466 19952
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 49698 15564 49754 15600
rect 49698 15544 49700 15564
rect 49700 15544 49752 15564
rect 49752 15544 49754 15564
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 49882 17040 49938 17096
rect 50300 21242 50356 21244
rect 50380 21242 50436 21244
rect 50460 21242 50516 21244
rect 50540 21242 50596 21244
rect 50300 21190 50326 21242
rect 50326 21190 50356 21242
rect 50380 21190 50390 21242
rect 50390 21190 50436 21242
rect 50460 21190 50506 21242
rect 50506 21190 50516 21242
rect 50540 21190 50570 21242
rect 50570 21190 50596 21242
rect 50300 21188 50356 21190
rect 50380 21188 50436 21190
rect 50460 21188 50516 21190
rect 50540 21188 50596 21190
rect 50300 20154 50356 20156
rect 50380 20154 50436 20156
rect 50460 20154 50516 20156
rect 50540 20154 50596 20156
rect 50300 20102 50326 20154
rect 50326 20102 50356 20154
rect 50380 20102 50390 20154
rect 50390 20102 50436 20154
rect 50460 20102 50506 20154
rect 50506 20102 50516 20154
rect 50540 20102 50570 20154
rect 50570 20102 50596 20154
rect 50300 20100 50356 20102
rect 50380 20100 50436 20102
rect 50460 20100 50516 20102
rect 50540 20100 50596 20102
rect 50300 19066 50356 19068
rect 50380 19066 50436 19068
rect 50460 19066 50516 19068
rect 50540 19066 50596 19068
rect 50300 19014 50326 19066
rect 50326 19014 50356 19066
rect 50380 19014 50390 19066
rect 50390 19014 50436 19066
rect 50460 19014 50506 19066
rect 50506 19014 50516 19066
rect 50540 19014 50570 19066
rect 50570 19014 50596 19066
rect 50300 19012 50356 19014
rect 50380 19012 50436 19014
rect 50460 19012 50516 19014
rect 50540 19012 50596 19014
rect 50618 18808 50674 18864
rect 50158 18400 50214 18456
rect 50300 17978 50356 17980
rect 50380 17978 50436 17980
rect 50460 17978 50516 17980
rect 50540 17978 50596 17980
rect 50300 17926 50326 17978
rect 50326 17926 50356 17978
rect 50380 17926 50390 17978
rect 50390 17926 50436 17978
rect 50460 17926 50506 17978
rect 50506 17926 50516 17978
rect 50540 17926 50570 17978
rect 50570 17926 50596 17978
rect 50300 17924 50356 17926
rect 50380 17924 50436 17926
rect 50460 17924 50516 17926
rect 50540 17924 50596 17926
rect 50526 17312 50582 17368
rect 50300 16890 50356 16892
rect 50380 16890 50436 16892
rect 50460 16890 50516 16892
rect 50540 16890 50596 16892
rect 50300 16838 50326 16890
rect 50326 16838 50356 16890
rect 50380 16838 50390 16890
rect 50390 16838 50436 16890
rect 50460 16838 50506 16890
rect 50506 16838 50516 16890
rect 50540 16838 50570 16890
rect 50570 16838 50596 16890
rect 50300 16836 50356 16838
rect 50380 16836 50436 16838
rect 50460 16836 50516 16838
rect 50540 16836 50596 16838
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 49146 14048 49202 14104
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 2870 1264 2926 1320
rect 4066 2216 4122 2272
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 45006 4528 45062 4584
rect 47214 3984 47270 4040
rect 49330 11620 49386 11656
rect 49330 11600 49332 11620
rect 49332 11600 49384 11620
rect 49384 11600 49386 11620
rect 48686 7792 48742 7848
rect 48410 7656 48466 7712
rect 48778 6860 48834 6896
rect 48778 6840 48780 6860
rect 48780 6840 48832 6860
rect 48832 6840 48834 6860
rect 48686 6740 48688 6760
rect 48688 6740 48740 6760
rect 48740 6740 48742 6760
rect 48686 6704 48742 6740
rect 48134 4548 48190 4584
rect 48134 4528 48136 4548
rect 48136 4528 48188 4548
rect 48188 4528 48190 4548
rect 49330 7928 49386 7984
rect 50300 15802 50356 15804
rect 50380 15802 50436 15804
rect 50460 15802 50516 15804
rect 50540 15802 50596 15804
rect 50300 15750 50326 15802
rect 50326 15750 50356 15802
rect 50380 15750 50390 15802
rect 50390 15750 50436 15802
rect 50460 15750 50506 15802
rect 50506 15750 50516 15802
rect 50540 15750 50570 15802
rect 50570 15750 50596 15802
rect 50300 15748 50356 15750
rect 50380 15748 50436 15750
rect 50460 15748 50516 15750
rect 50540 15748 50596 15750
rect 50300 14714 50356 14716
rect 50380 14714 50436 14716
rect 50460 14714 50516 14716
rect 50540 14714 50596 14716
rect 50300 14662 50326 14714
rect 50326 14662 50356 14714
rect 50380 14662 50390 14714
rect 50390 14662 50436 14714
rect 50460 14662 50506 14714
rect 50506 14662 50516 14714
rect 50540 14662 50570 14714
rect 50570 14662 50596 14714
rect 50300 14660 50356 14662
rect 50380 14660 50436 14662
rect 50460 14660 50516 14662
rect 50540 14660 50596 14662
rect 50434 14456 50490 14512
rect 49698 6840 49754 6896
rect 50300 13626 50356 13628
rect 50380 13626 50436 13628
rect 50460 13626 50516 13628
rect 50540 13626 50596 13628
rect 50300 13574 50326 13626
rect 50326 13574 50356 13626
rect 50380 13574 50390 13626
rect 50390 13574 50436 13626
rect 50460 13574 50506 13626
rect 50506 13574 50516 13626
rect 50540 13574 50570 13626
rect 50570 13574 50596 13626
rect 50300 13572 50356 13574
rect 50380 13572 50436 13574
rect 50460 13572 50516 13574
rect 50540 13572 50596 13574
rect 50300 12538 50356 12540
rect 50380 12538 50436 12540
rect 50460 12538 50516 12540
rect 50540 12538 50596 12540
rect 50300 12486 50326 12538
rect 50326 12486 50356 12538
rect 50380 12486 50390 12538
rect 50390 12486 50436 12538
rect 50460 12486 50506 12538
rect 50506 12486 50516 12538
rect 50540 12486 50570 12538
rect 50570 12486 50596 12538
rect 50300 12484 50356 12486
rect 50380 12484 50436 12486
rect 50460 12484 50516 12486
rect 50540 12484 50596 12486
rect 50710 18536 50766 18592
rect 52550 33496 52606 33552
rect 51814 31884 51870 31920
rect 51814 31864 51816 31884
rect 51816 31864 51868 31884
rect 51868 31864 51870 31884
rect 50710 13640 50766 13696
rect 50526 12300 50582 12336
rect 50526 12280 50528 12300
rect 50528 12280 50580 12300
rect 50580 12280 50582 12300
rect 51078 18944 51134 19000
rect 51262 18536 51318 18592
rect 53286 33804 53288 33824
rect 53288 33804 53340 33824
rect 53340 33804 53342 33824
rect 53286 33768 53342 33804
rect 52182 28620 52238 28656
rect 52182 28600 52184 28620
rect 52184 28600 52236 28620
rect 52236 28600 52238 28620
rect 51906 25880 51962 25936
rect 51722 22772 51778 22808
rect 51722 22752 51724 22772
rect 51724 22752 51776 22772
rect 51776 22752 51778 22772
rect 51630 20848 51686 20904
rect 51998 20440 52054 20496
rect 51538 19352 51594 19408
rect 51814 18808 51870 18864
rect 51354 17620 51356 17640
rect 51356 17620 51408 17640
rect 51408 17620 51410 17640
rect 51354 17584 51410 17620
rect 51446 17312 51502 17368
rect 52090 17448 52146 17504
rect 50986 14184 51042 14240
rect 50986 13912 51042 13968
rect 50300 11450 50356 11452
rect 50380 11450 50436 11452
rect 50460 11450 50516 11452
rect 50540 11450 50596 11452
rect 50300 11398 50326 11450
rect 50326 11398 50356 11450
rect 50380 11398 50390 11450
rect 50390 11398 50436 11450
rect 50460 11398 50506 11450
rect 50506 11398 50516 11450
rect 50540 11398 50570 11450
rect 50570 11398 50596 11450
rect 50300 11396 50356 11398
rect 50380 11396 50436 11398
rect 50460 11396 50516 11398
rect 50540 11396 50596 11398
rect 50300 10362 50356 10364
rect 50380 10362 50436 10364
rect 50460 10362 50516 10364
rect 50540 10362 50596 10364
rect 50300 10310 50326 10362
rect 50326 10310 50356 10362
rect 50380 10310 50390 10362
rect 50390 10310 50436 10362
rect 50460 10310 50506 10362
rect 50506 10310 50516 10362
rect 50540 10310 50570 10362
rect 50570 10310 50596 10362
rect 50300 10308 50356 10310
rect 50380 10308 50436 10310
rect 50460 10308 50516 10310
rect 50540 10308 50596 10310
rect 50300 9274 50356 9276
rect 50380 9274 50436 9276
rect 50460 9274 50516 9276
rect 50540 9274 50596 9276
rect 50300 9222 50326 9274
rect 50326 9222 50356 9274
rect 50380 9222 50390 9274
rect 50390 9222 50436 9274
rect 50460 9222 50506 9274
rect 50506 9222 50516 9274
rect 50540 9222 50570 9274
rect 50570 9222 50596 9274
rect 50300 9220 50356 9222
rect 50380 9220 50436 9222
rect 50460 9220 50516 9222
rect 50540 9220 50596 9222
rect 49790 6704 49846 6760
rect 49238 5108 49240 5128
rect 49240 5108 49292 5128
rect 49292 5108 49294 5128
rect 49238 5072 49294 5108
rect 49146 3304 49202 3360
rect 49606 5772 49662 5808
rect 49606 5752 49608 5772
rect 49608 5752 49660 5772
rect 49660 5752 49662 5772
rect 49422 5208 49478 5264
rect 49606 3032 49662 3088
rect 50300 8186 50356 8188
rect 50380 8186 50436 8188
rect 50460 8186 50516 8188
rect 50540 8186 50596 8188
rect 50300 8134 50326 8186
rect 50326 8134 50356 8186
rect 50380 8134 50390 8186
rect 50390 8134 50436 8186
rect 50460 8134 50506 8186
rect 50506 8134 50516 8186
rect 50540 8134 50570 8186
rect 50570 8134 50596 8186
rect 50300 8132 50356 8134
rect 50380 8132 50436 8134
rect 50460 8132 50516 8134
rect 50540 8132 50596 8134
rect 50300 7098 50356 7100
rect 50380 7098 50436 7100
rect 50460 7098 50516 7100
rect 50540 7098 50596 7100
rect 50300 7046 50326 7098
rect 50326 7046 50356 7098
rect 50380 7046 50390 7098
rect 50390 7046 50436 7098
rect 50460 7046 50506 7098
rect 50506 7046 50516 7098
rect 50540 7046 50570 7098
rect 50570 7046 50596 7098
rect 50300 7044 50356 7046
rect 50380 7044 50436 7046
rect 50460 7044 50516 7046
rect 50540 7044 50596 7046
rect 49974 5480 50030 5536
rect 55218 40432 55274 40488
rect 55218 38972 55220 38992
rect 55220 38972 55272 38992
rect 55272 38972 55274 38992
rect 55218 38936 55274 38972
rect 55218 37304 55274 37360
rect 54390 35436 54392 35456
rect 54392 35436 54444 35456
rect 54444 35436 54446 35456
rect 54390 35400 54446 35436
rect 55218 35828 55274 35864
rect 55218 35808 55220 35828
rect 55220 35808 55272 35828
rect 55272 35808 55274 35828
rect 54942 35128 54998 35184
rect 54574 34312 54630 34368
rect 55218 34176 55274 34232
rect 57058 56480 57114 56536
rect 55494 54440 55550 54496
rect 57058 54848 57114 54904
rect 58162 57024 58218 57080
rect 58162 55392 58218 55448
rect 56966 53352 57022 53408
rect 58162 53896 58218 53952
rect 55586 52808 55642 52864
rect 55494 51312 55550 51368
rect 57058 51876 57114 51912
rect 57886 52264 57942 52320
rect 57058 51856 57060 51876
rect 57060 51856 57112 51876
rect 57112 51856 57114 51876
rect 57058 50244 57114 50280
rect 57058 50224 57060 50244
rect 57060 50224 57112 50244
rect 57112 50224 57114 50244
rect 55494 48184 55550 48240
rect 58162 50788 58218 50824
rect 58162 50768 58164 50788
rect 58164 50768 58216 50788
rect 58216 50768 58218 50788
rect 58162 49292 58218 49328
rect 58162 49272 58164 49292
rect 58164 49272 58216 49292
rect 58216 49272 58218 49292
rect 57058 48764 57060 48784
rect 57060 48764 57112 48784
rect 57112 48764 57114 48784
rect 57058 48728 57114 48764
rect 57058 47660 57114 47696
rect 57058 47640 57060 47660
rect 57060 47640 57112 47660
rect 57112 47640 57114 47660
rect 57426 47116 57482 47152
rect 57426 47096 57428 47116
rect 57428 47096 57480 47116
rect 57480 47096 57482 47116
rect 55494 34312 55550 34368
rect 54758 33768 54814 33824
rect 54666 33496 54722 33552
rect 53838 31864 53894 31920
rect 53654 30796 53710 30832
rect 53654 30776 53656 30796
rect 53656 30776 53708 30796
rect 53708 30776 53710 30796
rect 53838 30796 53894 30832
rect 53838 30776 53840 30796
rect 53840 30776 53892 30796
rect 53892 30776 53894 30796
rect 55402 33768 55458 33824
rect 55586 33496 55642 33552
rect 54758 30796 54814 30832
rect 54758 30776 54760 30796
rect 54760 30776 54812 30796
rect 54812 30776 54814 30796
rect 52918 26444 52974 26480
rect 52918 26424 52920 26444
rect 52920 26424 52972 26444
rect 52972 26424 52974 26444
rect 55218 31204 55274 31240
rect 55218 31184 55220 31204
rect 55220 31184 55272 31204
rect 55272 31184 55274 31204
rect 52734 22752 52790 22808
rect 54206 27512 54262 27568
rect 55494 29552 55550 29608
rect 55310 28056 55366 28112
rect 55218 24948 55274 24984
rect 55218 24928 55220 24948
rect 55220 24928 55272 24948
rect 55272 24928 55274 24948
rect 52642 21004 52698 21040
rect 52642 20984 52644 21004
rect 52644 20984 52696 21004
rect 52696 20984 52698 21004
rect 52550 19236 52606 19272
rect 52550 19216 52552 19236
rect 52552 19216 52604 19236
rect 52604 19216 52606 19236
rect 52274 18808 52330 18864
rect 53102 19916 53158 19952
rect 53102 19896 53104 19916
rect 53104 19896 53156 19916
rect 53156 19896 53158 19916
rect 53010 19760 53066 19816
rect 55218 23432 55274 23488
rect 54298 21004 54354 21040
rect 54298 20984 54300 21004
rect 54300 20984 54352 21004
rect 54352 20984 54354 21004
rect 53286 20460 53342 20496
rect 53286 20440 53288 20460
rect 53288 20440 53340 20460
rect 53340 20440 53342 20460
rect 53194 18808 53250 18864
rect 53378 19216 53434 19272
rect 53102 17720 53158 17776
rect 54666 19896 54722 19952
rect 55494 26424 55550 26480
rect 55218 21836 55220 21856
rect 55220 21836 55272 21856
rect 55272 21836 55274 21856
rect 55218 21800 55274 21836
rect 54574 19760 54630 19816
rect 54758 19352 54814 19408
rect 57058 45600 57114 45656
rect 57886 46144 57942 46200
rect 57058 44104 57114 44160
rect 58162 44512 58218 44568
rect 56966 42508 56968 42528
rect 56968 42508 57020 42528
rect 57020 42508 57022 42528
rect 56966 42472 57022 42508
rect 58162 43016 58218 43072
rect 58162 41520 58218 41576
rect 57426 40996 57482 41032
rect 57426 40976 57428 40996
rect 57428 40976 57480 40996
rect 57480 40976 57482 40996
rect 56966 39364 57022 39400
rect 56966 39344 56968 39364
rect 56968 39344 57020 39364
rect 57020 39344 57022 39364
rect 57886 39888 57942 39944
rect 57058 37204 57060 37224
rect 57060 37204 57112 37224
rect 57112 37204 57114 37224
rect 57058 37168 57114 37204
rect 57886 37848 57942 37904
rect 56966 36372 57022 36408
rect 56966 36352 56968 36372
rect 56968 36352 57020 36372
rect 57020 36352 57022 36372
rect 56598 35436 56600 35456
rect 56600 35436 56652 35456
rect 56652 35436 56654 35456
rect 56598 35400 56654 35436
rect 56414 34720 56470 34776
rect 58162 38412 58218 38448
rect 58162 38392 58164 38412
rect 58164 38392 58216 38412
rect 58216 38392 58218 38412
rect 58162 36780 58218 36816
rect 58162 36760 58164 36780
rect 58164 36760 58216 36780
rect 58216 36760 58218 36780
rect 56966 35284 57022 35320
rect 56966 35264 56968 35284
rect 56968 35264 57020 35284
rect 57020 35264 57022 35284
rect 57058 34604 57114 34640
rect 57058 34584 57060 34604
rect 57060 34584 57112 34604
rect 57112 34584 57114 34604
rect 56874 34484 56876 34504
rect 56876 34484 56928 34504
rect 56928 34484 56930 34504
rect 56874 34448 56930 34484
rect 56782 34076 56784 34096
rect 56784 34076 56836 34096
rect 56836 34076 56838 34096
rect 56782 34040 56838 34076
rect 57334 33260 57336 33280
rect 57336 33260 57388 33280
rect 57388 33260 57390 33280
rect 57334 33224 57390 33260
rect 55954 29144 56010 29200
rect 57426 31592 57482 31648
rect 57426 30912 57482 30968
rect 56690 25356 56746 25392
rect 56690 25336 56692 25356
rect 56692 25336 56744 25356
rect 56744 25336 56746 25356
rect 55494 20848 55550 20904
rect 55310 20304 55366 20360
rect 55218 18672 55274 18728
rect 52826 16496 52882 16552
rect 52550 14456 52606 14512
rect 52366 13912 52422 13968
rect 52550 13812 52552 13832
rect 52552 13812 52604 13832
rect 52604 13812 52606 13832
rect 52550 13776 52606 13812
rect 53194 16632 53250 16688
rect 53930 17448 53986 17504
rect 54942 17740 54998 17776
rect 54942 17720 54944 17740
rect 54944 17720 54996 17740
rect 54996 17720 54998 17740
rect 54022 17312 54078 17368
rect 54758 17584 54814 17640
rect 54206 16652 54262 16688
rect 54206 16632 54208 16652
rect 54208 16632 54260 16652
rect 54260 16632 54262 16652
rect 52274 12300 52330 12336
rect 52274 12280 52276 12300
rect 52276 12280 52328 12300
rect 52328 12280 52330 12300
rect 53930 14456 53986 14512
rect 54482 16496 54538 16552
rect 55218 17176 55274 17232
rect 55678 17332 55734 17368
rect 55678 17312 55680 17332
rect 55680 17312 55732 17332
rect 55732 17312 55734 17332
rect 55218 13776 55274 13832
rect 50300 6010 50356 6012
rect 50380 6010 50436 6012
rect 50460 6010 50516 6012
rect 50540 6010 50596 6012
rect 50300 5958 50326 6010
rect 50326 5958 50356 6010
rect 50380 5958 50390 6010
rect 50390 5958 50436 6010
rect 50460 5958 50506 6010
rect 50506 5958 50516 6010
rect 50540 5958 50570 6010
rect 50570 5958 50596 6010
rect 50300 5956 50356 5958
rect 50380 5956 50436 5958
rect 50460 5956 50516 5958
rect 50540 5956 50596 5958
rect 50300 4922 50356 4924
rect 50380 4922 50436 4924
rect 50460 4922 50516 4924
rect 50540 4922 50596 4924
rect 50300 4870 50326 4922
rect 50326 4870 50356 4922
rect 50380 4870 50390 4922
rect 50390 4870 50436 4922
rect 50460 4870 50506 4922
rect 50506 4870 50516 4922
rect 50540 4870 50570 4922
rect 50570 4870 50596 4922
rect 50300 4868 50356 4870
rect 50380 4868 50436 4870
rect 50460 4868 50516 4870
rect 50540 4868 50596 4870
rect 50710 4564 50712 4584
rect 50712 4564 50764 4584
rect 50764 4564 50766 4584
rect 50710 4528 50766 4564
rect 50066 4120 50122 4176
rect 50300 3834 50356 3836
rect 50380 3834 50436 3836
rect 50460 3834 50516 3836
rect 50540 3834 50596 3836
rect 50300 3782 50326 3834
rect 50326 3782 50356 3834
rect 50380 3782 50390 3834
rect 50390 3782 50436 3834
rect 50460 3782 50506 3834
rect 50506 3782 50516 3834
rect 50540 3782 50570 3834
rect 50570 3782 50596 3834
rect 50300 3780 50356 3782
rect 50380 3780 50436 3782
rect 50460 3780 50516 3782
rect 50540 3780 50596 3782
rect 50300 2746 50356 2748
rect 50380 2746 50436 2748
rect 50460 2746 50516 2748
rect 50540 2746 50596 2748
rect 50300 2694 50326 2746
rect 50326 2694 50356 2746
rect 50380 2694 50390 2746
rect 50390 2694 50436 2746
rect 50460 2694 50506 2746
rect 50506 2694 50516 2746
rect 50540 2694 50570 2746
rect 50570 2694 50596 2746
rect 50300 2692 50356 2694
rect 50380 2692 50436 2694
rect 50460 2692 50516 2694
rect 50540 2692 50596 2694
rect 50986 6704 51042 6760
rect 50986 5752 51042 5808
rect 50894 5652 50896 5672
rect 50896 5652 50948 5672
rect 50948 5652 50950 5672
rect 50894 5616 50950 5652
rect 51170 5208 51226 5264
rect 50894 5072 50950 5128
rect 51078 5072 51134 5128
rect 50894 4428 50896 4448
rect 50896 4428 50948 4448
rect 50948 4428 50950 4448
rect 50894 4392 50950 4428
rect 51078 4428 51080 4448
rect 51080 4428 51132 4448
rect 51132 4428 51134 4448
rect 51078 4392 51134 4428
rect 53930 12280 53986 12336
rect 55218 12552 55274 12608
rect 55494 14592 55550 14648
rect 55218 10956 55220 10976
rect 55220 10956 55272 10976
rect 55272 10956 55274 10976
rect 55218 10920 55274 10956
rect 52826 5616 52882 5672
rect 52458 3984 52514 4040
rect 52734 4020 52736 4040
rect 52736 4020 52788 4040
rect 52788 4020 52790 4040
rect 52734 3984 52790 4020
rect 55218 9444 55274 9480
rect 55218 9424 55220 9444
rect 55220 9424 55272 9444
rect 55272 9424 55274 9444
rect 55218 7928 55274 7984
rect 56506 21256 56562 21312
rect 56046 14184 56102 14240
rect 56138 13676 56140 13696
rect 56140 13676 56192 13696
rect 56192 13676 56194 13696
rect 56138 13640 56194 13676
rect 57426 30096 57482 30152
rect 57058 28620 57114 28656
rect 58162 33768 58218 33824
rect 58162 32136 58218 32192
rect 58162 30660 58218 30696
rect 58162 30640 58164 30660
rect 58164 30640 58216 30660
rect 58216 30640 58218 30660
rect 58162 29028 58218 29064
rect 58162 29008 58164 29028
rect 58164 29008 58216 29028
rect 58216 29008 58218 29028
rect 57058 28600 57060 28620
rect 57060 28600 57112 28620
rect 57112 28600 57114 28620
rect 57058 27548 57060 27568
rect 57060 27548 57112 27568
rect 57112 27548 57114 27568
rect 57058 27512 57114 27548
rect 57334 26968 57390 27024
rect 57886 26016 57942 26072
rect 57702 25880 57758 25936
rect 58162 25472 58218 25528
rect 56966 23840 57022 23896
rect 57150 23180 57206 23216
rect 57150 23160 57152 23180
rect 57152 23160 57204 23180
rect 57204 23160 57206 23180
rect 57058 19216 57114 19272
rect 56966 18944 57022 19000
rect 58162 24384 58218 24440
rect 57886 22888 57942 22944
rect 57426 22344 57482 22400
rect 57518 20848 57574 20904
rect 58162 19760 58218 19816
rect 56782 18400 56838 18456
rect 58162 18264 58218 18320
rect 57058 17720 57114 17776
rect 57150 17040 57206 17096
rect 58162 16632 58218 16688
rect 57426 16088 57482 16144
rect 57886 15136 57942 15192
rect 57058 13504 57114 13560
rect 57334 13096 57390 13152
rect 57150 11636 57152 11656
rect 57152 11636 57204 11656
rect 57204 11636 57206 11656
rect 57150 11600 57206 11636
rect 57058 9988 57114 10024
rect 57058 9968 57060 9988
rect 57060 9968 57112 9988
rect 57112 9968 57114 9988
rect 56598 8064 56654 8120
rect 55402 7656 55458 7712
rect 55310 6296 55366 6352
rect 57334 7828 57336 7848
rect 57336 7828 57388 7848
rect 57388 7828 57390 7848
rect 54390 5108 54392 5128
rect 54392 5108 54444 5128
rect 54444 5108 54446 5128
rect 54390 5072 54446 5108
rect 55218 4820 55274 4856
rect 55218 4800 55220 4820
rect 55220 4800 55272 4820
rect 55272 4800 55274 4820
rect 55218 3984 55274 4040
rect 54206 3884 54208 3904
rect 54208 3884 54260 3904
rect 54260 3884 54262 3904
rect 54206 3848 54262 3884
rect 55218 3168 55274 3224
rect 54850 2896 54906 2952
rect 55494 3304 55550 3360
rect 55218 1672 55274 1728
rect 2962 448 3018 504
rect 55954 3984 56010 4040
rect 56046 3712 56102 3768
rect 55862 2916 55918 2952
rect 55862 2896 55864 2916
rect 55864 2896 55916 2916
rect 55916 2896 55918 2916
rect 56690 5480 56746 5536
rect 56690 4140 56746 4176
rect 56690 4120 56692 4140
rect 56692 4120 56744 4140
rect 56744 4120 56746 4140
rect 56782 3848 56838 3904
rect 57334 7792 57390 7828
rect 57150 6840 57206 6896
rect 57886 12008 57942 12064
rect 58162 11464 58218 11520
rect 58162 10532 58218 10568
rect 58162 10512 58164 10532
rect 58164 10512 58216 10532
rect 58216 10512 58218 10532
rect 58162 8880 58218 8936
rect 58162 8356 58218 8392
rect 58162 8336 58164 8356
rect 58164 8336 58216 8356
rect 58216 8336 58218 8356
rect 58162 7404 58218 7440
rect 58162 7384 58164 7404
rect 58164 7384 58216 7404
rect 58216 7384 58218 7404
rect 56966 5364 57022 5400
rect 56966 5344 56968 5364
rect 56968 5344 57020 5364
rect 57020 5344 57022 5364
rect 57242 4564 57244 4584
rect 57244 4564 57296 4584
rect 57296 4564 57298 4584
rect 57242 4528 57298 4564
rect 56966 4256 57022 4312
rect 55770 2216 55826 2272
rect 55218 176 55274 232
rect 57058 3052 57114 3088
rect 57058 3032 57060 3052
rect 57060 3032 57112 3052
rect 57112 3032 57114 3052
rect 58162 5772 58218 5808
rect 58162 5752 58164 5772
rect 58164 5752 58216 5772
rect 58216 5752 58218 5772
rect 58162 2760 58218 2816
rect 57886 1128 57942 1184
rect 56414 584 56470 640
<< metal3 >>
rect 56501 59666 56567 59669
rect 59200 59666 60000 59696
rect 56501 59664 60000 59666
rect 56501 59608 56506 59664
rect 56562 59608 60000 59664
rect 56501 59606 60000 59608
rect 56501 59603 56567 59606
rect 59200 59576 60000 59606
rect 0 59530 800 59560
rect 2773 59530 2839 59533
rect 0 59528 2839 59530
rect 0 59472 2778 59528
rect 2834 59472 2839 59528
rect 0 59470 2839 59472
rect 0 59440 800 59470
rect 2773 59467 2839 59470
rect 56317 59122 56383 59125
rect 59200 59122 60000 59152
rect 56317 59120 60000 59122
rect 56317 59064 56322 59120
rect 56378 59064 60000 59120
rect 56317 59062 60000 59064
rect 56317 59059 56383 59062
rect 59200 59032 60000 59062
rect 0 58578 800 58608
rect 2037 58578 2103 58581
rect 0 58576 2103 58578
rect 0 58520 2042 58576
rect 2098 58520 2103 58576
rect 0 58518 2103 58520
rect 0 58488 800 58518
rect 2037 58515 2103 58518
rect 55489 58578 55555 58581
rect 59200 58578 60000 58608
rect 55489 58576 60000 58578
rect 55489 58520 55494 58576
rect 55550 58520 60000 58576
rect 55489 58518 60000 58520
rect 55489 58515 55555 58518
rect 59200 58488 60000 58518
rect 55029 58442 55095 58445
rect 56317 58442 56383 58445
rect 55029 58440 56383 58442
rect 55029 58384 55034 58440
rect 55090 58384 56322 58440
rect 56378 58384 56383 58440
rect 55029 58382 56383 58384
rect 55029 58379 55095 58382
rect 56317 58379 56383 58382
rect 54937 58170 55003 58173
rect 56501 58170 56567 58173
rect 54937 58168 56567 58170
rect 54937 58112 54942 58168
rect 54998 58112 56506 58168
rect 56562 58112 56567 58168
rect 54937 58110 56567 58112
rect 54937 58107 55003 58110
rect 56501 58107 56567 58110
rect 56501 58034 56567 58037
rect 59200 58034 60000 58064
rect 56501 58032 60000 58034
rect 56501 57976 56506 58032
rect 56562 57976 60000 58032
rect 56501 57974 60000 57976
rect 56501 57971 56567 57974
rect 59200 57944 60000 57974
rect 4208 57696 4528 57697
rect 0 57626 800 57656
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 1393 57626 1459 57629
rect 0 57624 1459 57626
rect 0 57568 1398 57624
rect 1454 57568 1459 57624
rect 0 57566 1459 57568
rect 0 57536 800 57566
rect 1393 57563 1459 57566
rect 55581 57490 55647 57493
rect 59200 57490 60000 57520
rect 55581 57488 60000 57490
rect 55581 57432 55586 57488
rect 55642 57432 60000 57488
rect 55581 57430 60000 57432
rect 55581 57427 55647 57430
rect 59200 57400 60000 57430
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 50288 57152 50608 57153
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 57087 50608 57088
rect 58157 57082 58223 57085
rect 59200 57082 60000 57112
rect 58157 57080 60000 57082
rect 58157 57024 58162 57080
rect 58218 57024 60000 57080
rect 58157 57022 60000 57024
rect 58157 57019 58223 57022
rect 59200 56992 60000 57022
rect 0 56674 800 56704
rect 1393 56674 1459 56677
rect 0 56672 1459 56674
rect 0 56616 1398 56672
rect 1454 56616 1459 56672
rect 0 56614 1459 56616
rect 0 56584 800 56614
rect 1393 56611 1459 56614
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 57053 56538 57119 56541
rect 59200 56538 60000 56568
rect 57053 56536 60000 56538
rect 57053 56480 57058 56536
rect 57114 56480 60000 56536
rect 57053 56478 60000 56480
rect 57053 56475 57119 56478
rect 59200 56448 60000 56478
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect 50288 56064 50608 56065
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 55999 50608 56000
rect 55673 55994 55739 55997
rect 59200 55994 60000 56024
rect 55673 55992 60000 55994
rect 55673 55936 55678 55992
rect 55734 55936 60000 55992
rect 55673 55934 60000 55936
rect 55673 55931 55739 55934
rect 59200 55904 60000 55934
rect 0 55722 800 55752
rect 1393 55722 1459 55725
rect 0 55720 1459 55722
rect 0 55664 1398 55720
rect 1454 55664 1459 55720
rect 0 55662 1459 55664
rect 0 55632 800 55662
rect 1393 55659 1459 55662
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 58157 55450 58223 55453
rect 59200 55450 60000 55480
rect 58157 55448 60000 55450
rect 58157 55392 58162 55448
rect 58218 55392 60000 55448
rect 58157 55390 60000 55392
rect 58157 55387 58223 55390
rect 59200 55360 60000 55390
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 50288 54976 50608 54977
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 54911 50608 54912
rect 57053 54906 57119 54909
rect 59200 54906 60000 54936
rect 57053 54904 60000 54906
rect 57053 54848 57058 54904
rect 57114 54848 60000 54904
rect 57053 54846 60000 54848
rect 57053 54843 57119 54846
rect 59200 54816 60000 54846
rect 0 54770 800 54800
rect 1393 54770 1459 54773
rect 0 54768 1459 54770
rect 0 54712 1398 54768
rect 1454 54712 1459 54768
rect 0 54710 1459 54712
rect 0 54680 800 54710
rect 1393 54707 1459 54710
rect 55489 54498 55555 54501
rect 59200 54498 60000 54528
rect 55489 54496 60000 54498
rect 55489 54440 55494 54496
rect 55550 54440 60000 54496
rect 55489 54438 60000 54440
rect 55489 54435 55555 54438
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 59200 54408 60000 54438
rect 34928 54367 35248 54368
rect 58157 53954 58223 53957
rect 59200 53954 60000 53984
rect 58157 53952 60000 53954
rect 58157 53896 58162 53952
rect 58218 53896 60000 53952
rect 58157 53894 60000 53896
rect 58157 53891 58223 53894
rect 19568 53888 19888 53889
rect 0 53818 800 53848
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 50288 53888 50608 53889
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 59200 53864 60000 53894
rect 50288 53823 50608 53824
rect 1393 53818 1459 53821
rect 0 53816 1459 53818
rect 0 53760 1398 53816
rect 1454 53760 1459 53816
rect 0 53758 1459 53760
rect 0 53728 800 53758
rect 1393 53755 1459 53758
rect 56961 53410 57027 53413
rect 59200 53410 60000 53440
rect 56961 53408 60000 53410
rect 56961 53352 56966 53408
rect 57022 53352 60000 53408
rect 56961 53350 60000 53352
rect 56961 53347 57027 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 59200 53320 60000 53350
rect 34928 53279 35248 53280
rect 0 52866 800 52896
rect 1393 52866 1459 52869
rect 0 52864 1459 52866
rect 0 52808 1398 52864
rect 1454 52808 1459 52864
rect 0 52806 1459 52808
rect 0 52776 800 52806
rect 1393 52803 1459 52806
rect 55581 52866 55647 52869
rect 59200 52866 60000 52896
rect 55581 52864 60000 52866
rect 55581 52808 55586 52864
rect 55642 52808 60000 52864
rect 55581 52806 60000 52808
rect 55581 52803 55647 52806
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 50288 52800 50608 52801
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 59200 52776 60000 52806
rect 50288 52735 50608 52736
rect 57881 52322 57947 52325
rect 59200 52322 60000 52352
rect 57881 52320 60000 52322
rect 57881 52264 57886 52320
rect 57942 52264 60000 52320
rect 57881 52262 60000 52264
rect 57881 52259 57947 52262
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 59200 52232 60000 52262
rect 34928 52191 35248 52192
rect 0 51914 800 51944
rect 1393 51914 1459 51917
rect 0 51912 1459 51914
rect 0 51856 1398 51912
rect 1454 51856 1459 51912
rect 0 51854 1459 51856
rect 0 51824 800 51854
rect 1393 51851 1459 51854
rect 57053 51914 57119 51917
rect 59200 51914 60000 51944
rect 57053 51912 60000 51914
rect 57053 51856 57058 51912
rect 57114 51856 60000 51912
rect 57053 51854 60000 51856
rect 57053 51851 57119 51854
rect 59200 51824 60000 51854
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 50288 51712 50608 51713
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 51647 50608 51648
rect 55489 51370 55555 51373
rect 59200 51370 60000 51400
rect 55489 51368 60000 51370
rect 55489 51312 55494 51368
rect 55550 51312 60000 51368
rect 55489 51310 60000 51312
rect 55489 51307 55555 51310
rect 59200 51280 60000 51310
rect 4208 51168 4528 51169
rect 0 51098 800 51128
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 51103 35248 51104
rect 1393 51098 1459 51101
rect 0 51096 1459 51098
rect 0 51040 1398 51096
rect 1454 51040 1459 51096
rect 0 51038 1459 51040
rect 0 51008 800 51038
rect 1393 51035 1459 51038
rect 58157 50826 58223 50829
rect 59200 50826 60000 50856
rect 58157 50824 60000 50826
rect 58157 50768 58162 50824
rect 58218 50768 60000 50824
rect 58157 50766 60000 50768
rect 58157 50763 58223 50766
rect 59200 50736 60000 50766
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 50559 19888 50560
rect 50288 50624 50608 50625
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 50559 50608 50560
rect 57053 50282 57119 50285
rect 59200 50282 60000 50312
rect 57053 50280 60000 50282
rect 57053 50224 57058 50280
rect 57114 50224 60000 50280
rect 57053 50222 60000 50224
rect 57053 50219 57119 50222
rect 59200 50192 60000 50222
rect 0 50146 800 50176
rect 1393 50146 1459 50149
rect 0 50144 1459 50146
rect 0 50088 1398 50144
rect 1454 50088 1459 50144
rect 0 50086 1459 50088
rect 0 50056 800 50086
rect 1393 50083 1459 50086
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 55213 49738 55279 49741
rect 59200 49738 60000 49768
rect 55213 49736 60000 49738
rect 55213 49680 55218 49736
rect 55274 49680 60000 49736
rect 55213 49678 60000 49680
rect 55213 49675 55279 49678
rect 59200 49648 60000 49678
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 50288 49536 50608 49537
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 49471 50608 49472
rect 58157 49330 58223 49333
rect 59200 49330 60000 49360
rect 58157 49328 60000 49330
rect 58157 49272 58162 49328
rect 58218 49272 60000 49328
rect 58157 49270 60000 49272
rect 58157 49267 58223 49270
rect 59200 49240 60000 49270
rect 0 49194 800 49224
rect 1393 49194 1459 49197
rect 0 49192 1459 49194
rect 0 49136 1398 49192
rect 1454 49136 1459 49192
rect 0 49134 1459 49136
rect 0 49104 800 49134
rect 1393 49131 1459 49134
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 57053 48786 57119 48789
rect 59200 48786 60000 48816
rect 57053 48784 60000 48786
rect 57053 48728 57058 48784
rect 57114 48728 60000 48784
rect 57053 48726 60000 48728
rect 57053 48723 57119 48726
rect 59200 48696 60000 48726
rect 19568 48448 19888 48449
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 50288 48448 50608 48449
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 48383 50608 48384
rect 0 48242 800 48272
rect 1393 48242 1459 48245
rect 0 48240 1459 48242
rect 0 48184 1398 48240
rect 1454 48184 1459 48240
rect 0 48182 1459 48184
rect 0 48152 800 48182
rect 1393 48179 1459 48182
rect 55489 48242 55555 48245
rect 59200 48242 60000 48272
rect 55489 48240 60000 48242
rect 55489 48184 55494 48240
rect 55550 48184 60000 48240
rect 55489 48182 60000 48184
rect 55489 48179 55555 48182
rect 59200 48152 60000 48182
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 57053 47698 57119 47701
rect 59200 47698 60000 47728
rect 57053 47696 60000 47698
rect 57053 47640 57058 47696
rect 57114 47640 60000 47696
rect 57053 47638 60000 47640
rect 57053 47635 57119 47638
rect 59200 47608 60000 47638
rect 19568 47360 19888 47361
rect 0 47290 800 47320
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 50288 47360 50608 47361
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 47295 50608 47296
rect 1393 47290 1459 47293
rect 0 47288 1459 47290
rect 0 47232 1398 47288
rect 1454 47232 1459 47288
rect 0 47230 1459 47232
rect 0 47200 800 47230
rect 1393 47227 1459 47230
rect 57421 47154 57487 47157
rect 59200 47154 60000 47184
rect 57421 47152 60000 47154
rect 57421 47096 57426 47152
rect 57482 47096 60000 47152
rect 57421 47094 60000 47096
rect 57421 47091 57487 47094
rect 59200 47064 60000 47094
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 55213 46746 55279 46749
rect 59200 46746 60000 46776
rect 55213 46744 60000 46746
rect 55213 46688 55218 46744
rect 55274 46688 60000 46744
rect 55213 46686 60000 46688
rect 55213 46683 55279 46686
rect 59200 46656 60000 46686
rect 0 46338 800 46368
rect 1393 46338 1459 46341
rect 0 46336 1459 46338
rect 0 46280 1398 46336
rect 1454 46280 1459 46336
rect 0 46278 1459 46280
rect 0 46248 800 46278
rect 1393 46275 1459 46278
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 50288 46272 50608 46273
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 46207 50608 46208
rect 57881 46202 57947 46205
rect 59200 46202 60000 46232
rect 57881 46200 60000 46202
rect 57881 46144 57886 46200
rect 57942 46144 60000 46200
rect 57881 46142 60000 46144
rect 57881 46139 57947 46142
rect 59200 46112 60000 46142
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 57053 45658 57119 45661
rect 59200 45658 60000 45688
rect 57053 45656 60000 45658
rect 57053 45600 57058 45656
rect 57114 45600 60000 45656
rect 57053 45598 60000 45600
rect 57053 45595 57119 45598
rect 59200 45568 60000 45598
rect 0 45386 800 45416
rect 1393 45386 1459 45389
rect 0 45384 1459 45386
rect 0 45328 1398 45384
rect 1454 45328 1459 45384
rect 0 45326 1459 45328
rect 0 45296 800 45326
rect 1393 45323 1459 45326
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 50288 45184 50608 45185
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 45119 50608 45120
rect 55029 45114 55095 45117
rect 59200 45114 60000 45144
rect 55029 45112 60000 45114
rect 55029 45056 55034 45112
rect 55090 45056 60000 45112
rect 55029 45054 60000 45056
rect 55029 45051 55095 45054
rect 59200 45024 60000 45054
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 58157 44570 58223 44573
rect 59200 44570 60000 44600
rect 58157 44568 60000 44570
rect 58157 44512 58162 44568
rect 58218 44512 60000 44568
rect 58157 44510 60000 44512
rect 58157 44507 58223 44510
rect 59200 44480 60000 44510
rect 0 44434 800 44464
rect 1393 44434 1459 44437
rect 0 44432 1459 44434
rect 0 44376 1398 44432
rect 1454 44376 1459 44432
rect 0 44374 1459 44376
rect 0 44344 800 44374
rect 1393 44371 1459 44374
rect 57053 44162 57119 44165
rect 59200 44162 60000 44192
rect 57053 44160 60000 44162
rect 57053 44104 57058 44160
rect 57114 44104 60000 44160
rect 57053 44102 60000 44104
rect 57053 44099 57119 44102
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 59200 44072 60000 44102
rect 50288 44031 50608 44032
rect 54753 43618 54819 43621
rect 59200 43618 60000 43648
rect 54753 43616 60000 43618
rect 54753 43560 54758 43616
rect 54814 43560 60000 43616
rect 54753 43558 60000 43560
rect 54753 43555 54819 43558
rect 4208 43552 4528 43553
rect 0 43482 800 43512
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 59200 43528 60000 43558
rect 34928 43487 35248 43488
rect 1393 43482 1459 43485
rect 0 43480 1459 43482
rect 0 43424 1398 43480
rect 1454 43424 1459 43480
rect 0 43422 1459 43424
rect 0 43392 800 43422
rect 1393 43419 1459 43422
rect 58157 43074 58223 43077
rect 59200 43074 60000 43104
rect 58157 43072 60000 43074
rect 58157 43016 58162 43072
rect 58218 43016 60000 43072
rect 58157 43014 60000 43016
rect 58157 43011 58223 43014
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 59200 42984 60000 43014
rect 50288 42943 50608 42944
rect 0 42666 800 42696
rect 1393 42666 1459 42669
rect 0 42664 1459 42666
rect 0 42608 1398 42664
rect 1454 42608 1459 42664
rect 0 42606 1459 42608
rect 0 42576 800 42606
rect 1393 42603 1459 42606
rect 56961 42530 57027 42533
rect 59200 42530 60000 42560
rect 56961 42528 60000 42530
rect 56961 42472 56966 42528
rect 57022 42472 60000 42528
rect 56961 42470 60000 42472
rect 56961 42467 57027 42470
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 59200 42440 60000 42470
rect 34928 42399 35248 42400
rect 50429 42258 50495 42261
rect 52177 42258 52243 42261
rect 50429 42256 52243 42258
rect 50429 42200 50434 42256
rect 50490 42200 52182 42256
rect 52238 42200 52243 42256
rect 50429 42198 52243 42200
rect 50429 42195 50495 42198
rect 52177 42195 52243 42198
rect 49417 42122 49483 42125
rect 49417 42120 57990 42122
rect 49417 42064 49422 42120
rect 49478 42064 57990 42120
rect 49417 42062 57990 42064
rect 49417 42059 49483 42062
rect 57930 41986 57990 42062
rect 59200 41986 60000 42016
rect 57930 41926 60000 41986
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 59200 41896 60000 41926
rect 50288 41855 50608 41856
rect 0 41714 800 41744
rect 1393 41714 1459 41717
rect 0 41712 1459 41714
rect 0 41656 1398 41712
rect 1454 41656 1459 41712
rect 0 41654 1459 41656
rect 0 41624 800 41654
rect 1393 41651 1459 41654
rect 58157 41578 58223 41581
rect 59200 41578 60000 41608
rect 58157 41576 60000 41578
rect 58157 41520 58162 41576
rect 58218 41520 60000 41576
rect 58157 41518 60000 41520
rect 58157 41515 58223 41518
rect 59200 41488 60000 41518
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 57421 41034 57487 41037
rect 59200 41034 60000 41064
rect 57421 41032 60000 41034
rect 57421 40976 57426 41032
rect 57482 40976 60000 41032
rect 57421 40974 60000 40976
rect 57421 40971 57487 40974
rect 59200 40944 60000 40974
rect 19568 40832 19888 40833
rect 0 40762 800 40792
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 1393 40762 1459 40765
rect 0 40760 1459 40762
rect 0 40704 1398 40760
rect 1454 40704 1459 40760
rect 0 40702 1459 40704
rect 0 40672 800 40702
rect 1393 40699 1459 40702
rect 55213 40490 55279 40493
rect 59200 40490 60000 40520
rect 55213 40488 60000 40490
rect 55213 40432 55218 40488
rect 55274 40432 60000 40488
rect 55213 40430 60000 40432
rect 55213 40427 55279 40430
rect 59200 40400 60000 40430
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 57881 39946 57947 39949
rect 59200 39946 60000 39976
rect 57881 39944 60000 39946
rect 57881 39888 57886 39944
rect 57942 39888 60000 39944
rect 57881 39886 60000 39888
rect 57881 39883 57947 39886
rect 59200 39856 60000 39886
rect 0 39810 800 39840
rect 1393 39810 1459 39813
rect 0 39808 1459 39810
rect 0 39752 1398 39808
rect 1454 39752 1459 39808
rect 0 39750 1459 39752
rect 0 39720 800 39750
rect 1393 39747 1459 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 56961 39402 57027 39405
rect 59200 39402 60000 39432
rect 56961 39400 60000 39402
rect 56961 39344 56966 39400
rect 57022 39344 60000 39400
rect 56961 39342 60000 39344
rect 56961 39339 57027 39342
rect 59200 39312 60000 39342
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 52545 38994 52611 38997
rect 53281 38994 53347 38997
rect 52545 38992 53347 38994
rect 52545 38936 52550 38992
rect 52606 38936 53286 38992
rect 53342 38936 53347 38992
rect 52545 38934 53347 38936
rect 52545 38931 52611 38934
rect 53281 38931 53347 38934
rect 55213 38994 55279 38997
rect 59200 38994 60000 39024
rect 55213 38992 60000 38994
rect 55213 38936 55218 38992
rect 55274 38936 60000 38992
rect 55213 38934 60000 38936
rect 55213 38931 55279 38934
rect 59200 38904 60000 38934
rect 0 38858 800 38888
rect 1393 38858 1459 38861
rect 0 38856 1459 38858
rect 0 38800 1398 38856
rect 1454 38800 1459 38856
rect 0 38798 1459 38800
rect 0 38768 800 38798
rect 1393 38795 1459 38798
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 50705 38586 50771 38589
rect 54201 38586 54267 38589
rect 50705 38584 54267 38586
rect 50705 38528 50710 38584
rect 50766 38528 54206 38584
rect 54262 38528 54267 38584
rect 50705 38526 54267 38528
rect 50705 38523 50771 38526
rect 54201 38523 54267 38526
rect 52453 38450 52519 38453
rect 53373 38450 53439 38453
rect 52453 38448 53439 38450
rect 52453 38392 52458 38448
rect 52514 38392 53378 38448
rect 53434 38392 53439 38448
rect 52453 38390 53439 38392
rect 52453 38387 52519 38390
rect 53373 38387 53439 38390
rect 58157 38450 58223 38453
rect 59200 38450 60000 38480
rect 58157 38448 60000 38450
rect 58157 38392 58162 38448
rect 58218 38392 60000 38448
rect 58157 38390 60000 38392
rect 58157 38387 58223 38390
rect 59200 38360 60000 38390
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 0 37906 800 37936
rect 1393 37906 1459 37909
rect 0 37904 1459 37906
rect 0 37848 1398 37904
rect 1454 37848 1459 37904
rect 0 37846 1459 37848
rect 0 37816 800 37846
rect 1393 37843 1459 37846
rect 57881 37906 57947 37909
rect 59200 37906 60000 37936
rect 57881 37904 60000 37906
rect 57881 37848 57886 37904
rect 57942 37848 60000 37904
rect 57881 37846 60000 37848
rect 57881 37843 57947 37846
rect 59200 37816 60000 37846
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 55213 37362 55279 37365
rect 59200 37362 60000 37392
rect 55213 37360 60000 37362
rect 55213 37304 55218 37360
rect 55274 37304 60000 37360
rect 55213 37302 60000 37304
rect 55213 37299 55279 37302
rect 59200 37272 60000 37302
rect 49785 37226 49851 37229
rect 57053 37226 57119 37229
rect 49785 37224 57119 37226
rect 49785 37168 49790 37224
rect 49846 37168 57058 37224
rect 57114 37168 57119 37224
rect 49785 37166 57119 37168
rect 49785 37163 49851 37166
rect 57053 37163 57119 37166
rect 51901 37090 51967 37093
rect 52637 37090 52703 37093
rect 51901 37088 52703 37090
rect 51901 37032 51906 37088
rect 51962 37032 52642 37088
rect 52698 37032 52703 37088
rect 51901 37030 52703 37032
rect 51901 37027 51967 37030
rect 52637 37027 52703 37030
rect 4208 37024 4528 37025
rect 0 36954 800 36984
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 1393 36954 1459 36957
rect 0 36952 1459 36954
rect 0 36896 1398 36952
rect 1454 36896 1459 36952
rect 0 36894 1459 36896
rect 0 36864 800 36894
rect 1393 36891 1459 36894
rect 58157 36818 58223 36821
rect 59200 36818 60000 36848
rect 58157 36816 60000 36818
rect 58157 36760 58162 36816
rect 58218 36760 60000 36816
rect 58157 36758 60000 36760
rect 58157 36755 58223 36758
rect 59200 36728 60000 36758
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 56961 36410 57027 36413
rect 59200 36410 60000 36440
rect 56961 36408 60000 36410
rect 56961 36352 56966 36408
rect 57022 36352 60000 36408
rect 56961 36350 60000 36352
rect 56961 36347 57027 36350
rect 59200 36320 60000 36350
rect 0 36002 800 36032
rect 1393 36002 1459 36005
rect 0 36000 1459 36002
rect 0 35944 1398 36000
rect 1454 35944 1459 36000
rect 0 35942 1459 35944
rect 0 35912 800 35942
rect 1393 35939 1459 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 55213 35866 55279 35869
rect 59200 35866 60000 35896
rect 55213 35864 60000 35866
rect 55213 35808 55218 35864
rect 55274 35808 60000 35864
rect 55213 35806 60000 35808
rect 55213 35803 55279 35806
rect 59200 35776 60000 35806
rect 54385 35458 54451 35461
rect 56593 35458 56659 35461
rect 54385 35456 56659 35458
rect 54385 35400 54390 35456
rect 54446 35400 56598 35456
rect 56654 35400 56659 35456
rect 54385 35398 56659 35400
rect 54385 35395 54451 35398
rect 56593 35395 56659 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 56961 35322 57027 35325
rect 59200 35322 60000 35352
rect 56961 35320 60000 35322
rect 56961 35264 56966 35320
rect 57022 35264 60000 35320
rect 56961 35262 60000 35264
rect 56961 35259 57027 35262
rect 59200 35232 60000 35262
rect 49877 35186 49943 35189
rect 54937 35186 55003 35189
rect 49877 35184 55003 35186
rect 49877 35128 49882 35184
rect 49938 35128 54942 35184
rect 54998 35128 55003 35184
rect 49877 35126 55003 35128
rect 49877 35123 49943 35126
rect 54937 35123 55003 35126
rect 0 35050 800 35080
rect 1393 35050 1459 35053
rect 0 35048 1459 35050
rect 0 34992 1398 35048
rect 1454 34992 1459 35048
rect 0 34990 1459 34992
rect 0 34960 800 34990
rect 1393 34987 1459 34990
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 56409 34778 56475 34781
rect 59200 34778 60000 34808
rect 56409 34776 60000 34778
rect 56409 34720 56414 34776
rect 56470 34720 60000 34776
rect 56409 34718 60000 34720
rect 56409 34715 56475 34718
rect 59200 34688 60000 34718
rect 50337 34642 50403 34645
rect 57053 34642 57119 34645
rect 50337 34640 57119 34642
rect 50337 34584 50342 34640
rect 50398 34584 57058 34640
rect 57114 34584 57119 34640
rect 50337 34582 57119 34584
rect 50337 34579 50403 34582
rect 57053 34579 57119 34582
rect 50613 34506 50679 34509
rect 56869 34506 56935 34509
rect 50613 34504 56935 34506
rect 50613 34448 50618 34504
rect 50674 34448 56874 34504
rect 56930 34448 56935 34504
rect 50613 34446 56935 34448
rect 50613 34443 50679 34446
rect 56869 34443 56935 34446
rect 54569 34370 54635 34373
rect 55489 34370 55555 34373
rect 54569 34368 55555 34370
rect 54569 34312 54574 34368
rect 54630 34312 55494 34368
rect 55550 34312 55555 34368
rect 54569 34310 55555 34312
rect 54569 34307 54635 34310
rect 55489 34307 55555 34310
rect 19568 34304 19888 34305
rect 0 34234 800 34264
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 1393 34234 1459 34237
rect 0 34232 1459 34234
rect 0 34176 1398 34232
rect 1454 34176 1459 34232
rect 0 34174 1459 34176
rect 0 34144 800 34174
rect 1393 34171 1459 34174
rect 55213 34234 55279 34237
rect 59200 34234 60000 34264
rect 55213 34232 60000 34234
rect 55213 34176 55218 34232
rect 55274 34176 60000 34232
rect 55213 34174 60000 34176
rect 55213 34171 55279 34174
rect 59200 34144 60000 34174
rect 50797 34098 50863 34101
rect 56777 34098 56843 34101
rect 50797 34096 56843 34098
rect 50797 34040 50802 34096
rect 50858 34040 56782 34096
rect 56838 34040 56843 34096
rect 50797 34038 56843 34040
rect 50797 34035 50863 34038
rect 56777 34035 56843 34038
rect 53281 33826 53347 33829
rect 54753 33826 54819 33829
rect 55397 33826 55463 33829
rect 53281 33824 55463 33826
rect 53281 33768 53286 33824
rect 53342 33768 54758 33824
rect 54814 33768 55402 33824
rect 55458 33768 55463 33824
rect 53281 33766 55463 33768
rect 53281 33763 53347 33766
rect 54753 33763 54819 33766
rect 55397 33763 55463 33766
rect 58157 33826 58223 33829
rect 59200 33826 60000 33856
rect 58157 33824 60000 33826
rect 58157 33768 58162 33824
rect 58218 33768 60000 33824
rect 58157 33766 60000 33768
rect 58157 33763 58223 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 59200 33736 60000 33766
rect 34928 33695 35248 33696
rect 52545 33554 52611 33557
rect 54661 33554 54727 33557
rect 55581 33554 55647 33557
rect 52545 33552 55647 33554
rect 52545 33496 52550 33552
rect 52606 33496 54666 33552
rect 54722 33496 55586 33552
rect 55642 33496 55647 33552
rect 52545 33494 55647 33496
rect 52545 33491 52611 33494
rect 54661 33491 54727 33494
rect 55581 33491 55647 33494
rect 0 33282 800 33312
rect 1393 33282 1459 33285
rect 0 33280 1459 33282
rect 0 33224 1398 33280
rect 1454 33224 1459 33280
rect 0 33222 1459 33224
rect 0 33192 800 33222
rect 1393 33219 1459 33222
rect 57329 33282 57395 33285
rect 59200 33282 60000 33312
rect 57329 33280 60000 33282
rect 57329 33224 57334 33280
rect 57390 33224 60000 33280
rect 57329 33222 60000 33224
rect 57329 33219 57395 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 59200 33192 60000 33222
rect 50288 33151 50608 33152
rect 49693 32738 49759 32741
rect 59200 32738 60000 32768
rect 49693 32736 60000 32738
rect 49693 32680 49698 32736
rect 49754 32680 60000 32736
rect 49693 32678 60000 32680
rect 49693 32675 49759 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 59200 32648 60000 32678
rect 34928 32607 35248 32608
rect 0 32330 800 32360
rect 1393 32330 1459 32333
rect 0 32328 1459 32330
rect 0 32272 1398 32328
rect 1454 32272 1459 32328
rect 0 32270 1459 32272
rect 0 32240 800 32270
rect 1393 32267 1459 32270
rect 58157 32194 58223 32197
rect 59200 32194 60000 32224
rect 58157 32192 60000 32194
rect 58157 32136 58162 32192
rect 58218 32136 60000 32192
rect 58157 32134 60000 32136
rect 58157 32131 58223 32134
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 59200 32104 60000 32134
rect 50288 32063 50608 32064
rect 51809 31922 51875 31925
rect 53833 31922 53899 31925
rect 51809 31920 53899 31922
rect 51809 31864 51814 31920
rect 51870 31864 53838 31920
rect 53894 31864 53899 31920
rect 51809 31862 53899 31864
rect 51809 31859 51875 31862
rect 53833 31859 53899 31862
rect 57421 31650 57487 31653
rect 59200 31650 60000 31680
rect 57421 31648 60000 31650
rect 57421 31592 57426 31648
rect 57482 31592 60000 31648
rect 57421 31590 60000 31592
rect 57421 31587 57487 31590
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 59200 31560 60000 31590
rect 34928 31519 35248 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 55213 31242 55279 31245
rect 59200 31242 60000 31272
rect 55213 31240 60000 31242
rect 55213 31184 55218 31240
rect 55274 31184 60000 31240
rect 55213 31182 60000 31184
rect 55213 31179 55279 31182
rect 59200 31152 60000 31182
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 50705 30970 50771 30973
rect 57421 30970 57487 30973
rect 50705 30968 57487 30970
rect 50705 30912 50710 30968
rect 50766 30912 57426 30968
rect 57482 30912 57487 30968
rect 50705 30910 57487 30912
rect 50705 30907 50771 30910
rect 57421 30907 57487 30910
rect 50521 30834 50587 30837
rect 53649 30834 53715 30837
rect 50521 30832 53715 30834
rect 50521 30776 50526 30832
rect 50582 30776 53654 30832
rect 53710 30776 53715 30832
rect 50521 30774 53715 30776
rect 50521 30771 50587 30774
rect 53649 30771 53715 30774
rect 53833 30834 53899 30837
rect 54753 30834 54819 30837
rect 53833 30832 54819 30834
rect 53833 30776 53838 30832
rect 53894 30776 54758 30832
rect 54814 30776 54819 30832
rect 53833 30774 54819 30776
rect 53833 30771 53899 30774
rect 54753 30771 54819 30774
rect 58157 30698 58223 30701
rect 59200 30698 60000 30728
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30608 60000 30638
rect 4208 30496 4528 30497
rect 0 30426 800 30456
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 1393 30426 1459 30429
rect 0 30424 1459 30426
rect 0 30368 1398 30424
rect 1454 30368 1459 30424
rect 0 30366 1459 30368
rect 0 30336 800 30366
rect 1393 30363 1459 30366
rect 57421 30154 57487 30157
rect 59200 30154 60000 30184
rect 57421 30152 60000 30154
rect 57421 30096 57426 30152
rect 57482 30096 60000 30152
rect 57421 30094 60000 30096
rect 57421 30091 57487 30094
rect 59200 30064 60000 30094
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 55489 29610 55555 29613
rect 59200 29610 60000 29640
rect 55489 29608 60000 29610
rect 55489 29552 55494 29608
rect 55550 29552 60000 29608
rect 55489 29550 60000 29552
rect 55489 29547 55555 29550
rect 59200 29520 60000 29550
rect 0 29474 800 29504
rect 1945 29474 2011 29477
rect 0 29472 2011 29474
rect 0 29416 1950 29472
rect 2006 29416 2011 29472
rect 0 29414 2011 29416
rect 0 29384 800 29414
rect 1945 29411 2011 29414
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 49509 29202 49575 29205
rect 55949 29202 56015 29205
rect 49509 29200 56015 29202
rect 49509 29144 49514 29200
rect 49570 29144 55954 29200
rect 56010 29144 56015 29200
rect 49509 29142 56015 29144
rect 49509 29139 49575 29142
rect 55949 29139 56015 29142
rect 58157 29066 58223 29069
rect 59200 29066 60000 29096
rect 58157 29064 60000 29066
rect 58157 29008 58162 29064
rect 58218 29008 60000 29064
rect 58157 29006 60000 29008
rect 58157 29003 58223 29006
rect 59200 28976 60000 29006
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 50288 28864 50608 28865
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 28799 50608 28800
rect 50705 28658 50771 28661
rect 52177 28658 52243 28661
rect 50705 28656 52243 28658
rect 50705 28600 50710 28656
rect 50766 28600 52182 28656
rect 52238 28600 52243 28656
rect 50705 28598 52243 28600
rect 50705 28595 50771 28598
rect 52177 28595 52243 28598
rect 57053 28658 57119 28661
rect 59200 28658 60000 28688
rect 57053 28656 60000 28658
rect 57053 28600 57058 28656
rect 57114 28600 60000 28656
rect 57053 28598 60000 28600
rect 57053 28595 57119 28598
rect 59200 28568 60000 28598
rect 0 28522 800 28552
rect 1393 28522 1459 28525
rect 0 28520 1459 28522
rect 0 28464 1398 28520
rect 1454 28464 1459 28520
rect 0 28462 1459 28464
rect 0 28432 800 28462
rect 1393 28459 1459 28462
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 55305 28114 55371 28117
rect 59200 28114 60000 28144
rect 55305 28112 60000 28114
rect 55305 28056 55310 28112
rect 55366 28056 60000 28112
rect 55305 28054 60000 28056
rect 55305 28051 55371 28054
rect 59200 28024 60000 28054
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 50288 27776 50608 27777
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 27711 50608 27712
rect 0 27570 800 27600
rect 1945 27570 2011 27573
rect 0 27568 2011 27570
rect 0 27512 1950 27568
rect 2006 27512 2011 27568
rect 0 27510 2011 27512
rect 0 27480 800 27510
rect 1945 27507 2011 27510
rect 50245 27570 50311 27573
rect 54201 27570 54267 27573
rect 50245 27568 54267 27570
rect 50245 27512 50250 27568
rect 50306 27512 54206 27568
rect 54262 27512 54267 27568
rect 50245 27510 54267 27512
rect 50245 27507 50311 27510
rect 54201 27507 54267 27510
rect 57053 27570 57119 27573
rect 59200 27570 60000 27600
rect 57053 27568 60000 27570
rect 57053 27512 57058 27568
rect 57114 27512 60000 27568
rect 57053 27510 60000 27512
rect 57053 27507 57119 27510
rect 59200 27480 60000 27510
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 57329 27026 57395 27029
rect 59200 27026 60000 27056
rect 57329 27024 60000 27026
rect 57329 26968 57334 27024
rect 57390 26968 60000 27024
rect 57329 26966 60000 26968
rect 57329 26963 57395 26966
rect 59200 26936 60000 26966
rect 19568 26688 19888 26689
rect 0 26618 800 26648
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 50288 26688 50608 26689
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 26623 50608 26624
rect 1945 26618 2011 26621
rect 0 26616 2011 26618
rect 0 26560 1950 26616
rect 2006 26560 2011 26616
rect 0 26558 2011 26560
rect 0 26528 800 26558
rect 1945 26555 2011 26558
rect 48405 26482 48471 26485
rect 52913 26482 52979 26485
rect 48405 26480 52979 26482
rect 48405 26424 48410 26480
rect 48466 26424 52918 26480
rect 52974 26424 52979 26480
rect 48405 26422 52979 26424
rect 48405 26419 48471 26422
rect 52913 26419 52979 26422
rect 55489 26482 55555 26485
rect 59200 26482 60000 26512
rect 55489 26480 60000 26482
rect 55489 26424 55494 26480
rect 55550 26424 60000 26480
rect 55489 26422 60000 26424
rect 55489 26419 55555 26422
rect 59200 26392 60000 26422
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 57881 26074 57947 26077
rect 59200 26074 60000 26104
rect 57881 26072 60000 26074
rect 57881 26016 57886 26072
rect 57942 26016 60000 26072
rect 57881 26014 60000 26016
rect 57881 26011 57947 26014
rect 59200 25984 60000 26014
rect 51901 25938 51967 25941
rect 57697 25938 57763 25941
rect 51901 25936 57763 25938
rect 51901 25880 51906 25936
rect 51962 25880 57702 25936
rect 57758 25880 57763 25936
rect 51901 25878 57763 25880
rect 51901 25875 51967 25878
rect 57697 25875 57763 25878
rect 0 25802 800 25832
rect 2037 25802 2103 25805
rect 0 25800 2103 25802
rect 0 25744 2042 25800
rect 2098 25744 2103 25800
rect 0 25742 2103 25744
rect 0 25712 800 25742
rect 2037 25739 2103 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 50288 25600 50608 25601
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 25535 50608 25536
rect 58157 25530 58223 25533
rect 59200 25530 60000 25560
rect 58157 25528 60000 25530
rect 58157 25472 58162 25528
rect 58218 25472 60000 25528
rect 58157 25470 60000 25472
rect 58157 25467 58223 25470
rect 59200 25440 60000 25470
rect 49601 25394 49667 25397
rect 56685 25394 56751 25397
rect 49601 25392 56751 25394
rect 49601 25336 49606 25392
rect 49662 25336 56690 25392
rect 56746 25336 56751 25392
rect 49601 25334 56751 25336
rect 49601 25331 49667 25334
rect 56685 25331 56751 25334
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 55213 24986 55279 24989
rect 59200 24986 60000 25016
rect 55213 24984 60000 24986
rect 55213 24928 55218 24984
rect 55274 24928 60000 24984
rect 55213 24926 60000 24928
rect 55213 24923 55279 24926
rect 59200 24896 60000 24926
rect 0 24850 800 24880
rect 2773 24850 2839 24853
rect 0 24848 2839 24850
rect 0 24792 2778 24848
rect 2834 24792 2839 24848
rect 0 24790 2839 24792
rect 0 24760 800 24790
rect 2773 24787 2839 24790
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 50288 24512 50608 24513
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 24447 50608 24448
rect 58157 24442 58223 24445
rect 59200 24442 60000 24472
rect 58157 24440 60000 24442
rect 58157 24384 58162 24440
rect 58218 24384 60000 24440
rect 58157 24382 60000 24384
rect 58157 24379 58223 24382
rect 59200 24352 60000 24382
rect 4208 23968 4528 23969
rect 0 23898 800 23928
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 1945 23898 2011 23901
rect 0 23896 2011 23898
rect 0 23840 1950 23896
rect 2006 23840 2011 23896
rect 0 23838 2011 23840
rect 0 23808 800 23838
rect 1945 23835 2011 23838
rect 56961 23898 57027 23901
rect 59200 23898 60000 23928
rect 56961 23896 60000 23898
rect 56961 23840 56966 23896
rect 57022 23840 60000 23896
rect 56961 23838 60000 23840
rect 56961 23835 57027 23838
rect 59200 23808 60000 23838
rect 55213 23490 55279 23493
rect 59200 23490 60000 23520
rect 55213 23488 60000 23490
rect 55213 23432 55218 23488
rect 55274 23432 60000 23488
rect 55213 23430 60000 23432
rect 55213 23427 55279 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 50288 23424 50608 23425
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 59200 23400 60000 23430
rect 50288 23359 50608 23360
rect 50429 23218 50495 23221
rect 57145 23218 57211 23221
rect 50429 23216 57211 23218
rect 50429 23160 50434 23216
rect 50490 23160 57150 23216
rect 57206 23160 57211 23216
rect 50429 23158 57211 23160
rect 50429 23155 50495 23158
rect 57145 23155 57211 23158
rect 0 22946 800 22976
rect 1945 22946 2011 22949
rect 0 22944 2011 22946
rect 0 22888 1950 22944
rect 2006 22888 2011 22944
rect 0 22886 2011 22888
rect 0 22856 800 22886
rect 1945 22883 2011 22886
rect 57881 22946 57947 22949
rect 59200 22946 60000 22976
rect 57881 22944 60000 22946
rect 57881 22888 57886 22944
rect 57942 22888 60000 22944
rect 57881 22886 60000 22888
rect 57881 22883 57947 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 59200 22856 60000 22886
rect 34928 22815 35248 22816
rect 51717 22810 51783 22813
rect 52729 22810 52795 22813
rect 51717 22808 52795 22810
rect 51717 22752 51722 22808
rect 51778 22752 52734 22808
rect 52790 22752 52795 22808
rect 51717 22750 52795 22752
rect 51717 22747 51783 22750
rect 52729 22747 52795 22750
rect 57421 22402 57487 22405
rect 59200 22402 60000 22432
rect 57421 22400 60000 22402
rect 57421 22344 57426 22400
rect 57482 22344 60000 22400
rect 57421 22342 60000 22344
rect 57421 22339 57487 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 50288 22336 50608 22337
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 59200 22312 60000 22342
rect 50288 22271 50608 22272
rect 0 21994 800 22024
rect 2037 21994 2103 21997
rect 0 21992 2103 21994
rect 0 21936 2042 21992
rect 2098 21936 2103 21992
rect 0 21934 2103 21936
rect 0 21904 800 21934
rect 2037 21931 2103 21934
rect 55213 21858 55279 21861
rect 59200 21858 60000 21888
rect 55213 21856 60000 21858
rect 55213 21800 55218 21856
rect 55274 21800 60000 21856
rect 55213 21798 60000 21800
rect 55213 21795 55279 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 59200 21768 60000 21798
rect 34928 21727 35248 21728
rect 56501 21314 56567 21317
rect 59200 21314 60000 21344
rect 56501 21312 60000 21314
rect 56501 21256 56506 21312
rect 56562 21256 60000 21312
rect 56501 21254 60000 21256
rect 56501 21251 56567 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 50288 21248 50608 21249
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 59200 21224 60000 21254
rect 50288 21183 50608 21184
rect 0 21042 800 21072
rect 2773 21042 2839 21045
rect 0 21040 2839 21042
rect 0 20984 2778 21040
rect 2834 20984 2839 21040
rect 0 20982 2839 20984
rect 0 20952 800 20982
rect 2773 20979 2839 20982
rect 52637 21042 52703 21045
rect 54293 21042 54359 21045
rect 52637 21040 54359 21042
rect 52637 20984 52642 21040
rect 52698 20984 54298 21040
rect 54354 20984 54359 21040
rect 52637 20982 54359 20984
rect 52637 20979 52703 20982
rect 54293 20979 54359 20982
rect 51625 20906 51691 20909
rect 55489 20906 55555 20909
rect 51625 20904 55555 20906
rect 51625 20848 51630 20904
rect 51686 20848 55494 20904
rect 55550 20848 55555 20904
rect 51625 20846 55555 20848
rect 51625 20843 51691 20846
rect 55489 20843 55555 20846
rect 57513 20906 57579 20909
rect 59200 20906 60000 20936
rect 57513 20904 60000 20906
rect 57513 20848 57518 20904
rect 57574 20848 60000 20904
rect 57513 20846 60000 20848
rect 57513 20843 57579 20846
rect 59200 20816 60000 20846
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 51993 20498 52059 20501
rect 53281 20498 53347 20501
rect 51993 20496 53347 20498
rect 51993 20440 51998 20496
rect 52054 20440 53286 20496
rect 53342 20440 53347 20496
rect 51993 20438 53347 20440
rect 51993 20435 52059 20438
rect 53281 20435 53347 20438
rect 55305 20362 55371 20365
rect 59200 20362 60000 20392
rect 55305 20360 60000 20362
rect 55305 20304 55310 20360
rect 55366 20304 60000 20360
rect 55305 20302 60000 20304
rect 55305 20299 55371 20302
rect 59200 20272 60000 20302
rect 19568 20160 19888 20161
rect 0 20090 800 20120
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 50288 20160 50608 20161
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 20095 50608 20096
rect 1945 20090 2011 20093
rect 0 20088 2011 20090
rect 0 20032 1950 20088
rect 2006 20032 2011 20088
rect 0 20030 2011 20032
rect 0 20000 800 20030
rect 1945 20027 2011 20030
rect 48405 19954 48471 19957
rect 53097 19954 53163 19957
rect 54661 19954 54727 19957
rect 48405 19952 54727 19954
rect 48405 19896 48410 19952
rect 48466 19896 53102 19952
rect 53158 19896 54666 19952
rect 54722 19896 54727 19952
rect 48405 19894 54727 19896
rect 48405 19891 48471 19894
rect 53097 19891 53163 19894
rect 54661 19891 54727 19894
rect 53005 19818 53071 19821
rect 54569 19818 54635 19821
rect 53005 19816 54635 19818
rect 53005 19760 53010 19816
rect 53066 19760 54574 19816
rect 54630 19760 54635 19816
rect 53005 19758 54635 19760
rect 53005 19755 53071 19758
rect 54569 19755 54635 19758
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 51533 19410 51599 19413
rect 54753 19410 54819 19413
rect 51533 19408 54819 19410
rect 51533 19352 51538 19408
rect 51594 19352 54758 19408
rect 54814 19352 54819 19408
rect 51533 19350 54819 19352
rect 51533 19347 51599 19350
rect 54753 19347 54819 19350
rect 52545 19274 52611 19277
rect 53373 19274 53439 19277
rect 52545 19272 53439 19274
rect 52545 19216 52550 19272
rect 52606 19216 53378 19272
rect 53434 19216 53439 19272
rect 52545 19214 53439 19216
rect 52545 19211 52611 19214
rect 53373 19211 53439 19214
rect 57053 19274 57119 19277
rect 59200 19274 60000 19304
rect 57053 19272 60000 19274
rect 57053 19216 57058 19272
rect 57114 19216 60000 19272
rect 57053 19214 60000 19216
rect 57053 19211 57119 19214
rect 59200 19184 60000 19214
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 50288 19072 50608 19073
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 19007 50608 19008
rect 51073 19002 51139 19005
rect 56961 19002 57027 19005
rect 51073 19000 57027 19002
rect 51073 18944 51078 19000
rect 51134 18944 56966 19000
rect 57022 18944 57027 19000
rect 51073 18942 57027 18944
rect 51073 18939 51139 18942
rect 56961 18939 57027 18942
rect 50613 18866 50679 18869
rect 51809 18866 51875 18869
rect 50613 18864 51875 18866
rect 50613 18808 50618 18864
rect 50674 18808 51814 18864
rect 51870 18808 51875 18864
rect 50613 18806 51875 18808
rect 50613 18803 50679 18806
rect 51809 18803 51875 18806
rect 52269 18866 52335 18869
rect 53189 18866 53255 18869
rect 52269 18864 53255 18866
rect 52269 18808 52274 18864
rect 52330 18808 53194 18864
rect 53250 18808 53255 18864
rect 52269 18806 53255 18808
rect 52269 18803 52335 18806
rect 53189 18803 53255 18806
rect 55213 18730 55279 18733
rect 59200 18730 60000 18760
rect 55213 18728 60000 18730
rect 55213 18672 55218 18728
rect 55274 18672 60000 18728
rect 55213 18670 60000 18672
rect 55213 18667 55279 18670
rect 59200 18640 60000 18670
rect 50705 18594 50771 18597
rect 51257 18594 51323 18597
rect 50705 18592 51323 18594
rect 50705 18536 50710 18592
rect 50766 18536 51262 18592
rect 51318 18536 51323 18592
rect 50705 18534 51323 18536
rect 50705 18531 50771 18534
rect 51257 18531 51323 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 50153 18458 50219 18461
rect 56777 18458 56843 18461
rect 50153 18456 56843 18458
rect 50153 18400 50158 18456
rect 50214 18400 56782 18456
rect 56838 18400 56843 18456
rect 50153 18398 56843 18400
rect 50153 18395 50219 18398
rect 56777 18395 56843 18398
rect 58157 18322 58223 18325
rect 59200 18322 60000 18352
rect 58157 18320 60000 18322
rect 58157 18264 58162 18320
rect 58218 18264 60000 18320
rect 58157 18262 60000 18264
rect 58157 18259 58223 18262
rect 59200 18232 60000 18262
rect 0 18186 800 18216
rect 1945 18186 2011 18189
rect 0 18184 2011 18186
rect 0 18128 1950 18184
rect 2006 18128 2011 18184
rect 0 18126 2011 18128
rect 0 18096 800 18126
rect 1945 18123 2011 18126
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 50288 17984 50608 17985
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 17919 50608 17920
rect 53097 17778 53163 17781
rect 54937 17778 55003 17781
rect 53097 17776 55003 17778
rect 53097 17720 53102 17776
rect 53158 17720 54942 17776
rect 54998 17720 55003 17776
rect 53097 17718 55003 17720
rect 53097 17715 53163 17718
rect 54937 17715 55003 17718
rect 57053 17778 57119 17781
rect 59200 17778 60000 17808
rect 57053 17776 60000 17778
rect 57053 17720 57058 17776
rect 57114 17720 60000 17776
rect 57053 17718 60000 17720
rect 57053 17715 57119 17718
rect 59200 17688 60000 17718
rect 51349 17642 51415 17645
rect 54753 17642 54819 17645
rect 51349 17640 54819 17642
rect 51349 17584 51354 17640
rect 51410 17584 54758 17640
rect 54814 17584 54819 17640
rect 51349 17582 54819 17584
rect 51349 17579 51415 17582
rect 54753 17579 54819 17582
rect 52085 17506 52151 17509
rect 53925 17506 53991 17509
rect 52085 17504 53991 17506
rect 52085 17448 52090 17504
rect 52146 17448 53930 17504
rect 53986 17448 53991 17504
rect 52085 17446 53991 17448
rect 52085 17443 52151 17446
rect 53925 17443 53991 17446
rect 4208 17440 4528 17441
rect 0 17370 800 17400
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 800 17310
rect 1945 17307 2011 17310
rect 50521 17370 50587 17373
rect 51441 17370 51507 17373
rect 54017 17370 54083 17373
rect 55673 17370 55739 17373
rect 50521 17368 55739 17370
rect 50521 17312 50526 17368
rect 50582 17312 51446 17368
rect 51502 17312 54022 17368
rect 54078 17312 55678 17368
rect 55734 17312 55739 17368
rect 50521 17310 55739 17312
rect 50521 17307 50587 17310
rect 51441 17307 51507 17310
rect 54017 17307 54083 17310
rect 55673 17307 55739 17310
rect 55213 17234 55279 17237
rect 59200 17234 60000 17264
rect 55213 17232 60000 17234
rect 55213 17176 55218 17232
rect 55274 17176 60000 17232
rect 55213 17174 60000 17176
rect 55213 17171 55279 17174
rect 59200 17144 60000 17174
rect 49877 17098 49943 17101
rect 57145 17098 57211 17101
rect 49877 17096 57211 17098
rect 49877 17040 49882 17096
rect 49938 17040 57150 17096
rect 57206 17040 57211 17096
rect 49877 17038 57211 17040
rect 49877 17035 49943 17038
rect 57145 17035 57211 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 50288 16896 50608 16897
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 16831 50608 16832
rect 53189 16690 53255 16693
rect 54201 16690 54267 16693
rect 53189 16688 54267 16690
rect 53189 16632 53194 16688
rect 53250 16632 54206 16688
rect 54262 16632 54267 16688
rect 53189 16630 54267 16632
rect 53189 16627 53255 16630
rect 54201 16627 54267 16630
rect 58157 16690 58223 16693
rect 59200 16690 60000 16720
rect 58157 16688 60000 16690
rect 58157 16632 58162 16688
rect 58218 16632 60000 16688
rect 58157 16630 60000 16632
rect 58157 16627 58223 16630
rect 59200 16600 60000 16630
rect 52821 16554 52887 16557
rect 54477 16554 54543 16557
rect 52821 16552 54543 16554
rect 52821 16496 52826 16552
rect 52882 16496 54482 16552
rect 54538 16496 54543 16552
rect 52821 16494 54543 16496
rect 52821 16491 52887 16494
rect 54477 16491 54543 16494
rect 0 16418 800 16448
rect 1945 16418 2011 16421
rect 0 16416 2011 16418
rect 0 16360 1950 16416
rect 2006 16360 2011 16416
rect 0 16358 2011 16360
rect 0 16328 800 16358
rect 1945 16355 2011 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 57421 16146 57487 16149
rect 59200 16146 60000 16176
rect 57421 16144 60000 16146
rect 57421 16088 57426 16144
rect 57482 16088 60000 16144
rect 57421 16086 60000 16088
rect 57421 16083 57487 16086
rect 59200 16056 60000 16086
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 50288 15808 50608 15809
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 15743 50608 15744
rect 59200 15738 60000 15768
rect 57930 15678 60000 15738
rect 49693 15602 49759 15605
rect 57930 15602 57990 15678
rect 59200 15648 60000 15678
rect 49693 15600 57990 15602
rect 49693 15544 49698 15600
rect 49754 15544 57990 15600
rect 49693 15542 57990 15544
rect 49693 15539 49759 15542
rect 0 15466 800 15496
rect 2773 15466 2839 15469
rect 0 15464 2839 15466
rect 0 15408 2778 15464
rect 2834 15408 2839 15464
rect 0 15406 2839 15408
rect 0 15376 800 15406
rect 2773 15403 2839 15406
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 57881 15194 57947 15197
rect 59200 15194 60000 15224
rect 57881 15192 60000 15194
rect 57881 15136 57886 15192
rect 57942 15136 60000 15192
rect 57881 15134 60000 15136
rect 57881 15131 57947 15134
rect 59200 15104 60000 15134
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 50288 14720 50608 14721
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 14655 50608 14656
rect 55489 14650 55555 14653
rect 59200 14650 60000 14680
rect 55489 14648 60000 14650
rect 55489 14592 55494 14648
rect 55550 14592 60000 14648
rect 55489 14590 60000 14592
rect 55489 14587 55555 14590
rect 59200 14560 60000 14590
rect 0 14514 800 14544
rect 1945 14514 2011 14517
rect 0 14512 2011 14514
rect 0 14456 1950 14512
rect 2006 14456 2011 14512
rect 0 14454 2011 14456
rect 0 14424 800 14454
rect 1945 14451 2011 14454
rect 50429 14514 50495 14517
rect 52545 14514 52611 14517
rect 53925 14514 53991 14517
rect 50429 14512 53991 14514
rect 50429 14456 50434 14512
rect 50490 14456 52550 14512
rect 52606 14456 53930 14512
rect 53986 14456 53991 14512
rect 50429 14454 53991 14456
rect 50429 14451 50495 14454
rect 52545 14451 52611 14454
rect 53925 14451 53991 14454
rect 50981 14242 51047 14245
rect 56041 14242 56107 14245
rect 50981 14240 56107 14242
rect 50981 14184 50986 14240
rect 51042 14184 56046 14240
rect 56102 14184 56107 14240
rect 50981 14182 56107 14184
rect 50981 14179 51047 14182
rect 56041 14179 56107 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 49141 14106 49207 14109
rect 59200 14106 60000 14136
rect 49141 14104 60000 14106
rect 49141 14048 49146 14104
rect 49202 14048 60000 14104
rect 49141 14046 60000 14048
rect 49141 14043 49207 14046
rect 59200 14016 60000 14046
rect 50981 13970 51047 13973
rect 52361 13970 52427 13973
rect 50981 13968 52427 13970
rect 50981 13912 50986 13968
rect 51042 13912 52366 13968
rect 52422 13912 52427 13968
rect 50981 13910 52427 13912
rect 50981 13907 51047 13910
rect 52361 13907 52427 13910
rect 52545 13834 52611 13837
rect 55213 13834 55279 13837
rect 52545 13832 55279 13834
rect 52545 13776 52550 13832
rect 52606 13776 55218 13832
rect 55274 13776 55279 13832
rect 52545 13774 55279 13776
rect 52545 13771 52611 13774
rect 55213 13771 55279 13774
rect 50705 13698 50771 13701
rect 56133 13698 56199 13701
rect 50705 13696 56199 13698
rect 50705 13640 50710 13696
rect 50766 13640 56138 13696
rect 56194 13640 56199 13696
rect 50705 13638 56199 13640
rect 50705 13635 50771 13638
rect 56133 13635 56199 13638
rect 19568 13632 19888 13633
rect 0 13562 800 13592
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 50288 13632 50608 13633
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 13567 50608 13568
rect 1945 13562 2011 13565
rect 0 13560 2011 13562
rect 0 13504 1950 13560
rect 2006 13504 2011 13560
rect 0 13502 2011 13504
rect 0 13472 800 13502
rect 1945 13499 2011 13502
rect 57053 13562 57119 13565
rect 59200 13562 60000 13592
rect 57053 13560 60000 13562
rect 57053 13504 57058 13560
rect 57114 13504 60000 13560
rect 57053 13502 60000 13504
rect 57053 13499 57119 13502
rect 59200 13472 60000 13502
rect 57329 13154 57395 13157
rect 59200 13154 60000 13184
rect 57329 13152 60000 13154
rect 57329 13096 57334 13152
rect 57390 13096 60000 13152
rect 57329 13094 60000 13096
rect 57329 13091 57395 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 59200 13064 60000 13094
rect 34928 13023 35248 13024
rect 0 12610 800 12640
rect 1945 12610 2011 12613
rect 0 12608 2011 12610
rect 0 12552 1950 12608
rect 2006 12552 2011 12608
rect 0 12550 2011 12552
rect 0 12520 800 12550
rect 1945 12547 2011 12550
rect 55213 12610 55279 12613
rect 59200 12610 60000 12640
rect 55213 12608 60000 12610
rect 55213 12552 55218 12608
rect 55274 12552 60000 12608
rect 55213 12550 60000 12552
rect 55213 12547 55279 12550
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 50288 12544 50608 12545
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 59200 12520 60000 12550
rect 50288 12479 50608 12480
rect 50521 12338 50587 12341
rect 52269 12338 52335 12341
rect 53925 12338 53991 12341
rect 50521 12336 53991 12338
rect 50521 12280 50526 12336
rect 50582 12280 52274 12336
rect 52330 12280 53930 12336
rect 53986 12280 53991 12336
rect 50521 12278 53991 12280
rect 50521 12275 50587 12278
rect 52269 12275 52335 12278
rect 53925 12275 53991 12278
rect 57881 12066 57947 12069
rect 59200 12066 60000 12096
rect 57881 12064 60000 12066
rect 57881 12008 57886 12064
rect 57942 12008 60000 12064
rect 57881 12006 60000 12008
rect 57881 12003 57947 12006
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 59200 11976 60000 12006
rect 34928 11935 35248 11936
rect 0 11658 800 11688
rect 2773 11658 2839 11661
rect 0 11656 2839 11658
rect 0 11600 2778 11656
rect 2834 11600 2839 11656
rect 0 11598 2839 11600
rect 0 11568 800 11598
rect 2773 11595 2839 11598
rect 49325 11658 49391 11661
rect 57145 11658 57211 11661
rect 49325 11656 57211 11658
rect 49325 11600 49330 11656
rect 49386 11600 57150 11656
rect 57206 11600 57211 11656
rect 49325 11598 57211 11600
rect 49325 11595 49391 11598
rect 57145 11595 57211 11598
rect 58157 11522 58223 11525
rect 59200 11522 60000 11552
rect 58157 11520 60000 11522
rect 58157 11464 58162 11520
rect 58218 11464 60000 11520
rect 58157 11462 60000 11464
rect 58157 11459 58223 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 50288 11456 50608 11457
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 59200 11432 60000 11462
rect 50288 11391 50608 11392
rect 55213 10978 55279 10981
rect 59200 10978 60000 11008
rect 55213 10976 60000 10978
rect 55213 10920 55218 10976
rect 55274 10920 60000 10976
rect 55213 10918 60000 10920
rect 55213 10915 55279 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 59200 10888 60000 10918
rect 34928 10847 35248 10848
rect 0 10706 800 10736
rect 1945 10706 2011 10709
rect 0 10704 2011 10706
rect 0 10648 1950 10704
rect 2006 10648 2011 10704
rect 0 10646 2011 10648
rect 0 10616 800 10646
rect 1945 10643 2011 10646
rect 58157 10570 58223 10573
rect 59200 10570 60000 10600
rect 58157 10568 60000 10570
rect 58157 10512 58162 10568
rect 58218 10512 60000 10568
rect 58157 10510 60000 10512
rect 58157 10507 58223 10510
rect 59200 10480 60000 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 50288 10368 50608 10369
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 10303 50608 10304
rect 57053 10026 57119 10029
rect 59200 10026 60000 10056
rect 57053 10024 60000 10026
rect 57053 9968 57058 10024
rect 57114 9968 60000 10024
rect 57053 9966 60000 9968
rect 57053 9963 57119 9966
rect 59200 9936 60000 9966
rect 4208 9824 4528 9825
rect 0 9754 800 9784
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 1945 9754 2011 9757
rect 0 9752 2011 9754
rect 0 9696 1950 9752
rect 2006 9696 2011 9752
rect 0 9694 2011 9696
rect 0 9664 800 9694
rect 1945 9691 2011 9694
rect 55213 9482 55279 9485
rect 59200 9482 60000 9512
rect 55213 9480 60000 9482
rect 55213 9424 55218 9480
rect 55274 9424 60000 9480
rect 55213 9422 60000 9424
rect 55213 9419 55279 9422
rect 59200 9392 60000 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 50288 9280 50608 9281
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 9215 50608 9216
rect 0 8938 800 8968
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8848 800 8878
rect 2773 8875 2839 8878
rect 58157 8938 58223 8941
rect 59200 8938 60000 8968
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8848 60000 8878
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 58157 8394 58223 8397
rect 59200 8394 60000 8424
rect 58157 8392 60000 8394
rect 58157 8336 58162 8392
rect 58218 8336 60000 8392
rect 58157 8334 60000 8336
rect 58157 8331 58223 8334
rect 59200 8304 60000 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 50288 8192 50608 8193
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 8127 50608 8128
rect 56593 8122 56659 8125
rect 51030 8120 56659 8122
rect 51030 8064 56598 8120
rect 56654 8064 56659 8120
rect 51030 8062 56659 8064
rect 0 7986 800 8016
rect 2037 7986 2103 7989
rect 0 7984 2103 7986
rect 0 7928 2042 7984
rect 2098 7928 2103 7984
rect 0 7926 2103 7928
rect 0 7896 800 7926
rect 2037 7923 2103 7926
rect 49325 7986 49391 7989
rect 51030 7986 51090 8062
rect 56593 8059 56659 8062
rect 49325 7984 51090 7986
rect 49325 7928 49330 7984
rect 49386 7928 51090 7984
rect 49325 7926 51090 7928
rect 55213 7986 55279 7989
rect 59200 7986 60000 8016
rect 55213 7984 60000 7986
rect 55213 7928 55218 7984
rect 55274 7928 60000 7984
rect 55213 7926 60000 7928
rect 49325 7923 49391 7926
rect 55213 7923 55279 7926
rect 59200 7896 60000 7926
rect 48681 7850 48747 7853
rect 57329 7850 57395 7853
rect 48681 7848 57395 7850
rect 48681 7792 48686 7848
rect 48742 7792 57334 7848
rect 57390 7792 57395 7848
rect 48681 7790 57395 7792
rect 48681 7787 48747 7790
rect 57329 7787 57395 7790
rect 48405 7714 48471 7717
rect 55397 7714 55463 7717
rect 48405 7712 55463 7714
rect 48405 7656 48410 7712
rect 48466 7656 55402 7712
rect 55458 7656 55463 7712
rect 48405 7654 55463 7656
rect 48405 7651 48471 7654
rect 55397 7651 55463 7654
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 58157 7442 58223 7445
rect 59200 7442 60000 7472
rect 58157 7440 60000 7442
rect 58157 7384 58162 7440
rect 58218 7384 60000 7440
rect 58157 7382 60000 7384
rect 58157 7379 58223 7382
rect 59200 7352 60000 7382
rect 19568 7104 19888 7105
rect 0 7034 800 7064
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 50288 7104 50608 7105
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 7039 50608 7040
rect 1945 7034 2011 7037
rect 0 7032 2011 7034
rect 0 6976 1950 7032
rect 2006 6976 2011 7032
rect 0 6974 2011 6976
rect 0 6944 800 6974
rect 1945 6971 2011 6974
rect 48773 6898 48839 6901
rect 49693 6898 49759 6901
rect 48773 6896 49759 6898
rect 48773 6840 48778 6896
rect 48834 6840 49698 6896
rect 49754 6840 49759 6896
rect 48773 6838 49759 6840
rect 48773 6835 48839 6838
rect 49693 6835 49759 6838
rect 57145 6898 57211 6901
rect 59200 6898 60000 6928
rect 57145 6896 60000 6898
rect 57145 6840 57150 6896
rect 57206 6840 60000 6896
rect 57145 6838 60000 6840
rect 57145 6835 57211 6838
rect 59200 6808 60000 6838
rect 48681 6762 48747 6765
rect 49785 6762 49851 6765
rect 50981 6762 51047 6765
rect 48681 6760 51047 6762
rect 48681 6704 48686 6760
rect 48742 6704 49790 6760
rect 49846 6704 50986 6760
rect 51042 6704 51047 6760
rect 48681 6702 51047 6704
rect 48681 6699 48747 6702
rect 49785 6699 49851 6702
rect 50981 6699 51047 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 55305 6354 55371 6357
rect 59200 6354 60000 6384
rect 55305 6352 60000 6354
rect 55305 6296 55310 6352
rect 55366 6296 60000 6352
rect 55305 6294 60000 6296
rect 55305 6291 55371 6294
rect 59200 6264 60000 6294
rect 0 6082 800 6112
rect 1945 6082 2011 6085
rect 0 6080 2011 6082
rect 0 6024 1950 6080
rect 2006 6024 2011 6080
rect 0 6022 2011 6024
rect 0 5992 800 6022
rect 1945 6019 2011 6022
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 50288 6016 50608 6017
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 5951 50608 5952
rect 49601 5810 49667 5813
rect 50981 5810 51047 5813
rect 49601 5808 51047 5810
rect 49601 5752 49606 5808
rect 49662 5752 50986 5808
rect 51042 5752 51047 5808
rect 49601 5750 51047 5752
rect 49601 5747 49667 5750
rect 50981 5747 51047 5750
rect 58157 5810 58223 5813
rect 59200 5810 60000 5840
rect 58157 5808 60000 5810
rect 58157 5752 58162 5808
rect 58218 5752 60000 5808
rect 58157 5750 60000 5752
rect 58157 5747 58223 5750
rect 59200 5720 60000 5750
rect 50889 5674 50955 5677
rect 52821 5674 52887 5677
rect 50889 5672 52887 5674
rect 50889 5616 50894 5672
rect 50950 5616 52826 5672
rect 52882 5616 52887 5672
rect 50889 5614 52887 5616
rect 50889 5611 50955 5614
rect 52821 5611 52887 5614
rect 49969 5538 50035 5541
rect 56685 5538 56751 5541
rect 49969 5536 56751 5538
rect 49969 5480 49974 5536
rect 50030 5480 56690 5536
rect 56746 5480 56751 5536
rect 49969 5478 56751 5480
rect 49969 5475 50035 5478
rect 56685 5475 56751 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 56961 5402 57027 5405
rect 59200 5402 60000 5432
rect 56961 5400 60000 5402
rect 56961 5344 56966 5400
rect 57022 5344 60000 5400
rect 56961 5342 60000 5344
rect 56961 5339 57027 5342
rect 59200 5312 60000 5342
rect 49417 5266 49483 5269
rect 51165 5266 51231 5269
rect 49417 5264 51231 5266
rect 49417 5208 49422 5264
rect 49478 5208 51170 5264
rect 51226 5208 51231 5264
rect 49417 5206 51231 5208
rect 49417 5203 49483 5206
rect 51165 5203 51231 5206
rect 0 5130 800 5160
rect 2773 5130 2839 5133
rect 0 5128 2839 5130
rect 0 5072 2778 5128
rect 2834 5072 2839 5128
rect 0 5070 2839 5072
rect 0 5040 800 5070
rect 2773 5067 2839 5070
rect 49233 5130 49299 5133
rect 50889 5130 50955 5133
rect 49233 5128 50955 5130
rect 49233 5072 49238 5128
rect 49294 5072 50894 5128
rect 50950 5072 50955 5128
rect 49233 5070 50955 5072
rect 49233 5067 49299 5070
rect 50889 5067 50955 5070
rect 51073 5130 51139 5133
rect 54385 5130 54451 5133
rect 51073 5128 54451 5130
rect 51073 5072 51078 5128
rect 51134 5072 54390 5128
rect 54446 5072 54451 5128
rect 51073 5070 54451 5072
rect 51073 5067 51139 5070
rect 54385 5067 54451 5070
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 50288 4928 50608 4929
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 4863 50608 4864
rect 55213 4858 55279 4861
rect 59200 4858 60000 4888
rect 55213 4856 60000 4858
rect 55213 4800 55218 4856
rect 55274 4800 60000 4856
rect 55213 4798 60000 4800
rect 55213 4795 55279 4798
rect 59200 4768 60000 4798
rect 45001 4586 45067 4589
rect 48129 4586 48195 4589
rect 45001 4584 48195 4586
rect 45001 4528 45006 4584
rect 45062 4528 48134 4584
rect 48190 4528 48195 4584
rect 45001 4526 48195 4528
rect 45001 4523 45067 4526
rect 48129 4523 48195 4526
rect 50705 4586 50771 4589
rect 57237 4586 57303 4589
rect 50705 4584 57303 4586
rect 50705 4528 50710 4584
rect 50766 4528 57242 4584
rect 57298 4528 57303 4584
rect 50705 4526 57303 4528
rect 50705 4523 50771 4526
rect 57237 4523 57303 4526
rect 50889 4450 50955 4453
rect 51073 4450 51139 4453
rect 50889 4448 51174 4450
rect 50889 4392 50894 4448
rect 50950 4392 51078 4448
rect 51134 4392 51174 4448
rect 50889 4390 51174 4392
rect 50889 4387 50955 4390
rect 51073 4387 51139 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 56961 4314 57027 4317
rect 59200 4314 60000 4344
rect 56961 4312 60000 4314
rect 56961 4256 56966 4312
rect 57022 4256 60000 4312
rect 56961 4254 60000 4256
rect 56961 4251 57027 4254
rect 59200 4224 60000 4254
rect 0 4178 800 4208
rect 2865 4178 2931 4181
rect 0 4176 2931 4178
rect 0 4120 2870 4176
rect 2926 4120 2931 4176
rect 0 4118 2931 4120
rect 0 4088 800 4118
rect 2865 4115 2931 4118
rect 50061 4178 50127 4181
rect 56685 4178 56751 4181
rect 50061 4176 56751 4178
rect 50061 4120 50066 4176
rect 50122 4120 56690 4176
rect 56746 4120 56751 4176
rect 50061 4118 56751 4120
rect 50061 4115 50127 4118
rect 56685 4115 56751 4118
rect 47209 4042 47275 4045
rect 52453 4042 52519 4045
rect 47209 4040 52519 4042
rect 47209 3984 47214 4040
rect 47270 3984 52458 4040
rect 52514 3984 52519 4040
rect 47209 3982 52519 3984
rect 47209 3979 47275 3982
rect 52453 3979 52519 3982
rect 52729 4042 52795 4045
rect 55213 4042 55279 4045
rect 55949 4042 56015 4045
rect 52729 4040 56015 4042
rect 52729 3984 52734 4040
rect 52790 3984 55218 4040
rect 55274 3984 55954 4040
rect 56010 3984 56015 4040
rect 52729 3982 56015 3984
rect 52729 3979 52795 3982
rect 55213 3979 55279 3982
rect 55949 3979 56015 3982
rect 54201 3906 54267 3909
rect 56777 3906 56843 3909
rect 54201 3904 56843 3906
rect 54201 3848 54206 3904
rect 54262 3848 56782 3904
rect 56838 3848 56843 3904
rect 54201 3846 56843 3848
rect 54201 3843 54267 3846
rect 56777 3843 56843 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 50288 3840 50608 3841
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 3775 50608 3776
rect 56041 3770 56107 3773
rect 59200 3770 60000 3800
rect 56041 3768 60000 3770
rect 56041 3712 56046 3768
rect 56102 3712 60000 3768
rect 56041 3710 60000 3712
rect 56041 3707 56107 3710
rect 59200 3680 60000 3710
rect 49141 3362 49207 3365
rect 55489 3362 55555 3365
rect 49141 3360 55555 3362
rect 49141 3304 49146 3360
rect 49202 3304 55494 3360
rect 55550 3304 55555 3360
rect 49141 3302 55555 3304
rect 49141 3299 49207 3302
rect 55489 3299 55555 3302
rect 4208 3296 4528 3297
rect 0 3226 800 3256
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 2773 3226 2839 3229
rect 0 3224 2839 3226
rect 0 3168 2778 3224
rect 2834 3168 2839 3224
rect 0 3166 2839 3168
rect 0 3136 800 3166
rect 2773 3163 2839 3166
rect 55213 3226 55279 3229
rect 59200 3226 60000 3256
rect 55213 3224 60000 3226
rect 55213 3168 55218 3224
rect 55274 3168 60000 3224
rect 55213 3166 60000 3168
rect 55213 3163 55279 3166
rect 59200 3136 60000 3166
rect 49601 3090 49667 3093
rect 57053 3090 57119 3093
rect 49601 3088 57119 3090
rect 49601 3032 49606 3088
rect 49662 3032 57058 3088
rect 57114 3032 57119 3088
rect 49601 3030 57119 3032
rect 49601 3027 49667 3030
rect 57053 3027 57119 3030
rect 54845 2954 54911 2957
rect 55857 2954 55923 2957
rect 54845 2952 55923 2954
rect 54845 2896 54850 2952
rect 54906 2896 55862 2952
rect 55918 2896 55923 2952
rect 54845 2894 55923 2896
rect 54845 2891 54911 2894
rect 55857 2891 55923 2894
rect 58157 2818 58223 2821
rect 59200 2818 60000 2848
rect 58157 2816 60000 2818
rect 58157 2760 58162 2816
rect 58218 2760 60000 2816
rect 58157 2758 60000 2760
rect 58157 2755 58223 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 50288 2752 50608 2753
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 59200 2728 60000 2758
rect 50288 2687 50608 2688
rect 0 2274 800 2304
rect 4061 2274 4127 2277
rect 0 2272 4127 2274
rect 0 2216 4066 2272
rect 4122 2216 4127 2272
rect 0 2214 4127 2216
rect 0 2184 800 2214
rect 4061 2211 4127 2214
rect 55765 2274 55831 2277
rect 59200 2274 60000 2304
rect 55765 2272 60000 2274
rect 55765 2216 55770 2272
rect 55826 2216 60000 2272
rect 55765 2214 60000 2216
rect 55765 2211 55831 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 59200 2184 60000 2214
rect 34928 2143 35248 2144
rect 55213 1730 55279 1733
rect 59200 1730 60000 1760
rect 55213 1728 60000 1730
rect 55213 1672 55218 1728
rect 55274 1672 60000 1728
rect 55213 1670 60000 1672
rect 55213 1667 55279 1670
rect 59200 1640 60000 1670
rect 0 1322 800 1352
rect 2865 1322 2931 1325
rect 0 1320 2931 1322
rect 0 1264 2870 1320
rect 2926 1264 2931 1320
rect 0 1262 2931 1264
rect 0 1232 800 1262
rect 2865 1259 2931 1262
rect 57881 1186 57947 1189
rect 59200 1186 60000 1216
rect 57881 1184 60000 1186
rect 57881 1128 57886 1184
rect 57942 1128 60000 1184
rect 57881 1126 60000 1128
rect 57881 1123 57947 1126
rect 59200 1096 60000 1126
rect 56409 642 56475 645
rect 59200 642 60000 672
rect 56409 640 60000 642
rect 56409 584 56414 640
rect 56470 584 60000 640
rect 56409 582 60000 584
rect 56409 579 56475 582
rect 59200 552 60000 582
rect 0 506 800 536
rect 2957 506 3023 509
rect 0 504 3023 506
rect 0 448 2962 504
rect 3018 448 3023 504
rect 0 446 3023 448
rect 0 416 800 446
rect 2957 443 3023 446
rect 55213 234 55279 237
rect 59200 234 60000 264
rect 55213 232 60000 234
rect 55213 176 55218 232
rect 55274 176 60000 232
rect 55213 174 60000 176
rect 55213 171 55279 174
rect 59200 144 60000 174
<< via3 >>
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 50296 57148 50360 57152
rect 50296 57092 50300 57148
rect 50300 57092 50356 57148
rect 50356 57092 50360 57148
rect 50296 57088 50360 57092
rect 50376 57148 50440 57152
rect 50376 57092 50380 57148
rect 50380 57092 50436 57148
rect 50436 57092 50440 57148
rect 50376 57088 50440 57092
rect 50456 57148 50520 57152
rect 50456 57092 50460 57148
rect 50460 57092 50516 57148
rect 50516 57092 50520 57148
rect 50456 57088 50520 57092
rect 50536 57148 50600 57152
rect 50536 57092 50540 57148
rect 50540 57092 50596 57148
rect 50596 57092 50600 57148
rect 50536 57088 50600 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 50296 56060 50360 56064
rect 50296 56004 50300 56060
rect 50300 56004 50356 56060
rect 50356 56004 50360 56060
rect 50296 56000 50360 56004
rect 50376 56060 50440 56064
rect 50376 56004 50380 56060
rect 50380 56004 50436 56060
rect 50436 56004 50440 56060
rect 50376 56000 50440 56004
rect 50456 56060 50520 56064
rect 50456 56004 50460 56060
rect 50460 56004 50516 56060
rect 50516 56004 50520 56060
rect 50456 56000 50520 56004
rect 50536 56060 50600 56064
rect 50536 56004 50540 56060
rect 50540 56004 50596 56060
rect 50596 56004 50600 56060
rect 50536 56000 50600 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 50296 54972 50360 54976
rect 50296 54916 50300 54972
rect 50300 54916 50356 54972
rect 50356 54916 50360 54972
rect 50296 54912 50360 54916
rect 50376 54972 50440 54976
rect 50376 54916 50380 54972
rect 50380 54916 50436 54972
rect 50436 54916 50440 54972
rect 50376 54912 50440 54916
rect 50456 54972 50520 54976
rect 50456 54916 50460 54972
rect 50460 54916 50516 54972
rect 50516 54916 50520 54972
rect 50456 54912 50520 54916
rect 50536 54972 50600 54976
rect 50536 54916 50540 54972
rect 50540 54916 50596 54972
rect 50596 54916 50600 54972
rect 50536 54912 50600 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 50296 53884 50360 53888
rect 50296 53828 50300 53884
rect 50300 53828 50356 53884
rect 50356 53828 50360 53884
rect 50296 53824 50360 53828
rect 50376 53884 50440 53888
rect 50376 53828 50380 53884
rect 50380 53828 50436 53884
rect 50436 53828 50440 53884
rect 50376 53824 50440 53828
rect 50456 53884 50520 53888
rect 50456 53828 50460 53884
rect 50460 53828 50516 53884
rect 50516 53828 50520 53884
rect 50456 53824 50520 53828
rect 50536 53884 50600 53888
rect 50536 53828 50540 53884
rect 50540 53828 50596 53884
rect 50596 53828 50600 53884
rect 50536 53824 50600 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 50296 52796 50360 52800
rect 50296 52740 50300 52796
rect 50300 52740 50356 52796
rect 50356 52740 50360 52796
rect 50296 52736 50360 52740
rect 50376 52796 50440 52800
rect 50376 52740 50380 52796
rect 50380 52740 50436 52796
rect 50436 52740 50440 52796
rect 50376 52736 50440 52740
rect 50456 52796 50520 52800
rect 50456 52740 50460 52796
rect 50460 52740 50516 52796
rect 50516 52740 50520 52796
rect 50456 52736 50520 52740
rect 50536 52796 50600 52800
rect 50536 52740 50540 52796
rect 50540 52740 50596 52796
rect 50596 52740 50600 52796
rect 50536 52736 50600 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 50296 51708 50360 51712
rect 50296 51652 50300 51708
rect 50300 51652 50356 51708
rect 50356 51652 50360 51708
rect 50296 51648 50360 51652
rect 50376 51708 50440 51712
rect 50376 51652 50380 51708
rect 50380 51652 50436 51708
rect 50436 51652 50440 51708
rect 50376 51648 50440 51652
rect 50456 51708 50520 51712
rect 50456 51652 50460 51708
rect 50460 51652 50516 51708
rect 50516 51652 50520 51708
rect 50456 51648 50520 51652
rect 50536 51708 50600 51712
rect 50536 51652 50540 51708
rect 50540 51652 50596 51708
rect 50596 51652 50600 51708
rect 50536 51648 50600 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 50296 50620 50360 50624
rect 50296 50564 50300 50620
rect 50300 50564 50356 50620
rect 50356 50564 50360 50620
rect 50296 50560 50360 50564
rect 50376 50620 50440 50624
rect 50376 50564 50380 50620
rect 50380 50564 50436 50620
rect 50436 50564 50440 50620
rect 50376 50560 50440 50564
rect 50456 50620 50520 50624
rect 50456 50564 50460 50620
rect 50460 50564 50516 50620
rect 50516 50564 50520 50620
rect 50456 50560 50520 50564
rect 50536 50620 50600 50624
rect 50536 50564 50540 50620
rect 50540 50564 50596 50620
rect 50596 50564 50600 50620
rect 50536 50560 50600 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 50296 49532 50360 49536
rect 50296 49476 50300 49532
rect 50300 49476 50356 49532
rect 50356 49476 50360 49532
rect 50296 49472 50360 49476
rect 50376 49532 50440 49536
rect 50376 49476 50380 49532
rect 50380 49476 50436 49532
rect 50436 49476 50440 49532
rect 50376 49472 50440 49476
rect 50456 49532 50520 49536
rect 50456 49476 50460 49532
rect 50460 49476 50516 49532
rect 50516 49476 50520 49532
rect 50456 49472 50520 49476
rect 50536 49532 50600 49536
rect 50536 49476 50540 49532
rect 50540 49476 50596 49532
rect 50596 49476 50600 49532
rect 50536 49472 50600 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 50296 48444 50360 48448
rect 50296 48388 50300 48444
rect 50300 48388 50356 48444
rect 50356 48388 50360 48444
rect 50296 48384 50360 48388
rect 50376 48444 50440 48448
rect 50376 48388 50380 48444
rect 50380 48388 50436 48444
rect 50436 48388 50440 48444
rect 50376 48384 50440 48388
rect 50456 48444 50520 48448
rect 50456 48388 50460 48444
rect 50460 48388 50516 48444
rect 50516 48388 50520 48444
rect 50456 48384 50520 48388
rect 50536 48444 50600 48448
rect 50536 48388 50540 48444
rect 50540 48388 50596 48444
rect 50596 48388 50600 48444
rect 50536 48384 50600 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 50296 47356 50360 47360
rect 50296 47300 50300 47356
rect 50300 47300 50356 47356
rect 50356 47300 50360 47356
rect 50296 47296 50360 47300
rect 50376 47356 50440 47360
rect 50376 47300 50380 47356
rect 50380 47300 50436 47356
rect 50436 47300 50440 47356
rect 50376 47296 50440 47300
rect 50456 47356 50520 47360
rect 50456 47300 50460 47356
rect 50460 47300 50516 47356
rect 50516 47300 50520 47356
rect 50456 47296 50520 47300
rect 50536 47356 50600 47360
rect 50536 47300 50540 47356
rect 50540 47300 50596 47356
rect 50596 47300 50600 47356
rect 50536 47296 50600 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 50296 46268 50360 46272
rect 50296 46212 50300 46268
rect 50300 46212 50356 46268
rect 50356 46212 50360 46268
rect 50296 46208 50360 46212
rect 50376 46268 50440 46272
rect 50376 46212 50380 46268
rect 50380 46212 50436 46268
rect 50436 46212 50440 46268
rect 50376 46208 50440 46212
rect 50456 46268 50520 46272
rect 50456 46212 50460 46268
rect 50460 46212 50516 46268
rect 50516 46212 50520 46268
rect 50456 46208 50520 46212
rect 50536 46268 50600 46272
rect 50536 46212 50540 46268
rect 50540 46212 50596 46268
rect 50596 46212 50600 46268
rect 50536 46208 50600 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 50296 45180 50360 45184
rect 50296 45124 50300 45180
rect 50300 45124 50356 45180
rect 50356 45124 50360 45180
rect 50296 45120 50360 45124
rect 50376 45180 50440 45184
rect 50376 45124 50380 45180
rect 50380 45124 50436 45180
rect 50436 45124 50440 45180
rect 50376 45120 50440 45124
rect 50456 45180 50520 45184
rect 50456 45124 50460 45180
rect 50460 45124 50516 45180
rect 50516 45124 50520 45180
rect 50456 45120 50520 45124
rect 50536 45180 50600 45184
rect 50536 45124 50540 45180
rect 50540 45124 50596 45180
rect 50596 45124 50600 45180
rect 50536 45120 50600 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 50296 28860 50360 28864
rect 50296 28804 50300 28860
rect 50300 28804 50356 28860
rect 50356 28804 50360 28860
rect 50296 28800 50360 28804
rect 50376 28860 50440 28864
rect 50376 28804 50380 28860
rect 50380 28804 50436 28860
rect 50436 28804 50440 28860
rect 50376 28800 50440 28804
rect 50456 28860 50520 28864
rect 50456 28804 50460 28860
rect 50460 28804 50516 28860
rect 50516 28804 50520 28860
rect 50456 28800 50520 28804
rect 50536 28860 50600 28864
rect 50536 28804 50540 28860
rect 50540 28804 50596 28860
rect 50596 28804 50600 28860
rect 50536 28800 50600 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 50296 27772 50360 27776
rect 50296 27716 50300 27772
rect 50300 27716 50356 27772
rect 50356 27716 50360 27772
rect 50296 27712 50360 27716
rect 50376 27772 50440 27776
rect 50376 27716 50380 27772
rect 50380 27716 50436 27772
rect 50436 27716 50440 27772
rect 50376 27712 50440 27716
rect 50456 27772 50520 27776
rect 50456 27716 50460 27772
rect 50460 27716 50516 27772
rect 50516 27716 50520 27772
rect 50456 27712 50520 27716
rect 50536 27772 50600 27776
rect 50536 27716 50540 27772
rect 50540 27716 50596 27772
rect 50596 27716 50600 27772
rect 50536 27712 50600 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 50296 26684 50360 26688
rect 50296 26628 50300 26684
rect 50300 26628 50356 26684
rect 50356 26628 50360 26684
rect 50296 26624 50360 26628
rect 50376 26684 50440 26688
rect 50376 26628 50380 26684
rect 50380 26628 50436 26684
rect 50436 26628 50440 26684
rect 50376 26624 50440 26628
rect 50456 26684 50520 26688
rect 50456 26628 50460 26684
rect 50460 26628 50516 26684
rect 50516 26628 50520 26684
rect 50456 26624 50520 26628
rect 50536 26684 50600 26688
rect 50536 26628 50540 26684
rect 50540 26628 50596 26684
rect 50596 26628 50600 26684
rect 50536 26624 50600 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 50296 25596 50360 25600
rect 50296 25540 50300 25596
rect 50300 25540 50356 25596
rect 50356 25540 50360 25596
rect 50296 25536 50360 25540
rect 50376 25596 50440 25600
rect 50376 25540 50380 25596
rect 50380 25540 50436 25596
rect 50436 25540 50440 25596
rect 50376 25536 50440 25540
rect 50456 25596 50520 25600
rect 50456 25540 50460 25596
rect 50460 25540 50516 25596
rect 50516 25540 50520 25596
rect 50456 25536 50520 25540
rect 50536 25596 50600 25600
rect 50536 25540 50540 25596
rect 50540 25540 50596 25596
rect 50596 25540 50600 25596
rect 50536 25536 50600 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 50296 24508 50360 24512
rect 50296 24452 50300 24508
rect 50300 24452 50356 24508
rect 50356 24452 50360 24508
rect 50296 24448 50360 24452
rect 50376 24508 50440 24512
rect 50376 24452 50380 24508
rect 50380 24452 50436 24508
rect 50436 24452 50440 24508
rect 50376 24448 50440 24452
rect 50456 24508 50520 24512
rect 50456 24452 50460 24508
rect 50460 24452 50516 24508
rect 50516 24452 50520 24508
rect 50456 24448 50520 24452
rect 50536 24508 50600 24512
rect 50536 24452 50540 24508
rect 50540 24452 50596 24508
rect 50596 24452 50600 24508
rect 50536 24448 50600 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 50296 23420 50360 23424
rect 50296 23364 50300 23420
rect 50300 23364 50356 23420
rect 50356 23364 50360 23420
rect 50296 23360 50360 23364
rect 50376 23420 50440 23424
rect 50376 23364 50380 23420
rect 50380 23364 50436 23420
rect 50436 23364 50440 23420
rect 50376 23360 50440 23364
rect 50456 23420 50520 23424
rect 50456 23364 50460 23420
rect 50460 23364 50516 23420
rect 50516 23364 50520 23420
rect 50456 23360 50520 23364
rect 50536 23420 50600 23424
rect 50536 23364 50540 23420
rect 50540 23364 50596 23420
rect 50596 23364 50600 23420
rect 50536 23360 50600 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 50296 22332 50360 22336
rect 50296 22276 50300 22332
rect 50300 22276 50356 22332
rect 50356 22276 50360 22332
rect 50296 22272 50360 22276
rect 50376 22332 50440 22336
rect 50376 22276 50380 22332
rect 50380 22276 50436 22332
rect 50436 22276 50440 22332
rect 50376 22272 50440 22276
rect 50456 22332 50520 22336
rect 50456 22276 50460 22332
rect 50460 22276 50516 22332
rect 50516 22276 50520 22332
rect 50456 22272 50520 22276
rect 50536 22332 50600 22336
rect 50536 22276 50540 22332
rect 50540 22276 50596 22332
rect 50596 22276 50600 22332
rect 50536 22272 50600 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 50296 21244 50360 21248
rect 50296 21188 50300 21244
rect 50300 21188 50356 21244
rect 50356 21188 50360 21244
rect 50296 21184 50360 21188
rect 50376 21244 50440 21248
rect 50376 21188 50380 21244
rect 50380 21188 50436 21244
rect 50436 21188 50440 21244
rect 50376 21184 50440 21188
rect 50456 21244 50520 21248
rect 50456 21188 50460 21244
rect 50460 21188 50516 21244
rect 50516 21188 50520 21244
rect 50456 21184 50520 21188
rect 50536 21244 50600 21248
rect 50536 21188 50540 21244
rect 50540 21188 50596 21244
rect 50596 21188 50600 21244
rect 50536 21184 50600 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 50296 20156 50360 20160
rect 50296 20100 50300 20156
rect 50300 20100 50356 20156
rect 50356 20100 50360 20156
rect 50296 20096 50360 20100
rect 50376 20156 50440 20160
rect 50376 20100 50380 20156
rect 50380 20100 50436 20156
rect 50436 20100 50440 20156
rect 50376 20096 50440 20100
rect 50456 20156 50520 20160
rect 50456 20100 50460 20156
rect 50460 20100 50516 20156
rect 50516 20100 50520 20156
rect 50456 20096 50520 20100
rect 50536 20156 50600 20160
rect 50536 20100 50540 20156
rect 50540 20100 50596 20156
rect 50596 20100 50600 20156
rect 50536 20096 50600 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 50296 19068 50360 19072
rect 50296 19012 50300 19068
rect 50300 19012 50356 19068
rect 50356 19012 50360 19068
rect 50296 19008 50360 19012
rect 50376 19068 50440 19072
rect 50376 19012 50380 19068
rect 50380 19012 50436 19068
rect 50436 19012 50440 19068
rect 50376 19008 50440 19012
rect 50456 19068 50520 19072
rect 50456 19012 50460 19068
rect 50460 19012 50516 19068
rect 50516 19012 50520 19068
rect 50456 19008 50520 19012
rect 50536 19068 50600 19072
rect 50536 19012 50540 19068
rect 50540 19012 50596 19068
rect 50596 19012 50600 19068
rect 50536 19008 50600 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 50296 17980 50360 17984
rect 50296 17924 50300 17980
rect 50300 17924 50356 17980
rect 50356 17924 50360 17980
rect 50296 17920 50360 17924
rect 50376 17980 50440 17984
rect 50376 17924 50380 17980
rect 50380 17924 50436 17980
rect 50436 17924 50440 17980
rect 50376 17920 50440 17924
rect 50456 17980 50520 17984
rect 50456 17924 50460 17980
rect 50460 17924 50516 17980
rect 50516 17924 50520 17980
rect 50456 17920 50520 17924
rect 50536 17980 50600 17984
rect 50536 17924 50540 17980
rect 50540 17924 50596 17980
rect 50596 17924 50600 17980
rect 50536 17920 50600 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 50296 16892 50360 16896
rect 50296 16836 50300 16892
rect 50300 16836 50356 16892
rect 50356 16836 50360 16892
rect 50296 16832 50360 16836
rect 50376 16892 50440 16896
rect 50376 16836 50380 16892
rect 50380 16836 50436 16892
rect 50436 16836 50440 16892
rect 50376 16832 50440 16836
rect 50456 16892 50520 16896
rect 50456 16836 50460 16892
rect 50460 16836 50516 16892
rect 50516 16836 50520 16892
rect 50456 16832 50520 16836
rect 50536 16892 50600 16896
rect 50536 16836 50540 16892
rect 50540 16836 50596 16892
rect 50596 16836 50600 16892
rect 50536 16832 50600 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 50296 15804 50360 15808
rect 50296 15748 50300 15804
rect 50300 15748 50356 15804
rect 50356 15748 50360 15804
rect 50296 15744 50360 15748
rect 50376 15804 50440 15808
rect 50376 15748 50380 15804
rect 50380 15748 50436 15804
rect 50436 15748 50440 15804
rect 50376 15744 50440 15748
rect 50456 15804 50520 15808
rect 50456 15748 50460 15804
rect 50460 15748 50516 15804
rect 50516 15748 50520 15804
rect 50456 15744 50520 15748
rect 50536 15804 50600 15808
rect 50536 15748 50540 15804
rect 50540 15748 50596 15804
rect 50596 15748 50600 15804
rect 50536 15744 50600 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 50296 14716 50360 14720
rect 50296 14660 50300 14716
rect 50300 14660 50356 14716
rect 50356 14660 50360 14716
rect 50296 14656 50360 14660
rect 50376 14716 50440 14720
rect 50376 14660 50380 14716
rect 50380 14660 50436 14716
rect 50436 14660 50440 14716
rect 50376 14656 50440 14660
rect 50456 14716 50520 14720
rect 50456 14660 50460 14716
rect 50460 14660 50516 14716
rect 50516 14660 50520 14716
rect 50456 14656 50520 14660
rect 50536 14716 50600 14720
rect 50536 14660 50540 14716
rect 50540 14660 50596 14716
rect 50596 14660 50600 14716
rect 50536 14656 50600 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 50296 13628 50360 13632
rect 50296 13572 50300 13628
rect 50300 13572 50356 13628
rect 50356 13572 50360 13628
rect 50296 13568 50360 13572
rect 50376 13628 50440 13632
rect 50376 13572 50380 13628
rect 50380 13572 50436 13628
rect 50436 13572 50440 13628
rect 50376 13568 50440 13572
rect 50456 13628 50520 13632
rect 50456 13572 50460 13628
rect 50460 13572 50516 13628
rect 50516 13572 50520 13628
rect 50456 13568 50520 13572
rect 50536 13628 50600 13632
rect 50536 13572 50540 13628
rect 50540 13572 50596 13628
rect 50596 13572 50600 13628
rect 50536 13568 50600 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 50296 12540 50360 12544
rect 50296 12484 50300 12540
rect 50300 12484 50356 12540
rect 50356 12484 50360 12540
rect 50296 12480 50360 12484
rect 50376 12540 50440 12544
rect 50376 12484 50380 12540
rect 50380 12484 50436 12540
rect 50436 12484 50440 12540
rect 50376 12480 50440 12484
rect 50456 12540 50520 12544
rect 50456 12484 50460 12540
rect 50460 12484 50516 12540
rect 50516 12484 50520 12540
rect 50456 12480 50520 12484
rect 50536 12540 50600 12544
rect 50536 12484 50540 12540
rect 50540 12484 50596 12540
rect 50596 12484 50600 12540
rect 50536 12480 50600 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 50296 11452 50360 11456
rect 50296 11396 50300 11452
rect 50300 11396 50356 11452
rect 50356 11396 50360 11452
rect 50296 11392 50360 11396
rect 50376 11452 50440 11456
rect 50376 11396 50380 11452
rect 50380 11396 50436 11452
rect 50436 11396 50440 11452
rect 50376 11392 50440 11396
rect 50456 11452 50520 11456
rect 50456 11396 50460 11452
rect 50460 11396 50516 11452
rect 50516 11396 50520 11452
rect 50456 11392 50520 11396
rect 50536 11452 50600 11456
rect 50536 11396 50540 11452
rect 50540 11396 50596 11452
rect 50596 11396 50600 11452
rect 50536 11392 50600 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 50296 10364 50360 10368
rect 50296 10308 50300 10364
rect 50300 10308 50356 10364
rect 50356 10308 50360 10364
rect 50296 10304 50360 10308
rect 50376 10364 50440 10368
rect 50376 10308 50380 10364
rect 50380 10308 50436 10364
rect 50436 10308 50440 10364
rect 50376 10304 50440 10308
rect 50456 10364 50520 10368
rect 50456 10308 50460 10364
rect 50460 10308 50516 10364
rect 50516 10308 50520 10364
rect 50456 10304 50520 10308
rect 50536 10364 50600 10368
rect 50536 10308 50540 10364
rect 50540 10308 50596 10364
rect 50596 10308 50600 10364
rect 50536 10304 50600 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 50296 9276 50360 9280
rect 50296 9220 50300 9276
rect 50300 9220 50356 9276
rect 50356 9220 50360 9276
rect 50296 9216 50360 9220
rect 50376 9276 50440 9280
rect 50376 9220 50380 9276
rect 50380 9220 50436 9276
rect 50436 9220 50440 9276
rect 50376 9216 50440 9220
rect 50456 9276 50520 9280
rect 50456 9220 50460 9276
rect 50460 9220 50516 9276
rect 50516 9220 50520 9276
rect 50456 9216 50520 9220
rect 50536 9276 50600 9280
rect 50536 9220 50540 9276
rect 50540 9220 50596 9276
rect 50596 9220 50600 9276
rect 50536 9216 50600 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 50296 8188 50360 8192
rect 50296 8132 50300 8188
rect 50300 8132 50356 8188
rect 50356 8132 50360 8188
rect 50296 8128 50360 8132
rect 50376 8188 50440 8192
rect 50376 8132 50380 8188
rect 50380 8132 50436 8188
rect 50436 8132 50440 8188
rect 50376 8128 50440 8132
rect 50456 8188 50520 8192
rect 50456 8132 50460 8188
rect 50460 8132 50516 8188
rect 50516 8132 50520 8188
rect 50456 8128 50520 8132
rect 50536 8188 50600 8192
rect 50536 8132 50540 8188
rect 50540 8132 50596 8188
rect 50596 8132 50600 8188
rect 50536 8128 50600 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 50296 7100 50360 7104
rect 50296 7044 50300 7100
rect 50300 7044 50356 7100
rect 50356 7044 50360 7100
rect 50296 7040 50360 7044
rect 50376 7100 50440 7104
rect 50376 7044 50380 7100
rect 50380 7044 50436 7100
rect 50436 7044 50440 7100
rect 50376 7040 50440 7044
rect 50456 7100 50520 7104
rect 50456 7044 50460 7100
rect 50460 7044 50516 7100
rect 50516 7044 50520 7100
rect 50456 7040 50520 7044
rect 50536 7100 50600 7104
rect 50536 7044 50540 7100
rect 50540 7044 50596 7100
rect 50596 7044 50600 7100
rect 50536 7040 50600 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 50296 6012 50360 6016
rect 50296 5956 50300 6012
rect 50300 5956 50356 6012
rect 50356 5956 50360 6012
rect 50296 5952 50360 5956
rect 50376 6012 50440 6016
rect 50376 5956 50380 6012
rect 50380 5956 50436 6012
rect 50436 5956 50440 6012
rect 50376 5952 50440 5956
rect 50456 6012 50520 6016
rect 50456 5956 50460 6012
rect 50460 5956 50516 6012
rect 50516 5956 50520 6012
rect 50456 5952 50520 5956
rect 50536 6012 50600 6016
rect 50536 5956 50540 6012
rect 50540 5956 50596 6012
rect 50596 5956 50600 6012
rect 50536 5952 50600 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 50296 4924 50360 4928
rect 50296 4868 50300 4924
rect 50300 4868 50356 4924
rect 50356 4868 50360 4924
rect 50296 4864 50360 4868
rect 50376 4924 50440 4928
rect 50376 4868 50380 4924
rect 50380 4868 50436 4924
rect 50436 4868 50440 4924
rect 50376 4864 50440 4868
rect 50456 4924 50520 4928
rect 50456 4868 50460 4924
rect 50460 4868 50516 4924
rect 50516 4868 50520 4924
rect 50456 4864 50520 4868
rect 50536 4924 50600 4928
rect 50536 4868 50540 4924
rect 50540 4868 50596 4924
rect 50596 4868 50600 4924
rect 50536 4864 50600 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 50296 3836 50360 3840
rect 50296 3780 50300 3836
rect 50300 3780 50356 3836
rect 50356 3780 50360 3836
rect 50296 3776 50360 3780
rect 50376 3836 50440 3840
rect 50376 3780 50380 3836
rect 50380 3780 50436 3836
rect 50436 3780 50440 3836
rect 50376 3776 50440 3780
rect 50456 3836 50520 3840
rect 50456 3780 50460 3836
rect 50460 3780 50516 3836
rect 50516 3780 50520 3836
rect 50456 3776 50520 3780
rect 50536 3836 50600 3840
rect 50536 3780 50540 3836
rect 50540 3780 50596 3836
rect 50596 3780 50600 3836
rect 50536 3776 50600 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 50296 2748 50360 2752
rect 50296 2692 50300 2748
rect 50300 2692 50356 2748
rect 50356 2692 50360 2748
rect 50296 2688 50360 2692
rect 50376 2748 50440 2752
rect 50376 2692 50380 2748
rect 50380 2692 50436 2748
rect 50436 2692 50440 2748
rect 50376 2688 50440 2692
rect 50456 2748 50520 2752
rect 50456 2692 50460 2748
rect 50460 2692 50516 2748
rect 50516 2692 50520 2748
rect 50456 2688 50520 2692
rect 50536 2748 50600 2752
rect 50536 2692 50540 2748
rect 50540 2692 50596 2748
rect 50596 2692 50600 2748
rect 50536 2688 50600 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 57696 4528 57712
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 57664
rect 5528 2176 5848 57664
rect 6188 2176 6508 57664
rect 19568 57152 19888 57712
rect 34928 57696 35248 57712
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 57664
rect 20888 2176 21208 57664
rect 21548 2176 21868 57664
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 57664
rect 36248 2176 36568 57664
rect 36908 2176 37228 57664
rect 50288 57152 50608 57712
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 56064 50608 57088
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 54976 50608 56000
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 53888 50608 54912
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 52800 50608 53824
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 51712 50608 52736
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 50624 50608 51648
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 49536 50608 50560
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 48448 50608 49472
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 47360 50608 48384
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 46272 50608 47296
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 45184 50608 46208
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 44096 50608 45120
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 28864 50608 29888
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 27776 50608 28800
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 26688 50608 27712
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 25600 50608 26624
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 24512 50608 25536
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 23424 50608 24448
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 22336 50608 23360
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 21248 50608 22272
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 20160 50608 21184
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 19072 50608 20096
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 17984 50608 19008
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 16896 50608 17920
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 15808 50608 16832
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 14720 50608 15744
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 13632 50608 14656
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 12544 50608 13568
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 11456 50608 12480
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 10368 50608 11392
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 9280 50608 10304
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 8192 50608 9216
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 7104 50608 8128
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 6016 50608 7040
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 4928 50608 5952
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 3840 50608 4864
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 2752 50608 3776
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 34928 2128 35248 2144
rect 50288 2128 50608 2688
rect 50948 2176 51268 57664
rect 51608 2176 51928 57664
rect 52268 2176 52588 57664
use sky130_fd_sc_hd__decap_3  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1621523292
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1621523292
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1656 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 2668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1932 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output288 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 2760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1207_
timestamp 1621523292
transform 1 0 2760 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp 1621523292
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1621523292
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28
timestamp 1621523292
transform 1 0 3680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3128 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output310
timestamp 1621523292
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1621523292
transform 1 0 4232 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1206_
timestamp 1621523292
transform 1 0 4232 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4600 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1621523292
transform 1 0 4876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1621523292
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1621523292
transform 1 0 5520 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49
timestamp 1621523292
transform 1 0 5612 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1052_
timestamp 1621523292
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1045_
timestamp 1621523292
transform 1 0 5336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1621523292
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1621523292
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1621523292
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1621523292
transform 1 0 6348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1621523292
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1621523292
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1621523292
transform 1 0 7084 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1621523292
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1621523292
transform 1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66
timestamp 1621523292
transform 1 0 7176 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1621523292
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1621523292
transform 1 0 7544 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1621523292
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80
timestamp 1621523292
transform 1 0 8464 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1621523292
transform 1 0 8832 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1621523292
transform 1 0 8188 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1621523292
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_87 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_72
timestamp 1621523292
transform 1 0 7728 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1621523292
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1621523292
transform 1 0 10764 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88
timestamp 1621523292
transform 1 0 9200 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 1621523292
transform 1 0 10028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_108
timestamp 1621523292
transform 1 0 11040 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_99
timestamp 1621523292
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_111
timestamp 1621523292
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1621523292
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1621523292
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1621523292
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1621523292
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1621523292
transform 1 0 12512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1621523292
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1621523292
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1621523292
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1621523292
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1621523292
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1621523292
transform 1 0 13524 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1621523292
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_138
timestamp 1621523292
transform 1 0 13800 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1621523292
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1621523292
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1621523292
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1621523292
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1621523292
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_160
timestamp 1621523292
transform 1 0 15824 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1621523292
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1621523292
transform 1 0 15548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1621523292
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1621523292
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1621523292
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1621523292
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1621523292
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1621523292
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1621523292
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1621523292
transform 1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1621523292
transform 1 0 19136 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1621523292
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1621523292
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1621523292
transform 1 0 18492 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1621523292
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1621523292
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1621523292
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1621523292
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1621523292
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1621523292
transform 1 0 21068 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1621523292
transform 1 0 19412 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1621523292
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1621523292
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1621523292
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_220
timestamp 1621523292
transform 1 0 21344 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1621523292
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_224
timestamp 1621523292
transform 1 0 21712 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1621523292
transform 1 0 21344 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1621523292
transform 1 0 21804 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1621523292
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_240
timestamp 1621523292
transform 1 0 23184 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1621523292
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1621523292
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1621523292
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1621523292
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1621523292
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1621523292
transform 1 0 23828 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_246
timestamp 1621523292
transform 1 0 23736 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_250
timestamp 1621523292
transform 1 0 24104 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_258
timestamp 1621523292
transform 1 0 24840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1621523292
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_241
timestamp 1621523292
transform 1 0 23276 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1621523292
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1621523292
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1621523292
transform 1 0 26220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1621523292
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1621523292
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1621523292
transform 1 0 26496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_283
timestamp 1621523292
transform 1 0 27140 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1621523292
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_277
timestamp 1621523292
transform 1 0 26588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1621523292
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1621523292
transform 1 0 27692 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1621523292
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1621523292
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_302
timestamp 1621523292
transform 1 0 28888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_298
timestamp 1621523292
transform 1 0 28520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_302
timestamp 1621523292
transform 1 0 28888 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1621523292
transform 1 0 28520 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output266
timestamp 1621523292
transform 1 0 28980 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1621523292
transform 1 0 28244 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 28612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_286
timestamp 1621523292
transform 1 0 27416 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_309
timestamp 1621523292
transform 1 0 29532 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_307
timestamp 1621523292
transform 1 0 29348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output255
timestamp 1621523292
transform 1 0 29716 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1238_
timestamp 1621523292
transform 1 0 29900 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1051_
timestamp 1621523292
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_321
timestamp 1621523292
transform 1 0 30636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1621523292
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_315
timestamp 1621523292
transform 1 0 30084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1621523292
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_325
timestamp 1621523292
transform 1 0 31004 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1239_
timestamp 1621523292
transform 1 0 30912 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1008_
timestamp 1621523292
transform 1 0 31096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_333
timestamp 1621523292
transform 1 0 31740 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_329
timestamp 1621523292
transform 1 0 31372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1621523292
transform 1 0 31648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output277
timestamp 1621523292
transform 1 0 31832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1240_
timestamp 1621523292
transform 1 0 32016 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1621523292
transform 1 0 32660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_338
timestamp 1621523292
transform 1 0 32200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1621523292
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1621523292
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1621523292
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1621523292
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1004_
timestamp 1621523292
transform 1 0 33028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1241_
timestamp 1621523292
transform 1 0 33580 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1242_
timestamp 1621523292
transform 1 0 33672 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1243_
timestamp 1621523292
transform 1 0 34684 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_361
timestamp 1621523292
transform 1 0 34316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_350
timestamp 1621523292
transform 1 0 33304 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_362
timestamp 1621523292
transform 1 0 34408 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_370 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 35144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1621523292
transform 1 0 36064 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1621523292
transform 1 0 35880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1621523292
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1621523292
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1244_
timestamp 1621523292
transform 1 0 35328 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1621523292
transform 1 0 36800 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output283
timestamp 1621523292
transform 1 0 36432 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1245_
timestamp 1621523292
transform 1 0 36248 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_390
timestamp 1621523292
transform 1 0 36984 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0994_
timestamp 1621523292
transform 1 0 37168 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_400
timestamp 1621523292
transform 1 0 37904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_395
timestamp 1621523292
transform 1 0 37444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output256
timestamp 1621523292
transform 1 0 37720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1621523292
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1621523292
transform 1 0 38548 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1621523292
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1621523292
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1246_
timestamp 1621523292
transform 1 0 38272 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1621523292
transform 1 0 39008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1247_
timestamp 1621523292
transform 1 0 38916 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_419
timestamp 1621523292
transform 1 0 39652 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_419
timestamp 1621523292
transform 1 0 39652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1249_
timestamp 1621523292
transform 1 0 40020 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1248_
timestamp 1621523292
transform 1 0 40020 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0996_
timestamp 1621523292
transform 1 0 39376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1621523292
transform 1 0 40756 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1621523292
transform 1 0 40756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_436
timestamp 1621523292
transform 1 0 41216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output257
timestamp 1621523292
transform 1 0 41124 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1621523292
transform 1 0 41124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1250_
timestamp 1621523292
transform 1 0 41584 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1251_
timestamp 1621523292
transform 1 0 42688 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1621523292
transform 1 0 43056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output258
timestamp 1621523292
transform 1 0 41860 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_448
timestamp 1621523292
transform 1 0 42320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_439
timestamp 1621523292
transform 1 0 41492 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_447
timestamp 1621523292
transform 1 0 42228 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_455
timestamp 1621523292
transform 1 0 42964 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1621523292
transform 1 0 43148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1252_
timestamp 1621523292
transform 1 0 43516 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1253_
timestamp 1621523292
transform 1 0 44252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1621523292
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output261
timestamp 1621523292
transform 1 0 44620 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_460
timestamp 1621523292
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_465
timestamp 1621523292
transform 1 0 43884 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1621523292
transform 1 0 44988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_469
timestamp 1621523292
transform 1 0 44252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_477
timestamp 1621523292
transform 1 0 44988 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _1254_
timestamp 1621523292
transform 1 0 45356 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1255_
timestamp 1621523292
transform 1 0 45540 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1256_
timestamp 1621523292
transform 1 0 46920 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1257_
timestamp 1621523292
transform 1 0 47196 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1621523292
transform 1 0 46460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1621523292
transform 1 0 46092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1621523292
transform 1 0 46552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_491
timestamp 1621523292
transform 1 0 46276 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_499
timestamp 1621523292
transform 1 0 47012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1258_
timestamp 1621523292
transform 1 0 48760 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1621523292
transform 1 0 49128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1621523292
transform 1 0 48300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output260
timestamp 1621523292
transform 1 0 48024 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_506
timestamp 1621523292
transform 1 0 47656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_514
timestamp 1621523292
transform 1 0 48392 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_523
timestamp 1621523292
transform 1 0 49220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_509
timestamp 1621523292
transform 1 0 47932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_514
timestamp 1621523292
transform 1 0 48392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1259_
timestamp 1621523292
transform 1 0 49588 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1260_
timestamp 1621523292
transform 1 0 50692 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output267
timestamp 1621523292
transform 1 0 49864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output268
timestamp 1621523292
transform 1 0 50600 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_535
timestamp 1621523292
transform 1 0 50324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_526
timestamp 1621523292
transform 1 0 49496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_534
timestamp 1621523292
transform 1 0 50232 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_542
timestamp 1621523292
transform 1 0 50968 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_550
timestamp 1621523292
transform 1 0 51704 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_552
timestamp 1621523292
transform 1 0 51888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_547
timestamp 1621523292
transform 1 0 51428 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output269
timestamp 1621523292
transform 1 0 51336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1621523292
transform 1 0 51796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_556
timestamp 1621523292
transform 1 0 52256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1262_
timestamp 1621523292
transform 1 0 52348 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1261_
timestamp 1621523292
transform 1 0 52256 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_565
timestamp 1621523292
transform 1 0 53084 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1621523292
transform 1 0 52992 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1621523292
transform 1 0 53636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_569
timestamp 1621523292
transform 1 0 53452 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_576
timestamp 1621523292
transform 1 0 54096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output272
timestamp 1621523292
transform 1 0 54004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1621523292
transform 1 0 53544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1263_
timestamp 1621523292
transform 1 0 53360 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_579
timestamp 1621523292
transform 1 0 54372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_581
timestamp 1621523292
transform 1 0 54556 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 54740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output273
timestamp 1621523292
transform 1 0 54740 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1621523292
transform 1 0 54464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1265_
timestamp 1621523292
transform 1 0 54924 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_587
timestamp 1621523292
transform 1 0 55108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1266_
timestamp 1621523292
transform 1 0 55568 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1267_
timestamp 1621523292
transform 1 0 56028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1269_
timestamp 1621523292
transform 1 0 56856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1621523292
transform 1 0 57132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1621523292
transform 1 0 55660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_605
timestamp 1621523292
transform 1 0 56764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_610
timestamp 1621523292
transform 1 0 57224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_591
timestamp 1621523292
transform 1 0 55476 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_600
timestamp 1621523292
transform 1 0 56304 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0922_
timestamp 1621523292
transform 1 0 57960 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1621523292
transform -1 0 58880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1621523292
transform -1 0 58880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output176
timestamp 1621523292
transform 1 0 57868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_616
timestamp 1621523292
transform 1 0 57776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1621523292
transform 1 0 58236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_614
timestamp 1621523292
transform 1 0 57592 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1621523292
transform 1 0 58236 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1209_
timestamp 1621523292
transform 1 0 1932 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1621523292
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output299
timestamp 1621523292
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1621523292
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1621523292
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1093_
timestamp 1621523292
transform 1 0 4232 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1095_
timestamp 1621523292
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1621523292
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1621523292
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_30
timestamp 1621523292
transform 1 0 3864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1621523292
transform 1 0 4508 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1621523292
transform 1 0 5520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1621523292
transform 1 0 6164 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_44
timestamp 1621523292
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1621523292
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_58
timestamp 1621523292
transform 1 0 6440 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1621523292
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70
timestamp 1621523292
transform 1 0 7544 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_82
timestamp 1621523292
transform 1 0 8648 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1621523292
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1621523292
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1621523292
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1621523292
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1621523292
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1621523292
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1621523292
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1621523292
transform 1 0 15456 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1621523292
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1621523292
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1621523292
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1621523292
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1621523292
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_213
timestamp 1621523292
transform 1 0 20700 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1621523292
transform 1 0 21804 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_237
timestamp 1621523292
transform 1 0 22908 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1621523292
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_249
timestamp 1621523292
transform 1 0 24012 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1621523292
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_270
timestamp 1621523292
transform 1 0 25944 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_282
timestamp 1621523292
transform 1 0 27048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1621523292
transform 1 0 28520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1621523292
transform 1 0 28152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1621523292
transform 1 0 28796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1009_
timestamp 1621523292
transform 1 0 30544 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1126_
timestamp 1621523292
transform 1 0 31188 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1621523292
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1621523292
transform 1 0 29348 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_310
timestamp 1621523292
transform 1 0 29624 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1621523292
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_319
timestamp 1621523292
transform 1 0 30452 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_323
timestamp 1621523292
transform 1 0 30820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1127_
timestamp 1621523292
transform 1 0 31832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1128_
timestamp 1621523292
transform 1 0 32568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1621523292
transform 1 0 33212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_330
timestamp 1621523292
transform 1 0 31464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_337
timestamp 1621523292
transform 1 0 32108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_341
timestamp 1621523292
transform 1 0 32476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_345
timestamp 1621523292
transform 1 0 32844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1621523292
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output281
timestamp 1621523292
transform 1 0 34132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_353
timestamp 1621523292
transform 1 0 33580 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_363
timestamp 1621523292
transform 1 0 34500 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output282
timestamp 1621523292
transform 1 0 35696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output284
timestamp 1621523292
transform 1 0 36984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1621523292
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_380
timestamp 1621523292
transform 1 0 36064 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_388
timestamp 1621523292
transform 1 0 36800 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output285
timestamp 1621523292
transform 1 0 37904 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output286
timestamp 1621523292
transform 1 0 38824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_394
timestamp 1621523292
transform 1 0 37352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_404
timestamp 1621523292
transform 1 0 38272 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_414
timestamp 1621523292
transform 1 0 39192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0995_
timestamp 1621523292
transform 1 0 40940 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0997_
timestamp 1621523292
transform 1 0 39560 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1621523292
transform 1 0 40480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_421
timestamp 1621523292
transform 1 0 39836 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_427
timestamp 1621523292
transform 1 0 40388 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1621523292
transform 1 0 40572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_436
timestamp 1621523292
transform 1 0 41216 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0992_
timestamp 1621523292
transform 1 0 41952 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output259
timestamp 1621523292
transform 1 0 42596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1621523292
transform 1 0 42228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_455
timestamp 1621523292
transform 1 0 42964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0985_
timestamp 1621523292
transform 1 0 45080 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0988_
timestamp 1621523292
transform 1 0 43332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0990_
timestamp 1621523292
transform 1 0 44436 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_462
timestamp 1621523292
transform 1 0 43608 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_470
timestamp 1621523292
transform 1 0 44344 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_474
timestamp 1621523292
transform 1 0 44712 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1621523292
transform 1 0 45724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output262
timestamp 1621523292
transform 1 0 46184 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output263
timestamp 1621523292
transform 1 0 46920 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_481
timestamp 1621523292
transform 1 0 45356 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_486
timestamp 1621523292
transform 1 0 45816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1621523292
transform 1 0 46552 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_502
timestamp 1621523292
transform 1 0 47288 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output264
timestamp 1621523292
transform 1 0 47656 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output265
timestamp 1621523292
transform 1 0 48392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1621523292
transform 1 0 48024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_518
timestamp 1621523292
transform 1 0 48760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0971_
timestamp 1621523292
transform 1 0 49588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0975_
timestamp 1621523292
transform 1 0 50232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1621523292
transform 1 0 50968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_526
timestamp 1621523292
transform 1 0 49496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_530
timestamp 1621523292
transform 1 0 49864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1621523292
transform 1 0 50600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_543
timestamp 1621523292
transform 1 0 51060 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output270
timestamp 1621523292
transform 1 0 51980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output271
timestamp 1621523292
transform 1 0 52900 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_551
timestamp 1621523292
transform 1 0 51796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_557
timestamp 1621523292
transform 1 0 52348 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_567
timestamp 1621523292
transform 1 0 53268 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0923_
timestamp 1621523292
transform 1 0 54832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1264_
timestamp 1621523292
transform 1 0 53728 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_571
timestamp 1621523292
transform 1 0 53636 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_580
timestamp 1621523292
transform 1 0 54464 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_587
timestamp 1621523292
transform 1 0 55108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1621523292
transform 1 0 56212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output214
timestamp 1621523292
transform 1 0 56764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output225
timestamp 1621523292
transform 1 0 55476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1621523292
transform 1 0 57316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_595
timestamp 1621523292
transform 1 0 55844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_600
timestamp 1621523292
transform 1 0 56304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_604
timestamp 1621523292
transform 1 0 56672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_609
timestamp 1621523292
transform 1 0 57132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1308_
timestamp 1621523292
transform 1 0 57500 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1621523292
transform -1 0 58880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1621523292
transform 1 0 58236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1210_
timestamp 1621523292
transform 1 0 1564 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1621523292
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output314
timestamp 1621523292
transform 1 0 2668 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1621523292
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1621523292
transform 1 0 2300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1621523292
transform 1 0 3036 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1621523292
transform 1 0 3404 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1094_
timestamp 1621523292
transform 1 0 4048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1621523292
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1621523292
transform 1 0 3680 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1621523292
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1621523292
transform 1 0 4968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1621523292
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_54
timestamp 1621523292
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1621523292
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1621523292
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1621523292
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1621523292
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1621523292
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1621523292
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1621523292
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1621523292
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1621523292
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1621523292
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1621523292
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1621523292
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1621523292
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1621523292
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1621523292
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1621523292
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1621523292
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_220
timestamp 1621523292
transform 1 0 21344 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_229
timestamp 1621523292
transform 1 0 22172 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_241
timestamp 1621523292
transform 1 0 23276 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1621523292
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1621523292
transform 1 0 25484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_277
timestamp 1621523292
transform 1 0 26588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1621523292
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_286
timestamp 1621523292
transform 1 0 27416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_298
timestamp 1621523292
transform 1 0 28520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_310
timestamp 1621523292
transform 1 0 29624 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_322
timestamp 1621523292
transform 1 0 30728 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1005_
timestamp 1621523292
transform 1 0 33120 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1621523292
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_334
timestamp 1621523292
transform 1 0 31832 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_343
timestamp 1621523292
transform 1 0 32660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_347
timestamp 1621523292
transform 1 0 33028 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1003_
timestamp 1621523292
transform 1 0 34408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1129_
timestamp 1621523292
transform 1 0 33764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_351
timestamp 1621523292
transform 1 0 33396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_358
timestamp 1621523292
transform 1 0 34040 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_365
timestamp 1621523292
transform 1 0 34684 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1000_
timestamp 1621523292
transform 1 0 36800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1001_
timestamp 1621523292
transform 1 0 36156 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1002_
timestamp 1621523292
transform 1 0 35512 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_373
timestamp 1621523292
transform 1 0 35420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_377
timestamp 1621523292
transform 1 0 35788 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_384
timestamp 1621523292
transform 1 0 36432 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_391
timestamp 1621523292
transform 1 0 37076 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0998_
timestamp 1621523292
transform 1 0 38272 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1133_
timestamp 1621523292
transform 1 0 38916 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1621523292
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_400
timestamp 1621523292
transform 1 0 37904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_407
timestamp 1621523292
transform 1 0 38548 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_414
timestamp 1621523292
transform 1 0 39192 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1135_
timestamp 1621523292
transform 1 0 39560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1136_
timestamp 1621523292
transform 1 0 40296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1137_
timestamp 1621523292
transform 1 0 40940 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_421
timestamp 1621523292
transform 1 0 39836 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_425
timestamp 1621523292
transform 1 0 40204 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_429
timestamp 1621523292
transform 1 0 40572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_436
timestamp 1621523292
transform 1 0 41216 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0993_
timestamp 1621523292
transform 1 0 42412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1138_
timestamp 1621523292
transform 1 0 41768 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1621523292
transform 1 0 43056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_445
timestamp 1621523292
transform 1 0 42044 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_452
timestamp 1621523292
transform 1 0 42688 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_457
timestamp 1621523292
transform 1 0 43148 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0989_
timestamp 1621523292
transform 1 0 45080 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0991_
timestamp 1621523292
transform 1 0 43976 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_465
timestamp 1621523292
transform 1 0 43884 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_469
timestamp 1621523292
transform 1 0 44252 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_477
timestamp 1621523292
transform 1 0 44988 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0979_
timestamp 1621523292
transform 1 0 47012 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0982_
timestamp 1621523292
transform 1 0 46368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0987_
timestamp 1621523292
transform 1 0 45724 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_481
timestamp 1621523292
transform 1 0 45356 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_488
timestamp 1621523292
transform 1 0 46000 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_495
timestamp 1621523292
transform 1 0 46644 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_502
timestamp 1621523292
transform 1 0 47288 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0973_
timestamp 1621523292
transform 1 0 48944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0977_
timestamp 1621523292
transform 1 0 47656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1621523292
transform 1 0 48300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_509
timestamp 1621523292
transform 1 0 47932 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_514
timestamp 1621523292
transform 1 0 48392 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_523
timestamp 1621523292
transform 1 0 49220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1621523292
transform 1 0 50876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0970_
timestamp 1621523292
transform 1 0 50232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0972_
timestamp 1621523292
transform 1 0 49588 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_530
timestamp 1621523292
transform 1 0 49864 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_537
timestamp 1621523292
transform 1 0 50508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_544
timestamp 1621523292
transform 1 0 51152 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0924_
timestamp 1621523292
transform 1 0 52164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0968_
timestamp 1621523292
transform 1 0 51520 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output279
timestamp 1621523292
transform 1 0 52808 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_551
timestamp 1621523292
transform 1 0 51796 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_558
timestamp 1621523292
transform 1 0 52440 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_566
timestamp 1621523292
transform 1 0 53176 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1621523292
transform 1 0 53544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output274
timestamp 1621523292
transform 1 0 55016 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output275
timestamp 1621523292
transform 1 0 54280 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_571
timestamp 1621523292
transform 1 0 53636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_577
timestamp 1621523292
transform 1 0 54188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_582
timestamp 1621523292
transform 1 0 54648 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1268_
timestamp 1621523292
transform 1 0 56488 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output236
timestamp 1621523292
transform 1 0 55752 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1621523292
transform 1 0 56304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1621523292
transform 1 0 55384 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_598
timestamp 1621523292
transform 1 0 56120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_610
timestamp 1621523292
transform 1 0 57224 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1621523292
transform -1 0 58880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output187
timestamp 1621523292
transform 1 0 57868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_616
timestamp 1621523292
transform 1 0 57776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1621523292
transform 1 0 58236 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1042_
timestamp 1621523292
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1211_
timestamp 1621523292
transform 1 0 1932 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1621523292
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1621523292
transform 1 0 1380 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1621523292
transform 1 0 2668 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1097_
timestamp 1621523292
transform 1 0 4232 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1621523292
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1621523292
transform 1 0 3312 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1621523292
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_30
timestamp 1621523292
transform 1 0 3864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_37
timestamp 1621523292
transform 1 0 4508 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_49
timestamp 1621523292
transform 1 0 5612 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_61
timestamp 1621523292
transform 1 0 6716 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1621523292
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_73
timestamp 1621523292
transform 1 0 7820 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1621523292
transform 1 0 8924 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1621523292
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1621523292
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1621523292
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1621523292
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1621523292
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1621523292
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1621523292
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1621523292
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1621523292
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1621523292
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1621523292
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1621523292
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1621523292
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_213
timestamp 1621523292
transform 1 0 20700 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1621523292
transform 1 0 21804 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1621523292
transform 1 0 22908 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1621523292
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_249
timestamp 1621523292
transform 1 0 24012 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1621523292
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_270
timestamp 1621523292
transform 1 0 25944 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_282
timestamp 1621523292
transform 1 0 27048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_294
timestamp 1621523292
transform 1 0 28152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1621523292
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_306
timestamp 1621523292
transform 1 0 29256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_315
timestamp 1621523292
transform 1 0 30084 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_327
timestamp 1621523292
transform 1 0 31188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_339
timestamp 1621523292
transform 1 0 32292 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1130_
timestamp 1621523292
transform 1 0 34316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1621523292
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_351
timestamp 1621523292
transform 1 0 33396 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_359
timestamp 1621523292
transform 1 0 34132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_364
timestamp 1621523292
transform 1 0 34592 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_370
timestamp 1621523292
transform 1 0 35144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1131_
timestamp 1621523292
transform 1 0 35696 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1132_
timestamp 1621523292
transform 1 0 36524 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_372
timestamp 1621523292
transform 1 0 35328 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_379
timestamp 1621523292
transform 1 0 35972 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_388
timestamp 1621523292
transform 1 0 36800 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0999_
timestamp 1621523292
transform 1 0 37904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1134_
timestamp 1621523292
transform 1 0 38548 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1621523292
transform 1 0 38180 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_410
timestamp 1621523292
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1621523292
transform 1 0 40480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_422
timestamp 1621523292
transform 1 0 39928 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_429
timestamp 1621523292
transform 1 0 40572 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1139_
timestamp 1621523292
transform 1 0 42596 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_441
timestamp 1621523292
transform 1 0 41676 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_449
timestamp 1621523292
transform 1 0 42412 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_454
timestamp 1621523292
transform 1 0 42872 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_458
timestamp 1621523292
transform 1 0 43240 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1140_
timestamp 1621523292
transform 1 0 43976 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1141_
timestamp 1621523292
transform 1 0 44896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1156_
timestamp 1621523292
transform 1 0 43332 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_462
timestamp 1621523292
transform 1 0 43608 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1621523292
transform 1 0 44252 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1621523292
transform 1 0 44804 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_479
timestamp 1621523292
transform 1 0 45172 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0981_
timestamp 1621523292
transform 1 0 47288 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0986_
timestamp 1621523292
transform 1 0 46644 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1621523292
transform 1 0 45724 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_486
timestamp 1621523292
transform 1 0 45816 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_494
timestamp 1621523292
transform 1 0 46552 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_498
timestamp 1621523292
transform 1 0 46920 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0974_
timestamp 1621523292
transform 1 0 49220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0976_
timestamp 1621523292
transform 1 0 48576 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0978_
timestamp 1621523292
transform 1 0 47932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_505
timestamp 1621523292
transform 1 0 47564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1621523292
transform 1 0 48208 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_519
timestamp 1621523292
transform 1 0 48852 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0653_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 49864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1621523292
transform 1 0 50968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_526
timestamp 1621523292
transform 1 0 49496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_533
timestamp 1621523292
transform 1 0 50140 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_541
timestamp 1621523292
transform 1 0 50876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_543
timestamp 1621523292
transform 1 0 51060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1351_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51520 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_547
timestamp 1621523292
transform 1 0 51428 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_564
timestamp 1621523292
transform 1 0 52992 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0944_
timestamp 1621523292
transform 1 0 55200 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1621523292
transform 1 0 53360 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_4_584
timestamp 1621523292
transform 1 0 54832 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1621523292
transform 1 0 56212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output198
timestamp 1621523292
transform 1 0 56764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1621523292
transform 1 0 57316 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_592
timestamp 1621523292
transform 1 0 55568 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_598
timestamp 1621523292
transform 1 0 56120 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_600
timestamp 1621523292
transform 1 0 56304 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_604
timestamp 1621523292
transform 1 0 56672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_609
timestamp 1621523292
transform 1 0 57132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1309_
timestamp 1621523292
transform 1 0 57500 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1621523292
transform -1 0 58880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1621523292
transform 1 0 58236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1621523292
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output313
timestamp 1621523292
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output315
timestamp 1621523292
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1621523292
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1621523292
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_19
timestamp 1621523292
transform 1 0 2852 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1621523292
transform 1 0 3220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1096_
timestamp 1621523292
transform 1 0 3864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1621523292
transform 1 0 3496 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_33
timestamp 1621523292
transform 1 0 4140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1621523292
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_45
timestamp 1621523292
transform 1 0 5244 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1621523292
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1621523292
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1621523292
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1621523292
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1621523292
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1621523292
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1621523292
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1621523292
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1621523292
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1621523292
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1621523292
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1621523292
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1621523292
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1621523292
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1621523292
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1621523292
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1621523292
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1621523292
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_229
timestamp 1621523292
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_241
timestamp 1621523292
transform 1 0 23276 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1621523292
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_265
timestamp 1621523292
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_277
timestamp 1621523292
transform 1 0 26588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1621523292
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_286
timestamp 1621523292
transform 1 0 27416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_298
timestamp 1621523292
transform 1 0 28520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_310
timestamp 1621523292
transform 1 0 29624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_322
timestamp 1621523292
transform 1 0 30728 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1621523292
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_334
timestamp 1621523292
transform 1 0 31832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1621523292
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_355
timestamp 1621523292
transform 1 0 33764 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1621523292
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1621523292
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_391
timestamp 1621523292
transform 1 0 37076 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1621523292
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_400
timestamp 1621523292
transform 1 0 37904 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_412
timestamp 1621523292
transform 1 0 39008 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_424
timestamp 1621523292
transform 1 0 40112 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_436
timestamp 1621523292
transform 1 0 41216 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1621523292
transform 1 0 43056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_448
timestamp 1621523292
transform 1 0 42320 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_457
timestamp 1621523292
transform 1 0 43148 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1149_
timestamp 1621523292
transform 1 0 44804 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1153_
timestamp 1621523292
transform 1 0 44160 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1621523292
transform 1 0 43516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_464
timestamp 1621523292
transform 1 0 43792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_471
timestamp 1621523292
transform 1 0 44436 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_478
timestamp 1621523292
transform 1 0 45080 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 1621523292
transform 1 0 47012 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1142_
timestamp 1621523292
transform 1 0 45448 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1143_
timestamp 1621523292
transform 1 0 46368 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_485
timestamp 1621523292
transform 1 0 45724 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_491
timestamp 1621523292
transform 1 0 46276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_495
timestamp 1621523292
transform 1 0 46644 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_502
timestamp 1621523292
transform 1 0 47288 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1621523292
transform 1 0 47656 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1621523292
transform 1 0 49312 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1621523292
transform 1 0 48300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_509
timestamp 1621523292
transform 1 0 47932 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_514
timestamp 1621523292
transform 1 0 48392 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_522
timestamp 1621523292
transform 1 0 49128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0730_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51152 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_540
timestamp 1621523292
transform 1 0 50784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0650_
timestamp 1621523292
transform 1 0 52900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0865_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_547
timestamp 1621523292
transform 1 0 51428 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_551
timestamp 1621523292
transform 1 0 51796 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_555
timestamp 1621523292
transform 1 0 52164 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_566
timestamp 1621523292
transform 1 0 53176 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1621523292
transform 1 0 54004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1621523292
transform 1 0 53544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output278
timestamp 1621523292
transform 1 0 54648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_571
timestamp 1621523292
transform 1 0 53636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_578
timestamp 1621523292
transform 1 0 54280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_586
timestamp 1621523292
transform 1 0 55016 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1271_
timestamp 1621523292
transform 1 0 55384 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output245
timestamp 1621523292
transform 1 0 56764 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1621523292
transform 1 0 57316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_598
timestamp 1621523292
transform 1 0 56120 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_604
timestamp 1621523292
transform 1 0 56672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_609
timestamp 1621523292
transform 1 0 57132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1310_
timestamp 1621523292
transform 1 0 57500 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1621523292
transform -1 0 58880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1621523292
transform 1 0 58236 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1621523292
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1621523292
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output316
timestamp 1621523292
transform 1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1621523292
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1621523292
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1212_
timestamp 1621523292
transform 1 0 1656 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1621523292
transform 1 0 2116 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1621523292
transform 1 0 2392 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1621523292
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1621523292
transform 1 0 2760 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_21
timestamp 1621523292
transform 1 0 3036 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1040_
timestamp 1621523292
transform 1 0 2760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1098_
timestamp 1621523292
transform 1 0 3128 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1099_
timestamp 1621523292
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1621523292
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1621523292
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_37
timestamp 1621523292
transform 1 0 4508 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_25
timestamp 1621523292
transform 1 0 3404 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_37
timestamp 1621523292
transform 1 0 4508 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1621523292
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_49
timestamp 1621523292
transform 1 0 5612 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_61
timestamp 1621523292
transform 1 0 6716 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_49
timestamp 1621523292
transform 1 0 5612 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1621523292
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1621523292
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_73
timestamp 1621523292
transform 1 0 7820 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1621523292
transform 1 0 8924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1621523292
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1621523292
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1621523292
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1621523292
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1621523292
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1621523292
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1621523292
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1621523292
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1621523292
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1621523292
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1621523292
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1621523292
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1621523292
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1621523292
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1621523292
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1621523292
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1621523292
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1621523292
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1621523292
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1621523292
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1621523292
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1621523292
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1621523292
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1621523292
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1621523292
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1621523292
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1621523292
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1621523292
transform 1 0 20700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1621523292
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1621523292
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1621523292
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_237
timestamp 1621523292
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_220
timestamp 1621523292
transform 1 0 21344 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1621523292
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1621523292
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_249
timestamp 1621523292
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1621523292
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_241
timestamp 1621523292
transform 1 0 23276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1621523292
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_270
timestamp 1621523292
transform 1 0 25944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1621523292
transform 1 0 27048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1621523292
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1621523292
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1621523292
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_294
timestamp 1621523292
transform 1 0 28152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1621523292
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_298
timestamp 1621523292
transform 1 0 28520 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1621523292
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_306
timestamp 1621523292
transform 1 0 29256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_315
timestamp 1621523292
transform 1 0 30084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_327
timestamp 1621523292
transform 1 0 31188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_310
timestamp 1621523292
transform 1 0 29624 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_322
timestamp 1621523292
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1621523292
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_339
timestamp 1621523292
transform 1 0 32292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_334
timestamp 1621523292
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_343
timestamp 1621523292
transform 1 0 32660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1621523292
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_351
timestamp 1621523292
transform 1 0 33396 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_363
timestamp 1621523292
transform 1 0 34500 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_355
timestamp 1621523292
transform 1 0 33764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1621523292
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_372
timestamp 1621523292
transform 1 0 35328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_384
timestamp 1621523292
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1621523292
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_391
timestamp 1621523292
transform 1 0 37076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1621523292
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_396
timestamp 1621523292
transform 1 0 37536 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_408
timestamp 1621523292
transform 1 0 38640 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_400
timestamp 1621523292
transform 1 0 37904 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_412
timestamp 1621523292
transform 1 0 39008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1621523292
transform 1 0 40480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_420
timestamp 1621523292
transform 1 0 39744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_429
timestamp 1621523292
transform 1 0 40572 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_424
timestamp 1621523292
transform 1 0 40112 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_436
timestamp 1621523292
transform 1 0 41216 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1621523292
transform 1 0 43056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_441
timestamp 1621523292
transform 1 0 41676 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_453
timestamp 1621523292
transform 1 0 42780 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_448
timestamp 1621523292
transform 1 0 42320 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_457
timestamp 1621523292
transform 1 0 43148 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_461
timestamp 1621523292
transform 1 0 43516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1621523292
transform 1 0 43792 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_469
timestamp 1621523292
transform 1 0 44252 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_467
timestamp 1621523292
transform 1 0 44068 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1621523292
transform 1 0 44252 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1621523292
transform 1 0 44436 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1166_
timestamp 1621523292
transform 1 0 44436 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_474
timestamp 1621523292
transform 1 0 44712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1621523292
transform 1 0 44712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1621523292
transform 1 0 44896 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1621523292
transform 1 0 44896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _1165_
timestamp 1621523292
transform 1 0 45080 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1152_
timestamp 1621523292
transform 1 0 45080 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_481
timestamp 1621523292
transform 1 0 45356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_481
timestamp 1621523292
transform 1 0 45356 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1621523292
transform 1 0 45540 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1621523292
transform 1 0 45724 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1155_
timestamp 1621523292
transform 1 0 45724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_488
timestamp 1621523292
transform 1 0 46000 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_490
timestamp 1621523292
transform 1 0 46184 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_486
timestamp 1621523292
transform 1 0 45816 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_494
timestamp 1621523292
transform 1 0 46552 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1150_
timestamp 1621523292
transform 1 0 46368 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1148_
timestamp 1621523292
transform 1 0 46276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_495
timestamp 1621523292
transform 1 0 46644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1146_
timestamp 1621523292
transform 1 0 47012 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1144_
timestamp 1621523292
transform 1 0 46920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_502
timestamp 1621523292
transform 1 0 47288 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_501
timestamp 1621523292
transform 1 0 47196 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1059_
timestamp 1621523292
transform 1 0 47656 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1058_
timestamp 1621523292
transform 1 0 47564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_509
timestamp 1621523292
transform 1 0 47932 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_508
timestamp 1621523292
transform 1 0 47840 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_514
timestamp 1621523292
transform 1 0 48392 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_515
timestamp 1621523292
transform 1 0 48484 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1621523292
transform 1 0 48300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1049_
timestamp 1621523292
transform 1 0 48208 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_518
timestamp 1621523292
transform 1 0 48760 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0983_
timestamp 1621523292
transform 1 0 48852 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1621523292
transform 1 0 48852 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_522
timestamp 1621523292
transform 1 0 49128 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_522
timestamp 1621523292
transform 1 0 49128 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_529
timestamp 1621523292
transform 1 0 49772 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_529
timestamp 1621523292
transform 1 0 49772 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0967_
timestamp 1621523292
transform 1 0 49496 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1621523292
transform 1 0 49496 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_536
timestamp 1621523292
transform 1 0 50416 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0732_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 50140 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0652_
timestamp 1621523292
transform 1 0 50140 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_540
timestamp 1621523292
transform 1 0 50784 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_543
timestamp 1621523292
transform 1 0 51060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1621523292
transform 1 0 50968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _0734_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51152 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52716 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0738_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52348 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_547
timestamp 1621523292
transform 1 0 51428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_556
timestamp 1621523292
transform 1 0 52256 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_560
timestamp 1621523292
transform 1 0 52624 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_551
timestamp 1621523292
transform 1 0 51796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_564
timestamp 1621523292
transform 1 0 52992 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_571
timestamp 1621523292
transform 1 0 53636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_575
timestamp 1621523292
transform 1 0 54004 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_568
timestamp 1621523292
transform 1 0 53360 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1621523292
transform 1 0 53544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1621523292
transform 1 0 53728 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0736_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 54004 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_583
timestamp 1621523292
transform 1 0 54740 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_583
timestamp 1621523292
transform 1 0 54740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_579
timestamp 1621523292
transform 1 0 54372 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1621523292
transform 1 0 54464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_587
timestamp 1621523292
transform 1 0 55108 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1621523292
transform 1 0 55200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1272_
timestamp 1621523292
transform 1 0 56672 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1273_
timestamp 1621523292
transform 1 0 56396 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1621523292
transform 1 0 56212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output276
timestamp 1621523292
transform 1 0 55476 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_595
timestamp 1621523292
transform 1 0 55844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_600
timestamp 1621523292
transform 1 0 56304 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_591
timestamp 1621523292
transform 1 0 55476 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_599
timestamp 1621523292
transform 1 0 56212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_609
timestamp 1621523292
transform 1 0 57132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1311_
timestamp 1621523292
transform 1 0 57500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1621523292
transform -1 0 58880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1621523292
transform -1 0 58880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output207
timestamp 1621523292
transform 1 0 57868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_612
timestamp 1621523292
transform 1 0 57408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_616
timestamp 1621523292
transform 1 0 57776 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1621523292
transform 1 0 58236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1621523292
transform 1 0 58236 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1100_
timestamp 1621523292
transform 1 0 2760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1213_
timestamp 1621523292
transform 1 0 1656 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1621523292
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1621523292
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_14
timestamp 1621523292
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_21
timestamp 1621523292
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1621523292
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1621523292
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1621523292
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1621523292
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1621523292
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1621523292
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1621523292
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1621523292
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1621523292
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1621523292
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1621523292
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1621523292
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1621523292
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1621523292
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1621523292
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1621523292
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1621523292
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1621523292
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1621523292
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1621523292
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_213
timestamp 1621523292
transform 1 0 20700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_225
timestamp 1621523292
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_237
timestamp 1621523292
transform 1 0 22908 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1621523292
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1621523292
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_258
timestamp 1621523292
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_270
timestamp 1621523292
transform 1 0 25944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1621523292
transform 1 0 27048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_294
timestamp 1621523292
transform 1 0 28152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1621523292
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1621523292
transform 1 0 29256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_315
timestamp 1621523292
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_327
timestamp 1621523292
transform 1 0 31188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_339
timestamp 1621523292
transform 1 0 32292 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1621523292
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_351
timestamp 1621523292
transform 1 0 33396 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_363
timestamp 1621523292
transform 1 0 34500 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1621523292
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1621523292
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_396
timestamp 1621523292
transform 1 0 37536 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_408
timestamp 1621523292
transform 1 0 38640 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1621523292
transform 1 0 40480 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_420
timestamp 1621523292
transform 1 0 39744 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_429
timestamp 1621523292
transform 1 0 40572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_441
timestamp 1621523292
transform 1 0 41676 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_453
timestamp 1621523292
transform 1 0 42780 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1621523292
transform 1 0 45080 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_465
timestamp 1621523292
transform 1 0 43884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_477
timestamp 1621523292
transform 1 0 44988 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1154_
timestamp 1621523292
transform 1 0 46736 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1621523292
transform 1 0 45724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_481
timestamp 1621523292
transform 1 0 45356 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_486
timestamp 1621523292
transform 1 0 45816 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_494
timestamp 1621523292
transform 1 0 46552 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_499
timestamp 1621523292
transform 1 0 47012 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1145_
timestamp 1621523292
transform 1 0 48024 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1147_
timestamp 1621523292
transform 1 0 47380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1350_
timestamp 1621523292
transform 1 0 48668 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_506
timestamp 1621523292
transform 1 0 47656 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_513
timestamp 1621523292
transform 1 0 48300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1621523292
transform 1 0 50968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_533
timestamp 1621523292
transform 1 0 50140 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_541
timestamp 1621523292
transform 1 0 50876 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_543
timestamp 1621523292
transform 1 0 51060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0727_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 53176 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51612 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_556
timestamp 1621523292
transform 1 0 52256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_564
timestamp 1621523292
transform 1 0 52992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1621523292
transform 1 0 54188 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_573
timestamp 1621523292
transform 1 0 53820 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1621523292
transform 1 0 56212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output246
timestamp 1621523292
transform 1 0 56764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_593
timestamp 1621523292
transform 1 0 55660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_600
timestamp 1621523292
transform 1 0 56304 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_604
timestamp 1621523292
transform 1 0 56672 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_609
timestamp 1621523292
transform 1 0 57132 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1312_
timestamp 1621523292
transform 1 0 57500 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1621523292
transform -1 0 58880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_621
timestamp 1621523292
transform 1 0 58236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1101_
timestamp 1621523292
transform 1 0 2760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1214_
timestamp 1621523292
transform 1 0 1656 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1621523292
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1621523292
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1621523292
transform 1 0 2392 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_21
timestamp 1621523292
transform 1 0 3036 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_33
timestamp 1621523292
transform 1 0 4140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1621523292
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_45
timestamp 1621523292
transform 1 0 5244 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1621523292
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1621523292
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1621523292
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1621523292
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1621523292
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1621523292
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1621523292
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1621523292
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1621523292
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1621523292
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1621523292
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1621523292
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1621523292
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1621523292
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1621523292
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1621523292
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1621523292
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1621523292
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1621523292
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1621523292
transform 1 0 23276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1621523292
transform 1 0 24380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1621523292
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_277
timestamp 1621523292
transform 1 0 26588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1621523292
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_286
timestamp 1621523292
transform 1 0 27416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_298
timestamp 1621523292
transform 1 0 28520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_310
timestamp 1621523292
transform 1 0 29624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_322
timestamp 1621523292
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1621523292
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_334
timestamp 1621523292
transform 1 0 31832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1621523292
transform 1 0 32660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1621523292
transform 1 0 33764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1621523292
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1621523292
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1621523292
transform 1 0 37076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1621523292
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_400
timestamp 1621523292
transform 1 0 37904 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_412
timestamp 1621523292
transform 1 0 39008 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_424
timestamp 1621523292
transform 1 0 40112 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_436
timestamp 1621523292
transform 1 0 41216 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1621523292
transform 1 0 43056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_448
timestamp 1621523292
transform 1 0 42320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_457
timestamp 1621523292
transform 1 0 43148 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_469
timestamp 1621523292
transform 1 0 44252 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1164_
timestamp 1621523292
transform 1 0 47012 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1167_
timestamp 1621523292
transform 1 0 46368 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1621523292
transform 1 0 46828 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_481
timestamp 1621523292
transform 1 0 45356 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_489
timestamp 1621523292
transform 1 0 46092 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_495
timestamp 1621523292
transform 1 0 46644 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_502
timestamp 1621523292
transform 1 0 47288 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1621523292
transform 1 0 48760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1151_
timestamp 1621523292
transform 1 0 47656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1621523292
transform 1 0 48300 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_509
timestamp 1621523292
transform 1 0 47932 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_514
timestamp 1621523292
transform 1 0 48392 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_521
timestamp 1621523292
transform 1 0 49036 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 49404 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 50324 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_531
timestamp 1621523292
transform 1 0 49956 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_542
timestamp 1621523292
transform 1 0 50968 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0733_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51336 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0866_
timestamp 1621523292
transform 1 0 52348 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_551
timestamp 1621523292
transform 1 0 51796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_563
timestamp 1621523292
transform 1 0 52900 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0648_
timestamp 1621523292
transform 1 0 54004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1621523292
transform 1 0 54648 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1621523292
transform 1 0 53544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_569
timestamp 1621523292
transform 1 0 53452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_571
timestamp 1621523292
transform 1 0 53636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_578
timestamp 1621523292
transform 1 0 54280 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_585
timestamp 1621523292
transform 1 0 54924 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0919_
timestamp 1621523292
transform 1 0 55752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1274_
timestamp 1621523292
transform 1 0 56396 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_593
timestamp 1621523292
transform 1 0 55660 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_597
timestamp 1621523292
transform 1 0 56028 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_609
timestamp 1621523292
transform 1 0 57132 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1621523292
transform -1 0 58880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output208
timestamp 1621523292
transform 1 0 57868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1621523292
transform 1 0 58236 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1037_
timestamp 1621523292
transform 1 0 2484 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1621523292
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output317
timestamp 1621523292
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1621523292
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_11
timestamp 1621523292
transform 1 0 2116 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1621523292
transform 1 0 2760 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1038_
timestamp 1621523292
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1621523292
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_25
timestamp 1621523292
transform 1 0 3404 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1621523292
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1621523292
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1621523292
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1621523292
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1621523292
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1621523292
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1621523292
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1621523292
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1621523292
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1621523292
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1621523292
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1621523292
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1621523292
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1621523292
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1621523292
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1621523292
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1621523292
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1621523292
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1621523292
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_213
timestamp 1621523292
transform 1 0 20700 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_225
timestamp 1621523292
transform 1 0 21804 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1621523292
transform 1 0 22908 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1621523292
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_249
timestamp 1621523292
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1621523292
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_270
timestamp 1621523292
transform 1 0 25944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_282
timestamp 1621523292
transform 1 0 27048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_294
timestamp 1621523292
transform 1 0 28152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1621523292
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_306
timestamp 1621523292
transform 1 0 29256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1621523292
transform 1 0 30084 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_327
timestamp 1621523292
transform 1 0 31188 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_339
timestamp 1621523292
transform 1 0 32292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1621523292
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_351
timestamp 1621523292
transform 1 0 33396 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_363
timestamp 1621523292
transform 1 0 34500 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1621523292
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_384
timestamp 1621523292
transform 1 0 36432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_396
timestamp 1621523292
transform 1 0 37536 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_408
timestamp 1621523292
transform 1 0 38640 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1621523292
transform 1 0 40480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_420
timestamp 1621523292
transform 1 0 39744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_429
timestamp 1621523292
transform 1 0 40572 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_441
timestamp 1621523292
transform 1 0 41676 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_453
timestamp 1621523292
transform 1 0 42780 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_465
timestamp 1621523292
transform 1 0 43884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_477
timestamp 1621523292
transform 1 0 44988 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1168_
timestamp 1621523292
transform 1 0 46736 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1621523292
transform 1 0 45724 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_486
timestamp 1621523292
transform 1 0 45816 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_494
timestamp 1621523292
transform 1 0 46552 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_499
timestamp 1621523292
transform 1 0 47012 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0965_
timestamp 1621523292
transform 1 0 49312 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1050_
timestamp 1621523292
transform 1 0 48668 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1056_
timestamp 1621523292
transform 1 0 48024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1621523292
transform 1 0 47380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_506
timestamp 1621523292
transform 1 0 47656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_513
timestamp 1621523292
transform 1 0 48300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_520
timestamp 1621523292
transform 1 0 48944 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0655_
timestamp 1621523292
transform 1 0 49956 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1621523292
transform 1 0 50968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_527
timestamp 1621523292
transform 1 0 49588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_534
timestamp 1621523292
transform 1 0 50232 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_543
timestamp 1621523292
transform 1 0 51060 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1621523292
transform 1 0 51612 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_565
timestamp 1621523292
transform 1 0 53084 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1621523292
transform 1 0 55108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0726_
timestamp 1621523292
transform 1 0 53544 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0921_
timestamp 1621523292
transform 1 0 54464 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_569
timestamp 1621523292
transform 1 0 53452 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_573
timestamp 1621523292
transform 1 0 53820 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_579
timestamp 1621523292
transform 1 0 54372 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_583
timestamp 1621523292
transform 1 0 54740 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0917_
timestamp 1621523292
transform 1 0 56672 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1270_
timestamp 1621523292
transform 1 0 57316 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1621523292
transform 1 0 56212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_590
timestamp 1621523292
transform 1 0 55384 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_598
timestamp 1621523292
transform 1 0 56120 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_600
timestamp 1621523292
transform 1 0 56304 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_607
timestamp 1621523292
transform 1 0 56948 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1621523292
transform -1 0 58880 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_619
timestamp 1621523292
transform 1 0 58052 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1621523292
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output318
timestamp 1621523292
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output319
timestamp 1621523292
transform 1 0 2484 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1621523292
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1621523292
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1621523292
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_19
timestamp 1621523292
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_4  _1043_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3220 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _1102_
timestamp 1621523292
transform 1 0 4140 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_29
timestamp 1621523292
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_36
timestamp 1621523292
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1621523292
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1621523292
transform 1 0 5520 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1621523292
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1621523292
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1621523292
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1621523292
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1621523292
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1621523292
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1621523292
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1621523292
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1621523292
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1621523292
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1621523292
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1621523292
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1621523292
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1621523292
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1621523292
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1621523292
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1621523292
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1621523292
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1621523292
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_229
timestamp 1621523292
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_241
timestamp 1621523292
transform 1 0 23276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1621523292
transform 1 0 24380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1621523292
transform 1 0 25484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_277
timestamp 1621523292
transform 1 0 26588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1621523292
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1621523292
transform 1 0 27416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1621523292
transform 1 0 28520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1621523292
transform 1 0 29624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1621523292
transform 1 0 30728 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1621523292
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_334
timestamp 1621523292
transform 1 0 31832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_343
timestamp 1621523292
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1621523292
transform 1 0 33764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1621523292
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1621523292
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_391
timestamp 1621523292
transform 1 0 37076 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1621523292
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_400
timestamp 1621523292
transform 1 0 37904 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_412
timestamp 1621523292
transform 1 0 39008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_424
timestamp 1621523292
transform 1 0 40112 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_436
timestamp 1621523292
transform 1 0 41216 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1621523292
transform 1 0 43056 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_448
timestamp 1621523292
transform 1 0 42320 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_457
timestamp 1621523292
transform 1 0 43148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_469
timestamp 1621523292
transform 1 0 44252 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1621523292
transform 1 0 47012 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_481
timestamp 1621523292
transform 1 0 45356 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_493
timestamp 1621523292
transform 1 0 46460 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_502
timestamp 1621523292
transform 1 0 47288 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1621523292
transform 1 0 47656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1621523292
transform 1 0 48852 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1621523292
transform 1 0 48300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_509
timestamp 1621523292
transform 1 0 47932 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_514
timestamp 1621523292
transform 1 0 48392 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_518
timestamp 1621523292
transform 1 0 48760 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0654_
timestamp 1621523292
transform 1 0 50692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_535
timestamp 1621523292
transform 1 0 50324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_542
timestamp 1621523292
transform 1 0 50968 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1621523292
transform 1 0 51336 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0861_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1621523292
transform 1 0 51980 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_549
timestamp 1621523292
transform 1 0 51612 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_556
timestamp 1621523292
transform 1 0 52256 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_566
timestamp 1621523292
transform 1 0 53176 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1621523292
transform 1 0 54004 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1621523292
transform 1 0 53544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_571
timestamp 1621523292
transform 1 0 53636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1275_
timestamp 1621523292
transform 1 0 56396 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_591
timestamp 1621523292
transform 1 0 55476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_599
timestamp 1621523292
transform 1 0 56212 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_609
timestamp 1621523292
transform 1 0 57132 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1621523292
transform -1 0 58880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output247
timestamp 1621523292
transform 1 0 57868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_621
timestamp 1621523292
transform 1 0 58236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1036_
timestamp 1621523292
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1215_
timestamp 1621523292
transform 1 0 1656 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1621523292
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1621523292
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1621523292
transform 1 0 2392 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1621523292
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1621523292
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1621523292
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1621523292
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1621523292
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1621523292
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1621523292
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1621523292
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1621523292
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1621523292
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1621523292
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1621523292
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1621523292
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1621523292
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1621523292
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1621523292
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1621523292
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1621523292
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1621523292
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1621523292
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1621523292
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1621523292
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_225
timestamp 1621523292
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_237
timestamp 1621523292
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1621523292
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_249
timestamp 1621523292
transform 1 0 24012 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1621523292
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1621523292
transform 1 0 25944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1621523292
transform 1 0 27048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1621523292
transform 1 0 28152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1621523292
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_306
timestamp 1621523292
transform 1 0 29256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_315
timestamp 1621523292
transform 1 0 30084 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_327
timestamp 1621523292
transform 1 0 31188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_339
timestamp 1621523292
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1621523292
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1621523292
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1621523292
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1621523292
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1621523292
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_396
timestamp 1621523292
transform 1 0 37536 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_408
timestamp 1621523292
transform 1 0 38640 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1621523292
transform 1 0 40480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_420
timestamp 1621523292
transform 1 0 39744 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_429
timestamp 1621523292
transform 1 0 40572 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_441
timestamp 1621523292
transform 1 0 41676 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_453
timestamp 1621523292
transform 1 0 42780 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_465
timestamp 1621523292
transform 1 0 43884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1621523292
transform 1 0 44988 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1621523292
transform 1 0 45724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_486
timestamp 1621523292
transform 1 0 45816 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_498
timestamp 1621523292
transform 1 0 46920 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0964_
timestamp 1621523292
transform 1 0 49312 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1055_
timestamp 1621523292
transform 1 0 48668 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1621523292
transform 1 0 48024 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_513
timestamp 1621523292
transform 1 0 48300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_520
timestamp 1621523292
transform 1 0 48944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0872_
timestamp 1621523292
transform 1 0 49956 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1621523292
transform 1 0 50968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_527
timestamp 1621523292
transform 1 0 49588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_538
timestamp 1621523292
transform 1 0 50600 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_543
timestamp 1621523292
transform 1 0 51060 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0646_
timestamp 1621523292
transform 1 0 51428 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1621523292
transform 1 0 52256 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0860_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52900 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_12_551
timestamp 1621523292
transform 1 0 51796 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_555
timestamp 1621523292
transform 1 0 52164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_559
timestamp 1621523292
transform 1 0 52532 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0647_
timestamp 1621523292
transform 1 0 53728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0719_
timestamp 1621523292
transform 1 0 54464 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_568
timestamp 1621523292
transform 1 0 53360 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_575
timestamp 1621523292
transform 1 0 54004 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_579
timestamp 1621523292
transform 1 0 54372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_587
timestamp 1621523292
transform 1 0 55108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0645_
timestamp 1621523292
transform 1 0 55476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0916_
timestamp 1621523292
transform 1 0 56856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1621523292
transform 1 0 56212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_594
timestamp 1621523292
transform 1 0 55752 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_598
timestamp 1621523292
transform 1 0 56120 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_600
timestamp 1621523292
transform 1 0 56304 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_609
timestamp 1621523292
transform 1 0 57132 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1313_
timestamp 1621523292
transform 1 0 57500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1621523292
transform -1 0 58880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1621523292
transform 1 0 58236 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1621523292
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1621523292
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output289
timestamp 1621523292
transform 1 0 1748 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1621523292
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1621523292
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1216_
timestamp 1621523292
transform 1 0 1748 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1621523292
transform 1 0 2116 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1621523292
transform 1 0 2484 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1034_
timestamp 1621523292
transform 1 0 2484 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_18
timestamp 1621523292
transform 1 0 2760 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1621523292
transform 1 0 2852 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1103_
timestamp 1621523292
transform 1 0 3496 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1104_
timestamp 1621523292
transform 1 0 3128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1621523292
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_22
timestamp 1621523292
transform 1 0 3128 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_29
timestamp 1621523292
transform 1 0 3772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1621523292
transform 1 0 4876 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_25
timestamp 1621523292
transform 1 0 3404 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1621523292
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1621523292
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1621523292
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_53
timestamp 1621523292
transform 1 0 5980 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1621523292
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1621523292
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1621523292
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1621523292
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1621523292
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1621523292
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1621523292
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1621523292
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1621523292
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1621523292
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1621523292
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1621523292
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1621523292
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1621523292
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1621523292
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1621523292
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1621523292
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1621523292
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1621523292
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1621523292
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1621523292
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1621523292
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1621523292
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1621523292
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1621523292
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1621523292
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1621523292
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1621523292
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1621523292
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1621523292
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1621523292
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1621523292
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1621523292
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1621523292
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1621523292
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1621523292
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1621523292
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1621523292
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1621523292
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1621523292
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1621523292
transform 1 0 23276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1621523292
transform 1 0 24380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_249
timestamp 1621523292
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1621523292
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1621523292
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1621523292
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_270
timestamp 1621523292
transform 1 0 25944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_282
timestamp 1621523292
transform 1 0 27048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1621523292
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1621523292
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_298
timestamp 1621523292
transform 1 0 28520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_294
timestamp 1621523292
transform 1 0 28152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1621523292
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_310
timestamp 1621523292
transform 1 0 29624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_322
timestamp 1621523292
transform 1 0 30728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_306
timestamp 1621523292
transform 1 0 29256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_315
timestamp 1621523292
transform 1 0 30084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_327
timestamp 1621523292
transform 1 0 31188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1621523292
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_334
timestamp 1621523292
transform 1 0 31832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1621523292
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_339
timestamp 1621523292
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1621523292
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_355
timestamp 1621523292
transform 1 0 33764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1621523292
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1621523292
transform 1 0 33396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_363
timestamp 1621523292
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1621523292
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_391
timestamp 1621523292
transform 1 0 37076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1621523292
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1621523292
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1621523292
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_400
timestamp 1621523292
transform 1 0 37904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_412
timestamp 1621523292
transform 1 0 39008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_396
timestamp 1621523292
transform 1 0 37536 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_408
timestamp 1621523292
transform 1 0 38640 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1621523292
transform 1 0 40480 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_424
timestamp 1621523292
transform 1 0 40112 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_436
timestamp 1621523292
transform 1 0 41216 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_420
timestamp 1621523292
transform 1 0 39744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_429
timestamp 1621523292
transform 1 0 40572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1621523292
transform 1 0 43056 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_448
timestamp 1621523292
transform 1 0 42320 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_457
timestamp 1621523292
transform 1 0 43148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_441
timestamp 1621523292
transform 1 0 41676 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_453
timestamp 1621523292
transform 1 0 42780 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_469
timestamp 1621523292
transform 1 0 44252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_465
timestamp 1621523292
transform 1 0 43884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1621523292
transform 1 0 44988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1621523292
transform 1 0 45724 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_481
timestamp 1621523292
transform 1 0 45356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_493
timestamp 1621523292
transform 1 0 46460 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_486
timestamp 1621523292
transform 1 0 45816 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_498
timestamp 1621523292
transform 1 0 46920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1621523292
transform 1 0 49036 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1621523292
transform 1 0 48300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1621523292
transform 1 0 49312 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1621523292
transform 1 0 47564 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_514
timestamp 1621523292
transform 1 0 48392 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_520
timestamp 1621523292
transform 1 0 48944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1621523292
transform 1 0 48024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_522
timestamp 1621523292
transform 1 0 49128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _0863_
timestamp 1621523292
transform 1 0 51152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1621523292
transform 1 0 49956 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1621523292
transform 1 0 50968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_537
timestamp 1621523292
transform 1 0 50508 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_543
timestamp 1621523292
transform 1 0 51060 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_527
timestamp 1621523292
transform 1 0 49588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_536
timestamp 1621523292
transform 1 0 50416 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_543
timestamp 1621523292
transform 1 0 51060 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51888 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0864_
timestamp 1621523292
transform 1 0 53268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1621523292
transform 1 0 51428 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_547
timestamp 1621523292
transform 1 0 51428 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_551
timestamp 1621523292
transform 1 0 51796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_560
timestamp 1621523292
transform 1 0 52624 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_563
timestamp 1621523292
transform 1 0 52900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0643_
timestamp 1621523292
transform 1 0 54556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0717_
timestamp 1621523292
transform 1 0 55200 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1621523292
transform 1 0 54004 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1621523292
transform 1 0 53544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_568
timestamp 1621523292
transform 1 0 53360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_571
timestamp 1621523292
transform 1 0 53636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_575
timestamp 1621523292
transform 1 0 54004 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_584
timestamp 1621523292
transform 1 0 54832 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_595
timestamp 1621523292
transform 1 0 55844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_598
timestamp 1621523292
transform 1 0 56120 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_591
timestamp 1621523292
transform 1 0 55476 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1621523292
transform 1 0 55844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_604
timestamp 1621523292
transform 1 0 56672 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_600
timestamp 1621523292
transform 1 0 56304 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_604
timestamp 1621523292
transform 1 0 56672 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output248
timestamp 1621523292
transform 1 0 56764 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1621523292
transform 1 0 56212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1276_
timestamp 1621523292
transform 1 0 56764 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_609
timestamp 1621523292
transform 1 0 57132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1314_
timestamp 1621523292
transform 1 0 57500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1621523292
transform -1 0 58880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1621523292
transform -1 0 58880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output209
timestamp 1621523292
transform 1 0 57868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_613
timestamp 1621523292
transform 1 0 57500 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1621523292
transform 1 0 58236 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1621523292
transform 1 0 58236 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1217_
timestamp 1621523292
transform 1 0 1656 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1621523292
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1621523292
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_14
timestamp 1621523292
transform 1 0 2392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1621523292
transform 1 0 3496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1621523292
transform 1 0 4600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1621523292
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1621523292
transform 1 0 5704 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_56
timestamp 1621523292
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1621523292
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1621523292
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1621523292
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1621523292
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1621523292
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1621523292
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1621523292
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1621523292
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1621523292
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1621523292
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1621523292
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1621523292
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1621523292
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1621523292
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1621523292
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1621523292
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1621523292
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1621523292
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1621523292
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1621523292
transform 1 0 23276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1621523292
transform 1 0 24380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1621523292
transform 1 0 25484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_277
timestamp 1621523292
transform 1 0 26588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1621523292
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1621523292
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_298
timestamp 1621523292
transform 1 0 28520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_310
timestamp 1621523292
transform 1 0 29624 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_322
timestamp 1621523292
transform 1 0 30728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1621523292
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_334
timestamp 1621523292
transform 1 0 31832 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1621523292
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1621523292
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1621523292
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1621523292
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1621523292
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1621523292
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_400
timestamp 1621523292
transform 1 0 37904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_412
timestamp 1621523292
transform 1 0 39008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_424
timestamp 1621523292
transform 1 0 40112 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_436
timestamp 1621523292
transform 1 0 41216 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1621523292
transform 1 0 43056 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_448
timestamp 1621523292
transform 1 0 42320 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_457
timestamp 1621523292
transform 1 0 43148 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_469
timestamp 1621523292
transform 1 0 44252 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_481
timestamp 1621523292
transform 1 0 45356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_493
timestamp 1621523292
transform 1 0 46460 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1621523292
transform 1 0 48300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1621523292
transform 1 0 47564 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_514
timestamp 1621523292
transform 1 0 48392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1621523292
transform 1 0 51244 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1169_
timestamp 1621523292
transform 1 0 50600 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1170_
timestamp 1621523292
transform 1 0 49956 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_526
timestamp 1621523292
transform 1 0 49496 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_530
timestamp 1621523292
transform 1 0 49864 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_534
timestamp 1621523292
transform 1 0 50232 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_541
timestamp 1621523292
transform 1 0 50876 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1621523292
transform 1 0 52900 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0838_
timestamp 1621523292
transform 1 0 51888 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_548
timestamp 1621523292
transform 1 0 51520 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_556
timestamp 1621523292
transform 1 0 52256 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_562
timestamp 1621523292
transform 1 0 52808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_566
timestamp 1621523292
transform 1 0 53176 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0740_
timestamp 1621523292
transform 1 0 54464 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1621523292
transform 1 0 53544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_571
timestamp 1621523292
transform 1 0 53636 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_579
timestamp 1621523292
transform 1 0 54372 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_587
timestamp 1621523292
transform 1 0 55108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1621523292
transform 1 0 55476 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_607
timestamp 1621523292
transform 1 0 56948 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1621523292
transform -1 0 58880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output210
timestamp 1621523292
transform 1 0 57868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_615
timestamp 1621523292
transform 1 0 57684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1621523292
transform 1 0 58236 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1621523292
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1218_
timestamp 1621523292
transform 1 0 1840 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1621523292
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1621523292
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1621523292
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_16
timestamp 1621523292
transform 1 0 2576 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1621523292
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_23
timestamp 1621523292
transform 1 0 3220 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1621523292
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1621523292
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1621523292
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1621523292
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1621523292
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1621523292
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1621523292
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1621523292
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1621523292
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1621523292
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1621523292
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1621523292
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1621523292
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1621523292
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1621523292
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1621523292
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1621523292
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1621523292
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1621523292
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1621523292
transform 1 0 20700 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1621523292
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1621523292
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1621523292
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1621523292
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1621523292
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_270
timestamp 1621523292
transform 1 0 25944 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_282
timestamp 1621523292
transform 1 0 27048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_294
timestamp 1621523292
transform 1 0 28152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1621523292
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_306
timestamp 1621523292
transform 1 0 29256 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1621523292
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1621523292
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1621523292
transform 1 0 32292 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1621523292
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1621523292
transform 1 0 33396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_363
timestamp 1621523292
transform 1 0 34500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1621523292
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1621523292
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_396
timestamp 1621523292
transform 1 0 37536 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_408
timestamp 1621523292
transform 1 0 38640 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1621523292
transform 1 0 40480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_420
timestamp 1621523292
transform 1 0 39744 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_429
timestamp 1621523292
transform 1 0 40572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_441
timestamp 1621523292
transform 1 0 41676 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_453
timestamp 1621523292
transform 1 0 42780 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_465
timestamp 1621523292
transform 1 0 43884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_477
timestamp 1621523292
transform 1 0 44988 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1621523292
transform 1 0 45724 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_486
timestamp 1621523292
transform 1 0 45816 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_498
timestamp 1621523292
transform 1 0 46920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1621523292
transform 1 0 49036 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_510
timestamp 1621523292
transform 1 0 48024 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_518
timestamp 1621523292
transform 1 0 48760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_524
timestamp 1621523292
transform 1 0 49312 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1621523292
transform 1 0 50324 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1171_
timestamp 1621523292
transform 1 0 49680 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1621523292
transform 1 0 50968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_531
timestamp 1621523292
transform 1 0 49956 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_538
timestamp 1621523292
transform 1 0 50600 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_543
timestamp 1621523292
transform 1 0 51060 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1621523292
transform 1 0 51428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _0744_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52532 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_16_550
timestamp 1621523292
transform 1 0 51704 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_558
timestamp 1621523292
transform 1 0 52440 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _0741_
timestamp 1621523292
transform 1 0 55108 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 53820 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_569
timestamp 1621523292
transform 1 0 53452 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_583
timestamp 1621523292
transform 1 0 54740 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0644_
timestamp 1621523292
transform 1 0 56672 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1621523292
transform 1 0 56212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_594
timestamp 1621523292
transform 1 0 55752 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_598
timestamp 1621523292
transform 1 0 56120 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_600
timestamp 1621523292
transform 1 0 56304 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_607
timestamp 1621523292
transform 1 0 56948 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1621523292
transform -1 0 58880 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output249
timestamp 1621523292
transform 1 0 57868 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_615
timestamp 1621523292
transform 1 0 57684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1621523292
transform 1 0 58236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1621523292
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output290
timestamp 1621523292
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output291
timestamp 1621523292
transform 1 0 2484 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1621523292
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_11
timestamp 1621523292
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_19
timestamp 1621523292
transform 1 0 2852 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1032_
timestamp 1621523292
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1105_
timestamp 1621523292
transform 1 0 3864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1621523292
transform 1 0 3496 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_33
timestamp 1621523292
transform 1 0 4140 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1621523292
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_45
timestamp 1621523292
transform 1 0 5244 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1621523292
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1621523292
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1621523292
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1621523292
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1621523292
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1621523292
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1621523292
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1621523292
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1621523292
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1621523292
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1621523292
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1621523292
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1621523292
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1621523292
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1621523292
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1621523292
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1621523292
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1621523292
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1621523292
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1621523292
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1621523292
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1621523292
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1621523292
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1621523292
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1621523292
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_298
timestamp 1621523292
transform 1 0 28520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_310
timestamp 1621523292
transform 1 0 29624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1621523292
transform 1 0 30728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1621523292
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1621523292
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1621523292
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1621523292
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1621523292
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1621523292
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_391
timestamp 1621523292
transform 1 0 37076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1621523292
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_400
timestamp 1621523292
transform 1 0 37904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_412
timestamp 1621523292
transform 1 0 39008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_424
timestamp 1621523292
transform 1 0 40112 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_436
timestamp 1621523292
transform 1 0 41216 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1621523292
transform 1 0 43056 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_448
timestamp 1621523292
transform 1 0 42320 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_457
timestamp 1621523292
transform 1 0 43148 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_469
timestamp 1621523292
transform 1 0 44252 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_481
timestamp 1621523292
transform 1 0 45356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_493
timestamp 1621523292
transform 1 0 46460 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1064_
timestamp 1621523292
transform 1 0 49220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1621523292
transform 1 0 48300 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1621523292
transform 1 0 47564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_514
timestamp 1621523292
transform 1 0 48392 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_522
timestamp 1621523292
transform 1 0 49128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1621523292
transform 1 0 49864 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_526
timestamp 1621523292
transform 1 0 49496 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0639_
timestamp 1621523292
transform 1 0 51704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0743_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52348 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_546
timestamp 1621523292
transform 1 0 51336 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_553
timestamp 1621523292
transform 1 0 51980 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_566
timestamp 1621523292
transform 1 0 53176 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0724_
timestamp 1621523292
transform 1 0 54556 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1621523292
transform 1 0 53544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_571
timestamp 1621523292
transform 1 0 53636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_579
timestamp 1621523292
transform 1 0 54372 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_588
timestamp 1621523292
transform 1 0 55200 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0642_
timestamp 1621523292
transform 1 0 55568 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0914_
timestamp 1621523292
transform 1 0 56488 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1277_
timestamp 1621523292
transform 1 0 57132 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_595
timestamp 1621523292
transform 1 0 55844 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_601
timestamp 1621523292
transform 1 0 56396 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_605
timestamp 1621523292
transform 1 0 56764 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1621523292
transform -1 0 58880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_617
timestamp 1621523292
transform 1 0 57868 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1031_
timestamp 1621523292
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1219_
timestamp 1621523292
transform 1 0 1564 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1621523292
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1621523292
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1621523292
transform 1 0 2300 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1621523292
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1106_
timestamp 1621523292
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1621523292
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1621523292
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_30
timestamp 1621523292
transform 1 0 3864 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_37
timestamp 1621523292
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_49
timestamp 1621523292
transform 1 0 5612 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_61
timestamp 1621523292
transform 1 0 6716 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1621523292
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_73
timestamp 1621523292
transform 1 0 7820 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1621523292
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1621523292
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1621523292
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1621523292
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1621523292
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1621523292
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1621523292
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1621523292
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1621523292
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1621523292
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1621523292
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1621523292
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1621523292
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1621523292
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1621523292
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1621523292
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1621523292
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1621523292
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1621523292
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1621523292
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1621523292
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1621523292
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_294
timestamp 1621523292
transform 1 0 28152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1621523292
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_306
timestamp 1621523292
transform 1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1621523292
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_327
timestamp 1621523292
transform 1 0 31188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_339
timestamp 1621523292
transform 1 0 32292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1621523292
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1621523292
transform 1 0 33396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_363
timestamp 1621523292
transform 1 0 34500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1621523292
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1621523292
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_396
timestamp 1621523292
transform 1 0 37536 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_408
timestamp 1621523292
transform 1 0 38640 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1621523292
transform 1 0 40480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_420
timestamp 1621523292
transform 1 0 39744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_429
timestamp 1621523292
transform 1 0 40572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_441
timestamp 1621523292
transform 1 0 41676 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_453
timestamp 1621523292
transform 1 0 42780 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_465
timestamp 1621523292
transform 1 0 43884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1621523292
transform 1 0 44988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1621523292
transform 1 0 45724 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_486
timestamp 1621523292
transform 1 0 45816 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_498
timestamp 1621523292
transform 1 0 46920 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_510
timestamp 1621523292
transform 1 0 48024 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_522
timestamp 1621523292
transform 1 0 49128 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1621523292
transform 1 0 50324 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0962_
timestamp 1621523292
transform 1 0 49680 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1621523292
transform 1 0 50968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_531
timestamp 1621523292
transform 1 0 49956 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_538
timestamp 1621523292
transform 1 0 50600 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_543
timestamp 1621523292
transform 1 0 51060 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0722_
timestamp 1621523292
transform 1 0 51428 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0859_
timestamp 1621523292
transform 1 0 52532 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_554
timestamp 1621523292
transform 1 0 52072 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_558
timestamp 1621523292
transform 1 0 52440 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_567
timestamp 1621523292
transform 1 0 53268 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1621523292
transform 1 0 53636 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_587
timestamp 1621523292
transform 1 0 55108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0641_
timestamp 1621523292
transform 1 0 55476 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1621523292
transform 1 0 56672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1621523292
transform 1 0 56212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_594
timestamp 1621523292
transform 1 0 55752 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_598
timestamp 1621523292
transform 1 0 56120 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_600
timestamp 1621523292
transform 1 0 56304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_607
timestamp 1621523292
transform 1 0 56948 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _1315_
timestamp 1621523292
transform 1 0 57500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1621523292
transform -1 0 58880 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1621523292
transform 1 0 58236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1621523292
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1621523292
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output292
timestamp 1621523292
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1621523292
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1621523292
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1220_
timestamp 1621523292
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_14
timestamp 1621523292
transform 1 0 2392 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_17
timestamp 1621523292
transform 1 0 2668 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_11
timestamp 1621523292
transform 1 0 2116 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_21
timestamp 1621523292
transform 1 0 3036 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1107_
timestamp 1621523292
transform 1 0 2760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1006_
timestamp 1621523292
transform 1 0 2760 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _0874_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4968 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1621523292
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_22
timestamp 1621523292
transform 1 0 3128 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_34
timestamp 1621523292
transform 1 0 4232 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1621523292
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1621523292
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1621523292
transform 1 0 5336 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_54
timestamp 1621523292
transform 1 0 6072 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1621523292
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_49
timestamp 1621523292
transform 1 0 5612 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_61
timestamp 1621523292
transform 1 0 6716 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1621523292
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1621523292
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1621523292
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_73
timestamp 1621523292
transform 1 0 7820 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1621523292
transform 1 0 8924 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1621523292
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1621523292
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1621523292
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1621523292
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1621523292
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1621523292
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1621523292
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1621523292
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1621523292
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1621523292
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1621523292
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1621523292
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1621523292
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1621523292
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1621523292
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1621523292
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1621523292
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1621523292
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1621523292
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1621523292
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1621523292
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1621523292
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1621523292
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1621523292
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1621523292
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1621523292
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1621523292
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1621523292
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1621523292
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1621523292
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1621523292
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1621523292
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1621523292
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1621523292
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1621523292
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1621523292
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1621523292
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1621523292
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1621523292
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1621523292
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1621523292
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1621523292
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1621523292
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1621523292
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1621523292
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1621523292
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_310
timestamp 1621523292
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1621523292
transform 1 0 30728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_306
timestamp 1621523292
transform 1 0 29256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1621523292
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_327
timestamp 1621523292
transform 1 0 31188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1621523292
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_334
timestamp 1621523292
transform 1 0 31832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_343
timestamp 1621523292
transform 1 0 32660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1621523292
transform 1 0 32292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1621523292
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_355
timestamp 1621523292
transform 1 0 33764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1621523292
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1621523292
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1621523292
transform 1 0 34500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1621523292
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_391
timestamp 1621523292
transform 1 0 37076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1621523292
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1621523292
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1621523292
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_400
timestamp 1621523292
transform 1 0 37904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1621523292
transform 1 0 39008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_396
timestamp 1621523292
transform 1 0 37536 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1621523292
transform 1 0 38640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1621523292
transform 1 0 40480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_424
timestamp 1621523292
transform 1 0 40112 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_436
timestamp 1621523292
transform 1 0 41216 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_420
timestamp 1621523292
transform 1 0 39744 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_429
timestamp 1621523292
transform 1 0 40572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1621523292
transform 1 0 43056 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_448
timestamp 1621523292
transform 1 0 42320 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_457
timestamp 1621523292
transform 1 0 43148 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_441
timestamp 1621523292
transform 1 0 41676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_453
timestamp 1621523292
transform 1 0 42780 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_469
timestamp 1621523292
transform 1 0 44252 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_465
timestamp 1621523292
transform 1 0 43884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1621523292
transform 1 0 44988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1621523292
transform 1 0 45724 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_481
timestamp 1621523292
transform 1 0 45356 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_493
timestamp 1621523292
transform 1 0 46460 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_486
timestamp 1621523292
transform 1 0 45816 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_498
timestamp 1621523292
transform 1 0 46920 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0875_
timestamp 1621523292
transform 1 0 47748 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _1172_
timestamp 1621523292
transform 1 0 49128 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1621523292
transform 1 0 48300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1621523292
transform 1 0 47564 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_514
timestamp 1621523292
transform 1 0 48392 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_506
timestamp 1621523292
transform 1 0 47656 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_513
timestamp 1621523292
transform 1 0 48300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_531
timestamp 1621523292
transform 1 0 49956 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_525
timestamp 1621523292
transform 1 0 49404 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_525
timestamp 1621523292
transform 1 0 49404 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0961_
timestamp 1621523292
transform 1 0 49680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0858_
timestamp 1621523292
transform 1 0 50324 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_543
timestamp 1621523292
transform 1 0 51060 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_538
timestamp 1621523292
transform 1 0 50600 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_545
timestamp 1621523292
transform 1 0 51244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1621523292
transform 1 0 50968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1621523292
transform 1 0 49772 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1621523292
transform 1 0 51612 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0742_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52532 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0856_
timestamp 1621523292
transform 1 0 52624 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_1  _0857_
timestamp 1621523292
transform 1 0 51428 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_19_552
timestamp 1621523292
transform 1 0 51888 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_558
timestamp 1621523292
transform 1 0 52440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_566
timestamp 1621523292
transform 1 0 53176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_554
timestamp 1621523292
transform 1 0 52072 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_566
timestamp 1621523292
transform 1 0 53176 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_576
timestamp 1621523292
transform 1 0 54096 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_572
timestamp 1621523292
transform 1 0 53728 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_578
timestamp 1621523292
transform 1 0 54280 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_571
timestamp 1621523292
transform 1 0 53636 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1621523292
transform 1 0 53544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _0725_
timestamp 1621523292
transform 1 0 54004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1621523292
transform 1 0 53820 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_584
timestamp 1621523292
transform 1 0 54832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_580
timestamp 1621523292
transform 1 0 54464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1621523292
transform 1 0 54556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0636_
timestamp 1621523292
transform 1 0 55200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1621523292
transform 1 0 55016 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__ebufn_1  _1278_
timestamp 1621523292
transform 1 0 57040 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1621523292
transform 1 0 56212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output250
timestamp 1621523292
transform 1 0 57132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_602
timestamp 1621523292
transform 1 0 56488 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_608
timestamp 1621523292
transform 1 0 57040 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_591
timestamp 1621523292
transform 1 0 55476 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_600
timestamp 1621523292
transform 1 0 56304 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1621523292
transform -1 0 58880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1621523292
transform -1 0 58880 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output211
timestamp 1621523292
transform 1 0 57868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_613
timestamp 1621523292
transform 1 0 57500 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1621523292
transform 1 0 58236 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_616
timestamp 1621523292
transform 1 0 57776 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1621523292
transform 1 0 58512 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1621523292
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1621523292
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output293
timestamp 1621523292
transform 1 0 1748 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1621523292
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1621523292
transform 1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1621523292
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1030_
timestamp 1621523292
transform 1 0 3128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1108_
timestamp 1621523292
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1621523292
transform 1 0 3404 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1621523292
transform 1 0 4048 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1621523292
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1621523292
transform 1 0 5152 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1621523292
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1621523292
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1621523292
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1621523292
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1621523292
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1621523292
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1621523292
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1621523292
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1621523292
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1621523292
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1621523292
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1621523292
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1621523292
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1621523292
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1621523292
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1621523292
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1621523292
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1621523292
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1621523292
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1621523292
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1621523292
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1621523292
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1621523292
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1621523292
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1621523292
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1621523292
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1621523292
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1621523292
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1621523292
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1621523292
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1621523292
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1621523292
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_355
timestamp 1621523292
transform 1 0 33764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1621523292
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1621523292
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1621523292
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1621523292
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_400
timestamp 1621523292
transform 1 0 37904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1621523292
transform 1 0 39008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_424
timestamp 1621523292
transform 1 0 40112 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_436
timestamp 1621523292
transform 1 0 41216 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1621523292
transform 1 0 43056 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_448
timestamp 1621523292
transform 1 0 42320 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_457
timestamp 1621523292
transform 1 0 43148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_469
timestamp 1621523292
transform 1 0 44252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1621523292
transform 1 0 45356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_493
timestamp 1621523292
transform 1 0 46460 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1621523292
transform 1 0 48300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1621523292
transform 1 0 49128 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1621523292
transform 1 0 47564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_514
timestamp 1621523292
transform 1 0 48392 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0635_
timestamp 1621523292
transform 1 0 51060 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1065_
timestamp 1621523292
transform 1 0 50416 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1621523292
transform 1 0 49772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_525
timestamp 1621523292
transform 1 0 49404 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_532
timestamp 1621523292
transform 1 0 50048 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_539
timestamp 1621523292
transform 1 0 50692 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0638_
timestamp 1621523292
transform 1 0 52532 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0915_
timestamp 1621523292
transform 1 0 51888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_547
timestamp 1621523292
transform 1 0 51428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_551
timestamp 1621523292
transform 1 0 51796 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_555
timestamp 1621523292
transform 1 0 52164 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_562
timestamp 1621523292
transform 1 0 52808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0747_
timestamp 1621523292
transform 1 0 54188 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1621523292
transform 1 0 53544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output251
timestamp 1621523292
transform 1 0 55200 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_571
timestamp 1621523292
transform 1 0 53636 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_584
timestamp 1621523292
transform 1 0 54832 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1621523292
transform 1 0 55936 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output212
timestamp 1621523292
transform 1 0 56764 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_592
timestamp 1621523292
transform 1 0 55568 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_600
timestamp 1621523292
transform 1 0 56304 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_604
timestamp 1621523292
transform 1 0 56672 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_609
timestamp 1621523292
transform 1 0 57132 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1316_
timestamp 1621523292
transform 1 0 57500 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1621523292
transform -1 0 58880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_621
timestamp 1621523292
transform 1 0 58236 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1221_
timestamp 1621523292
transform 1 0 1840 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1621523292
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1621523292
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1621523292
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_16
timestamp 1621523292
transform 1 0 2576 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1621523292
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_28
timestamp 1621523292
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1621523292
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1621523292
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1621523292
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1621523292
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1621523292
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1621523292
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1621523292
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1621523292
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1621523292
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1621523292
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1621523292
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1621523292
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1621523292
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1621523292
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1621523292
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1621523292
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1621523292
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1621523292
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1621523292
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1621523292
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1621523292
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1621523292
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1621523292
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1621523292
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1621523292
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1621523292
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1621523292
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1621523292
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1621523292
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1621523292
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_315
timestamp 1621523292
transform 1 0 30084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_327
timestamp 1621523292
transform 1 0 31188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1621523292
transform 1 0 32292 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1621523292
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1621523292
transform 1 0 33396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1621523292
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1621523292
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_384
timestamp 1621523292
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_396
timestamp 1621523292
transform 1 0 37536 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_408
timestamp 1621523292
transform 1 0 38640 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1621523292
transform 1 0 40480 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_420
timestamp 1621523292
transform 1 0 39744 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_429
timestamp 1621523292
transform 1 0 40572 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_441
timestamp 1621523292
transform 1 0 41676 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_453
timestamp 1621523292
transform 1 0 42780 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_465
timestamp 1621523292
transform 1 0 43884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_477
timestamp 1621523292
transform 1 0 44988 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1621523292
transform 1 0 45724 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_486
timestamp 1621523292
transform 1 0 45816 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1621523292
transform 1 0 46920 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_510
timestamp 1621523292
transform 1 0 48024 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_522
timestamp 1621523292
transform 1 0 49128 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0960_
timestamp 1621523292
transform 1 0 50324 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1066_
timestamp 1621523292
transform 1 0 49680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1621523292
transform 1 0 50968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_531
timestamp 1621523292
transform 1 0 49956 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_538
timestamp 1621523292
transform 1 0 50600 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_543
timestamp 1621523292
transform 1 0 51060 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0852_
timestamp 1621523292
transform 1 0 51428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1621523292
transform 1 0 52348 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_550
timestamp 1621523292
transform 1 0 51704 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_556
timestamp 1621523292
transform 1 0 52256 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0711_
timestamp 1621523292
transform 1 0 54188 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0714_
timestamp 1621523292
transform 1 0 55200 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_573
timestamp 1621523292
transform 1 0 53820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_584
timestamp 1621523292
transform 1 0 54832 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1279_
timestamp 1621523292
transform 1 0 57224 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1621523292
transform 1 0 56212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_595
timestamp 1621523292
transform 1 0 55844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_600
timestamp 1621523292
transform 1 0 56304 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_608
timestamp 1621523292
transform 1 0 57040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1621523292
transform -1 0 58880 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_618
timestamp 1621523292
transform 1 0 57960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_624
timestamp 1621523292
transform 1 0 58512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1621523292
transform 1 0 2852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1222_
timestamp 1621523292
transform 1 0 1748 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1621523292
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1621523292
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_15
timestamp 1621523292
transform 1 0 2484 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_22
timestamp 1621523292
transform 1 0 3128 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_34
timestamp 1621523292
transform 1 0 4232 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1621523292
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1621523292
transform 1 0 5336 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_54
timestamp 1621523292
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1621523292
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1621523292
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1621523292
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1621523292
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1621523292
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1621523292
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1621523292
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1621523292
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1621523292
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1621523292
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1621523292
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1621523292
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1621523292
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1621523292
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1621523292
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1621523292
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1621523292
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_220
timestamp 1621523292
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1621523292
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1621523292
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1621523292
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1621523292
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1621523292
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1621523292
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1621523292
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1621523292
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1621523292
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1621523292
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1621523292
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1621523292
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1621523292
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1621523292
transform 1 0 33764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1621523292
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1621523292
transform 1 0 35972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_391
timestamp 1621523292
transform 1 0 37076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1621523292
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1621523292
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1621523292
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_424
timestamp 1621523292
transform 1 0 40112 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_436
timestamp 1621523292
transform 1 0 41216 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1621523292
transform 1 0 43056 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_448
timestamp 1621523292
transform 1 0 42320 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_457
timestamp 1621523292
transform 1 0 43148 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_469
timestamp 1621523292
transform 1 0 44252 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_481
timestamp 1621523292
transform 1 0 45356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_493
timestamp 1621523292
transform 1 0 46460 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1621523292
transform 1 0 48300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1621523292
transform 1 0 47564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_514
timestamp 1621523292
transform 1 0 48392 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1173_
timestamp 1621523292
transform 1 0 49772 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1621523292
transform 1 0 50416 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_23_526
timestamp 1621523292
transform 1 0 49496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_532
timestamp 1621523292
transform 1 0 50048 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0850_
timestamp 1621523292
transform 1 0 52256 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_552
timestamp 1621523292
transform 1 0 51888 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_562
timestamp 1621523292
transform 1 0 52808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _0748_
timestamp 1621523292
transform 1 0 54096 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1621523292
transform 1 0 55108 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1621523292
transform 1 0 53544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_571
timestamp 1621523292
transform 1 0 53636 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_575
timestamp 1621523292
transform 1 0 54004 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_583
timestamp 1621523292
transform 1 0 54740 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_603
timestamp 1621523292
transform 1 0 56580 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_611
timestamp 1621523292
transform 1 0 57316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1317_
timestamp 1621523292
transform 1 0 57500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1621523292
transform -1 0 58880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1621523292
transform 1 0 58236 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1621523292
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output294
timestamp 1621523292
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output295
timestamp 1621523292
transform 1 0 2484 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1621523292
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1621523292
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1621523292
transform 1 0 2852 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1621523292
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1621523292
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1621523292
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1621523292
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1621523292
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1621523292
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1621523292
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1621523292
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1621523292
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1621523292
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1621523292
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1621523292
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1621523292
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1621523292
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1621523292
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1621523292
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1621523292
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1621523292
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1621523292
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1621523292
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1621523292
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1621523292
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1621523292
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1621523292
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1621523292
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1621523292
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1621523292
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1621523292
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1621523292
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1621523292
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1621523292
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1621523292
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1621523292
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1621523292
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1621523292
transform 1 0 32292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1621523292
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1621523292
transform 1 0 33396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_363
timestamp 1621523292
transform 1 0 34500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_372
timestamp 1621523292
transform 1 0 35328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_384
timestamp 1621523292
transform 1 0 36432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_396
timestamp 1621523292
transform 1 0 37536 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_408
timestamp 1621523292
transform 1 0 38640 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1621523292
transform 1 0 40480 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_420
timestamp 1621523292
transform 1 0 39744 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_429
timestamp 1621523292
transform 1 0 40572 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_441
timestamp 1621523292
transform 1 0 41676 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_453
timestamp 1621523292
transform 1 0 42780 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_465
timestamp 1621523292
transform 1 0 43884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_477
timestamp 1621523292
transform 1 0 44988 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1621523292
transform 1 0 45724 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_486
timestamp 1621523292
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_498
timestamp 1621523292
transform 1 0 46920 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_510
timestamp 1621523292
transform 1 0 48024 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_522
timestamp 1621523292
transform 1 0 49128 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1621523292
transform 1 0 50324 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1621523292
transform 1 0 50968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1621523292
transform 1 0 49680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_531
timestamp 1621523292
transform 1 0 49956 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_538
timestamp 1621523292
transform 1 0 50600 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_543
timestamp 1621523292
transform 1 0 51060 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _0851_
timestamp 1621523292
transform 1 0 51428 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0853_
timestamp 1621523292
transform 1 0 52808 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_554
timestamp 1621523292
transform 1 0 52072 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0633_
timestamp 1621523292
transform 1 0 55016 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0637_
timestamp 1621523292
transform 1 0 53912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_570
timestamp 1621523292
transform 1 0 53544 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_577
timestamp 1621523292
transform 1 0 54188 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_585
timestamp 1621523292
transform 1 0 54924 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_589
timestamp 1621523292
transform 1 0 55292 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 56672 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1621523292
transform 1 0 56212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_597
timestamp 1621523292
transform 1 0 56028 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_600
timestamp 1621523292
transform 1 0 56304 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_608
timestamp 1621523292
transform 1 0 57040 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1621523292
transform -1 0 58880 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output213
timestamp 1621523292
transform 1 0 57868 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_616
timestamp 1621523292
transform 1 0 57776 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1621523292
transform 1 0 58236 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1223_
timestamp 1621523292
transform 1 0 1840 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1621523292
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1621523292
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1621523292
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_16
timestamp 1621523292
transform 1 0 2576 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1028_
timestamp 1621523292
transform 1 0 3220 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1109_
timestamp 1621523292
transform 1 0 3864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1110_
timestamp 1621523292
transform 1 0 4508 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_22
timestamp 1621523292
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1621523292
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_33
timestamp 1621523292
transform 1 0 4140 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_40
timestamp 1621523292
transform 1 0 4784 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1621523292
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1621523292
transform 1 0 5888 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_56
timestamp 1621523292
transform 1 0 6256 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1621523292
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1621523292
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1621523292
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1621523292
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1621523292
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1621523292
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1621523292
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1621523292
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1621523292
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1621523292
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1621523292
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1621523292
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1621523292
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1621523292
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1621523292
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1621523292
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1621523292
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1621523292
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1621523292
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1621523292
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1621523292
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1621523292
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_277
timestamp 1621523292
transform 1 0 26588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1621523292
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1621523292
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_298
timestamp 1621523292
transform 1 0 28520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_310
timestamp 1621523292
transform 1 0 29624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1621523292
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1621523292
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_334
timestamp 1621523292
transform 1 0 31832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1621523292
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1621523292
transform 1 0 33764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1621523292
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1621523292
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_391
timestamp 1621523292
transform 1 0 37076 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1621523292
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_400
timestamp 1621523292
transform 1 0 37904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_412
timestamp 1621523292
transform 1 0 39008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_424
timestamp 1621523292
transform 1 0 40112 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_436
timestamp 1621523292
transform 1 0 41216 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1621523292
transform 1 0 43056 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_448
timestamp 1621523292
transform 1 0 42320 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_457
timestamp 1621523292
transform 1 0 43148 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_469
timestamp 1621523292
transform 1 0 44252 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_481
timestamp 1621523292
transform 1 0 45356 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_493
timestamp 1621523292
transform 1 0 46460 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1621523292
transform 1 0 48300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1621523292
transform 1 0 47564 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_514
timestamp 1621523292
transform 1 0 48392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0840_
timestamp 1621523292
transform 1 0 50876 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1621523292
transform 1 0 50232 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0959_
timestamp 1621523292
transform 1 0 49588 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_526
timestamp 1621523292
transform 1 0 49496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_530
timestamp 1621523292
transform 1 0 49864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_537
timestamp 1621523292
transform 1 0 50508 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_545
timestamp 1621523292
transform 1 0 51244 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_4  _0715_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52072 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_553
timestamp 1621523292
transform 1 0 51980 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_563
timestamp 1621523292
transform 1 0 52900 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1621523292
transform 1 0 54004 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1621523292
transform 1 0 53544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_569
timestamp 1621523292
transform 1 0 53452 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_571
timestamp 1621523292
transform 1 0 53636 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0876_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 55844 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _1280_
timestamp 1621523292
transform 1 0 57040 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_591
timestamp 1621523292
transform 1 0 55476 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_604
timestamp 1621523292
transform 1 0 56672 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1621523292
transform -1 0 58880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_616
timestamp 1621523292
transform 1 0 57776 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_624
timestamp 1621523292
transform 1 0 58512 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1621523292
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1621523292
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output296
timestamp 1621523292
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1621523292
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1621523292
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1224_
timestamp 1621523292
transform 1 0 1564 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1621523292
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_18
timestamp 1621523292
transform 1 0 2760 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1621523292
transform 1 0 2116 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1111_
timestamp 1621523292
transform 1 0 2668 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1621523292
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_20
timestamp 1621523292
transform 1 0 2944 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1027_
timestamp 1621523292
transform 1 0 3128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1621523292
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_25
timestamp 1621523292
transform 1 0 3404 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1621523292
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1621523292
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1621523292
transform 1 0 4048 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1621523292
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1621523292
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1621523292
transform 1 0 5152 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1621523292
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1621523292
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1621523292
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1621523292
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1621523292
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1621523292
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1621523292
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_82
timestamp 1621523292
transform 1 0 8648 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_99
timestamp 1621523292
transform 1 0 10212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_94
timestamp 1621523292
transform 1 0 9752 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_106
timestamp 1621523292
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1621523292
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_111
timestamp 1621523292
transform 1 0 11316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_123
timestamp 1621523292
transform 1 0 12420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1621523292
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1621523292
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1621523292
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_135
timestamp 1621523292
transform 1 0 13524 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1621523292
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1621523292
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1621523292
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1621523292
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1621523292
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1621523292
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1621523292
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1621523292
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1621523292
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1621523292
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1621523292
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1621523292
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1621523292
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1621523292
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1621523292
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1621523292
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1621523292
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_225
timestamp 1621523292
transform 1 0 21804 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_237
timestamp 1621523292
transform 1 0 22908 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1621523292
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1621523292
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1621523292
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_249
timestamp 1621523292
transform 1 0 24012 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1621523292
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1621523292
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_253
timestamp 1621523292
transform 1 0 24380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1621523292
transform 1 0 25944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1621523292
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_265
timestamp 1621523292
transform 1 0 25484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_277
timestamp 1621523292
transform 1 0 26588 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1621523292
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1621523292
transform 1 0 28152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1621523292
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1621523292
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1621523292
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_306
timestamp 1621523292
transform 1 0 29256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1621523292
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1621523292
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1621523292
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1621523292
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1621523292
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1621523292
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1621523292
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1621523292
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1621523292
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1621523292
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1621523292
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1621523292
transform 1 0 33764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1621523292
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1621523292
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1621523292
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1621523292
transform 1 0 35972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_391
timestamp 1621523292
transform 1 0 37076 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1621523292
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_396
timestamp 1621523292
transform 1 0 37536 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_408
timestamp 1621523292
transform 1 0 38640 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1621523292
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1621523292
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1621523292
transform 1 0 40480 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_420
timestamp 1621523292
transform 1 0 39744 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_429
timestamp 1621523292
transform 1 0 40572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1621523292
transform 1 0 40112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1621523292
transform 1 0 41216 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1621523292
transform 1 0 43056 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_441
timestamp 1621523292
transform 1 0 41676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_453
timestamp 1621523292
transform 1 0 42780 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_448
timestamp 1621523292
transform 1 0 42320 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_457
timestamp 1621523292
transform 1 0 43148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_465
timestamp 1621523292
transform 1 0 43884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_477
timestamp 1621523292
transform 1 0 44988 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_469
timestamp 1621523292
transform 1 0 44252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1621523292
transform 1 0 45724 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_486
timestamp 1621523292
transform 1 0 45816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_498
timestamp 1621523292
transform 1 0 46920 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_481
timestamp 1621523292
transform 1 0 45356 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_493
timestamp 1621523292
transform 1 0 46460 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1174_
timestamp 1621523292
transform 1 0 49036 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1621523292
transform 1 0 48300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1621523292
transform 1 0 49128 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_510
timestamp 1621523292
transform 1 0 48024 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_518
timestamp 1621523292
transform 1 0 48760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_524
timestamp 1621523292
transform 1 0 49312 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1621523292
transform 1 0 47564 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_514
timestamp 1621523292
transform 1 0 48392 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1621523292
transform 1 0 50324 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0958_
timestamp 1621523292
transform 1 0 49680 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1621523292
transform 1 0 49772 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1621523292
transform 1 0 50968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_531
timestamp 1621523292
transform 1 0 49956 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_538
timestamp 1621523292
transform 1 0 50600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_543
timestamp 1621523292
transform 1 0 51060 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_525
timestamp 1621523292
transform 1 0 49404 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_545
timestamp 1621523292
transform 1 0 51244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0709_
timestamp 1621523292
transform 1 0 51428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0843_
timestamp 1621523292
transform 1 0 52900 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0845_
timestamp 1621523292
transform 1 0 52624 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2oi_1  _0846_
timestamp 1621523292
transform 1 0 51612 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0849_
timestamp 1621523292
transform 1 0 52072 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_26_550
timestamp 1621523292
transform 1 0 51704 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_559
timestamp 1621523292
transform 1 0 52532 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_556
timestamp 1621523292
transform 1 0 52256 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_566
timestamp 1621523292
transform 1 0 53176 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_575
timestamp 1621523292
transform 1 0 54004 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_571
timestamp 1621523292
transform 1 0 53636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_577
timestamp 1621523292
transform 1 0 54188 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_570
timestamp 1621523292
transform 1 0 53544 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1621523292
transform 1 0 53544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1621523292
transform 1 0 53912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_584
timestamp 1621523292
transform 1 0 54832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1621523292
transform 1 0 55200 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1621523292
transform 1 0 54556 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1621523292
transform 1 0 54096 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_1  _0708_
timestamp 1621523292
transform 1 0 55936 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1621523292
transform 1 0 56672 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1621523292
transform 1 0 56212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output215
timestamp 1621523292
transform 1 0 57132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_591
timestamp 1621523292
transform 1 0 55476 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_600
timestamp 1621523292
transform 1 0 56304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_608
timestamp 1621523292
transform 1 0 57040 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_592
timestamp 1621523292
transform 1 0 55568 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_603
timestamp 1621523292
transform 1 0 56580 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _1318_
timestamp 1621523292
transform 1 0 57500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1621523292
transform -1 0 58880 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1621523292
transform -1 0 58880 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output177
timestamp 1621523292
transform 1 0 57868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_612
timestamp 1621523292
transform 1 0 57408 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1621523292
transform 1 0 58236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_613
timestamp 1621523292
transform 1 0 57500 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1621523292
transform 1 0 58236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1024_
timestamp 1621523292
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1621523292
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output297
timestamp 1621523292
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1621523292
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_11
timestamp 1621523292
transform 1 0 2116 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1621523292
transform 1 0 2760 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1621523292
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1621523292
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1621523292
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1621523292
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1621523292
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1621523292
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1621523292
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1621523292
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1621523292
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1621523292
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1621523292
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1621523292
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1621523292
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1621523292
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1621523292
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1621523292
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1621523292
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1621523292
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1621523292
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1621523292
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1621523292
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_213
timestamp 1621523292
transform 1 0 20700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1621523292
transform 1 0 21804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1621523292
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1621523292
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1621523292
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1621523292
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_270
timestamp 1621523292
transform 1 0 25944 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_282
timestamp 1621523292
transform 1 0 27048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_294
timestamp 1621523292
transform 1 0 28152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1621523292
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_306
timestamp 1621523292
transform 1 0 29256 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1621523292
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1621523292
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1621523292
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1621523292
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1621523292
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1621523292
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1621523292
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1621523292
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_396
timestamp 1621523292
transform 1 0 37536 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_408
timestamp 1621523292
transform 1 0 38640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1621523292
transform 1 0 40480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_420
timestamp 1621523292
transform 1 0 39744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_429
timestamp 1621523292
transform 1 0 40572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_441
timestamp 1621523292
transform 1 0 41676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_453
timestamp 1621523292
transform 1 0 42780 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_465
timestamp 1621523292
transform 1 0 43884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 1621523292
transform 1 0 44988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1621523292
transform 1 0 45724 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_486
timestamp 1621523292
transform 1 0 45816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_498
timestamp 1621523292
transform 1 0 46920 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1175_
timestamp 1621523292
transform 1 0 49036 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_510
timestamp 1621523292
transform 1 0 48024 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_518
timestamp 1621523292
transform 1 0 48760 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_524
timestamp 1621523292
transform 1 0 49312 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 1621523292
transform 1 0 50324 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0912_
timestamp 1621523292
transform 1 0 49680 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1621523292
transform 1 0 50968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_531
timestamp 1621523292
transform 1 0 49956 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_538
timestamp 1621523292
transform 1 0 50600 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_543
timestamp 1621523292
transform 1 0 51060 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0706_
timestamp 1621523292
transform 1 0 51428 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0750_
timestamp 1621523292
transform 1 0 52440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_554
timestamp 1621523292
transform 1 0 52072 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_567
timestamp 1621523292
transform 1 0 53268 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0632_
timestamp 1621523292
transform 1 0 54740 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0848_
timestamp 1621523292
transform 1 0 53636 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_579
timestamp 1621523292
transform 1 0 54372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_586
timestamp 1621523292
transform 1 0 55016 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0631_
timestamp 1621523292
transform 1 0 55476 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1281_
timestamp 1621523292
transform 1 0 56948 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1621523292
transform 1 0 56212 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_590
timestamp 1621523292
transform 1 0 55384 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_594
timestamp 1621523292
transform 1 0 55752 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_598
timestamp 1621523292
transform 1 0 56120 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_600
timestamp 1621523292
transform 1 0 56304 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_606
timestamp 1621523292
transform 1 0 56856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1621523292
transform -1 0 58880 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_615
timestamp 1621523292
transform 1 0 57684 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_623
timestamp 1621523292
transform 1 0 58420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _1112_
timestamp 1621523292
transform 1 0 2668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1225_
timestamp 1621523292
transform 1 0 1564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1621523292
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1621523292
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1621523292
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1621523292
transform 1 0 2944 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1621523292
transform 1 0 4048 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1621523292
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1621523292
transform 1 0 5152 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_56
timestamp 1621523292
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1621523292
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1621523292
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1621523292
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1621523292
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1621523292
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1621523292
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1621523292
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1621523292
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1621523292
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1621523292
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1621523292
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1621523292
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1621523292
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1621523292
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1621523292
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1621523292
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1621523292
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1621523292
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1621523292
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1621523292
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1621523292
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1621523292
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1621523292
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1621523292
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1621523292
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_298
timestamp 1621523292
transform 1 0 28520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_310
timestamp 1621523292
transform 1 0 29624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1621523292
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1621523292
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1621523292
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1621523292
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_355
timestamp 1621523292
transform 1 0 33764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1621523292
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1621523292
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_391
timestamp 1621523292
transform 1 0 37076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1621523292
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1621523292
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_412
timestamp 1621523292
transform 1 0 39008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1621523292
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1621523292
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1621523292
transform 1 0 43056 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_448
timestamp 1621523292
transform 1 0 42320 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_457
timestamp 1621523292
transform 1 0 43148 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_469
timestamp 1621523292
transform 1 0 44252 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_481
timestamp 1621523292
transform 1 0 45356 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_493
timestamp 1621523292
transform 1 0 46460 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1621523292
transform 1 0 48300 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1621523292
transform 1 0 47564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_514
timestamp 1621523292
transform 1 0 48392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0629_
timestamp 1621523292
transform 1 0 51244 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0911_
timestamp 1621523292
transform 1 0 50600 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1068_
timestamp 1621523292
transform 1 0 49956 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_526
timestamp 1621523292
transform 1 0 49496 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_530
timestamp 1621523292
transform 1 0 49864 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_534
timestamp 1621523292
transform 1 0 50232 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_541
timestamp 1621523292
transform 1 0 50876 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0630_
timestamp 1621523292
transform 1 0 51888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0749_
timestamp 1621523292
transform 1 0 52532 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_548
timestamp 1621523292
transform 1 0 51520 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_555
timestamp 1621523292
transform 1 0 52164 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_566
timestamp 1621523292
transform 1 0 53176 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0834_
timestamp 1621523292
transform 1 0 54004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1621523292
transform 1 0 54740 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1621523292
transform 1 0 53544 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_571
timestamp 1621523292
transform 1 0 53636 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_578
timestamp 1621523292
transform 1 0 54280 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_582
timestamp 1621523292
transform 1 0 54648 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output216
timestamp 1621523292
transform 1 0 56764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_599
timestamp 1621523292
transform 1 0 56212 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_609
timestamp 1621523292
transform 1 0 57132 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1319_
timestamp 1621523292
transform 1 0 57500 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1621523292
transform -1 0 58880 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1621523292
transform 1 0 58236 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1023_
timestamp 1621523292
transform 1 0 3036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1226_
timestamp 1621523292
transform 1 0 1932 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1621523292
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_3
timestamp 1621523292
transform 1 0 1380 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_17
timestamp 1621523292
transform 1 0 2668 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1621523292
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1621523292
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1621523292
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1621523292
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1621523292
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1621523292
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1621523292
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1621523292
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1621523292
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1621523292
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1621523292
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1621523292
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1621523292
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1621523292
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1621523292
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1621523292
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1621523292
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1621523292
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1621523292
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1621523292
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1621523292
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1621523292
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1621523292
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1621523292
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1621523292
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1621523292
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1621523292
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1621523292
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_270
timestamp 1621523292
transform 1 0 25944 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_282
timestamp 1621523292
transform 1 0 27048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_294
timestamp 1621523292
transform 1 0 28152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1621523292
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_306
timestamp 1621523292
transform 1 0 29256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_315
timestamp 1621523292
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1621523292
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1621523292
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1621523292
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1621523292
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1621523292
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1621523292
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1621523292
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1621523292
transform 1 0 37536 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1621523292
transform 1 0 38640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1621523292
transform 1 0 40480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_420
timestamp 1621523292
transform 1 0 39744 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_429
timestamp 1621523292
transform 1 0 40572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_441
timestamp 1621523292
transform 1 0 41676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_453
timestamp 1621523292
transform 1 0 42780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_465
timestamp 1621523292
transform 1 0 43884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1621523292
transform 1 0 44988 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1621523292
transform 1 0 45724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_486
timestamp 1621523292
transform 1 0 45816 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_498
timestamp 1621523292
transform 1 0 46920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 49036 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_510
timestamp 1621523292
transform 1 0 48024 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_518
timestamp 1621523292
transform 1 0 48760 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_524
timestamp 1621523292
transform 1 0 49312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1069_
timestamp 1621523292
transform 1 0 50324 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1621523292
transform 1 0 50968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1621523292
transform 1 0 49680 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_531
timestamp 1621523292
transform 1 0 49956 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_538
timestamp 1621523292
transform 1 0 50600 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_543
timestamp 1621523292
transform 1 0 51060 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1621523292
transform 1 0 51612 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0826_
timestamp 1621523292
transform 1 0 52348 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_30_552
timestamp 1621523292
transform 1 0 51888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_556
timestamp 1621523292
transform 1 0 52256 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_564
timestamp 1621523292
transform 1 0 52992 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0701_
timestamp 1621523292
transform 1 0 53912 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1621523292
transform 1 0 54924 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_572
timestamp 1621523292
transform 1 0 53728 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_581
timestamp 1621523292
transform 1 0 54556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_588
timestamp 1621523292
transform 1 0 55200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0707_
timestamp 1621523292
transform 1 0 55568 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1054_
timestamp 1621523292
transform 1 0 56672 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1621523292
transform 1 0 56212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_595
timestamp 1621523292
transform 1 0 55844 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_600
timestamp 1621523292
transform 1 0 56304 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_608
timestamp 1621523292
transform 1 0 57040 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1621523292
transform -1 0 58880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output178
timestamp 1621523292
transform 1 0 57868 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_616
timestamp 1621523292
transform 1 0 57776 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1621523292
transform 1 0 58236 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1621523292
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output298
timestamp 1621523292
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output300
timestamp 1621523292
transform 1 0 2484 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1621523292
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1621523292
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_19
timestamp 1621523292
transform 1 0 2852 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1113_
timestamp 1621523292
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_26
timestamp 1621523292
transform 1 0 3496 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_38
timestamp 1621523292
transform 1 0 4600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1621523292
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1621523292
transform 1 0 5704 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_56
timestamp 1621523292
transform 1 0 6256 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1621523292
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1621523292
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_82
timestamp 1621523292
transform 1 0 8648 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_94
timestamp 1621523292
transform 1 0 9752 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_106
timestamp 1621523292
transform 1 0 10856 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1621523292
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1621523292
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1621523292
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1621523292
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1621523292
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1621523292
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1621523292
transform 1 0 16100 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1621523292
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1621523292
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1621523292
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1621523292
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1621523292
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1621523292
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1621523292
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1621523292
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1621523292
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1621523292
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1621523292
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1621523292
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1621523292
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1621523292
transform 1 0 28520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1621523292
transform 1 0 29624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1621523292
transform 1 0 30728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1621523292
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1621523292
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1621523292
transform 1 0 32660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1621523292
transform 1 0 33764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1621523292
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1621523292
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_391
timestamp 1621523292
transform 1 0 37076 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1621523292
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1621523292
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1621523292
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1621523292
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1621523292
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1621523292
transform 1 0 43056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_448
timestamp 1621523292
transform 1 0 42320 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_457
timestamp 1621523292
transform 1 0 43148 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_469
timestamp 1621523292
transform 1 0 44252 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_481
timestamp 1621523292
transform 1 0 45356 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_493
timestamp 1621523292
transform 1 0 46460 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1621523292
transform 1 0 48300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 48944 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1621523292
transform 1 0 47656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_505
timestamp 1621523292
transform 1 0 47564 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_509
timestamp 1621523292
transform 1 0 47932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_514
timestamp 1621523292
transform 1 0 48392 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_523
timestamp 1621523292
transform 1 0 49220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0910_
timestamp 1621523292
transform 1 0 49588 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1621523292
transform 1 0 50232 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_530
timestamp 1621523292
transform 1 0 49864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0839_
timestamp 1621523292
transform 1 0 52440 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_550
timestamp 1621523292
transform 1 0 51704 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_566
timestamp 1621523292
transform 1 0 53176 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1621523292
transform 1 0 54280 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1621523292
transform 1 0 54924 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1621523292
transform 1 0 53544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_571
timestamp 1621523292
transform 1 0 53636 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_577
timestamp 1621523292
transform 1 0 54188 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_581
timestamp 1621523292
transform 1 0 54556 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1282_
timestamp 1621523292
transform 1 0 56948 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_601
timestamp 1621523292
transform 1 0 56396 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1621523292
transform -1 0 58880 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_615
timestamp 1621523292
transform 1 0 57684 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1621523292
transform 1 0 58420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1019_
timestamp 1621523292
transform 1 0 2852 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1227_
timestamp 1621523292
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1621523292
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1621523292
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_15
timestamp 1621523292
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1114_
timestamp 1621523292
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1621523292
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1621523292
transform 1 0 3128 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_28
timestamp 1621523292
transform 1 0 3680 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_30
timestamp 1621523292
transform 1 0 3864 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_37
timestamp 1621523292
transform 1 0 4508 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_49
timestamp 1621523292
transform 1 0 5612 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_61
timestamp 1621523292
transform 1 0 6716 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1621523292
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_73
timestamp 1621523292
transform 1 0 7820 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1621523292
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1621523292
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1621523292
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1621523292
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1621523292
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1621523292
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1621523292
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1621523292
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1621523292
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1621523292
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_180
timestamp 1621523292
transform 1 0 17664 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1621523292
transform 1 0 18768 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1621523292
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1621523292
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1621523292
transform 1 0 20700 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1621523292
transform 1 0 21804 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_237
timestamp 1621523292
transform 1 0 22908 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1621523292
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_249
timestamp 1621523292
transform 1 0 24012 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1621523292
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1621523292
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1621523292
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1621523292
transform 1 0 28152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1621523292
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_306
timestamp 1621523292
transform 1 0 29256 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_315
timestamp 1621523292
transform 1 0 30084 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_327
timestamp 1621523292
transform 1 0 31188 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_339
timestamp 1621523292
transform 1 0 32292 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1621523292
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_351
timestamp 1621523292
transform 1 0 33396 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_363
timestamp 1621523292
transform 1 0 34500 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1621523292
transform 1 0 35328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1621523292
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_396
timestamp 1621523292
transform 1 0 37536 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_408
timestamp 1621523292
transform 1 0 38640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1621523292
transform 1 0 40480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_420
timestamp 1621523292
transform 1 0 39744 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_429
timestamp 1621523292
transform 1 0 40572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_441
timestamp 1621523292
transform 1 0 41676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_453
timestamp 1621523292
transform 1 0 42780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1621523292
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_477
timestamp 1621523292
transform 1 0 44988 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1621523292
transform 1 0 45724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_486
timestamp 1621523292
transform 1 0 45816 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_498
timestamp 1621523292
transform 1 0 46920 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 49036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_510
timestamp 1621523292
transform 1 0 48024 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_518
timestamp 1621523292
transform 1 0 48760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_524
timestamp 1621523292
transform 1 0 49312 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0956_
timestamp 1621523292
transform 1 0 50324 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1176_
timestamp 1621523292
transform 1 0 49680 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1621523292
transform 1 0 50968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_531
timestamp 1621523292
transform 1 0 49956 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_538
timestamp 1621523292
transform 1 0 50600 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_543
timestamp 1621523292
transform 1 0 51060 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0623_
timestamp 1621523292
transform 1 0 51428 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0835_
timestamp 1621523292
transform 1 0 52164 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1621523292
transform 1 0 53084 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_551
timestamp 1621523292
transform 1 0 51796 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_561
timestamp 1621523292
transform 1 0 52716 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0628_
timestamp 1621523292
transform 1 0 54924 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_581
timestamp 1621523292
transform 1 0 54556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_588
timestamp 1621523292
transform 1 0 55200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0700_
timestamp 1621523292
transform 1 0 55568 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1621523292
transform 1 0 56212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output217
timestamp 1621523292
transform 1 0 56764 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_595
timestamp 1621523292
transform 1 0 55844 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_600
timestamp 1621523292
transform 1 0 56304 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_604
timestamp 1621523292
transform 1 0 56672 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_609
timestamp 1621523292
transform 1 0 57132 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1320_
timestamp 1621523292
transform 1 0 57500 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1621523292
transform -1 0 58880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1621523292
transform 1 0 58236 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1621523292
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1621523292
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output301
timestamp 1621523292
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1621523292
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1621523292
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1228_
timestamp 1621523292
transform 1 0 1748 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1621523292
transform 1 0 2116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1621523292
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output302
timestamp 1621523292
transform 1 0 2484 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1621523292
transform 1 0 2852 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1020_
timestamp 1621523292
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1022_
timestamp 1621523292
transform 1 0 3864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1621523292
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1621523292
transform 1 0 3496 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_33
timestamp 1621523292
transform 1 0 4140 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1621523292
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1621523292
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1621523292
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1621523292
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_45
timestamp 1621523292
transform 1 0 5244 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1621523292
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1621523292
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1621523292
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1621523292
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1621523292
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1621523292
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1621523292
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1621523292
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1621523292
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1621523292
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1621523292
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1621523292
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1621523292
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1621523292
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1621523292
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1621523292
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1621523292
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1621523292
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1621523292
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1621523292
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1621523292
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1621523292
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1621523292
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1621523292
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1621523292
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1621523292
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1621523292
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1621523292
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1621523292
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1621523292
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1621523292
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1621523292
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_201
timestamp 1621523292
transform 1 0 19596 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_213
timestamp 1621523292
transform 1 0 20700 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1621523292
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1621523292
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_229
timestamp 1621523292
transform 1 0 22172 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_225
timestamp 1621523292
transform 1 0 21804 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_237
timestamp 1621523292
transform 1 0 22908 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1621523292
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_241
timestamp 1621523292
transform 1 0 23276 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_253
timestamp 1621523292
transform 1 0 24380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1621523292
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1621523292
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_265
timestamp 1621523292
transform 1 0 25484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_277
timestamp 1621523292
transform 1 0 26588 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1621523292
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_282
timestamp 1621523292
transform 1 0 27048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1621523292
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1621523292
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_298
timestamp 1621523292
transform 1 0 28520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_294
timestamp 1621523292
transform 1 0 28152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1621523292
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1621523292
transform 1 0 29624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_322
timestamp 1621523292
transform 1 0 30728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_306
timestamp 1621523292
transform 1 0 29256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_315
timestamp 1621523292
transform 1 0 30084 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_327
timestamp 1621523292
transform 1 0 31188 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1621523292
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_334
timestamp 1621523292
transform 1 0 31832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1621523292
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_339
timestamp 1621523292
transform 1 0 32292 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1621523292
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1621523292
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1621523292
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_351
timestamp 1621523292
transform 1 0 33396 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_363
timestamp 1621523292
transform 1 0 34500 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1621523292
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1621523292
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_372
timestamp 1621523292
transform 1 0 35328 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_384
timestamp 1621523292
transform 1 0 36432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1621523292
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_400
timestamp 1621523292
transform 1 0 37904 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_412
timestamp 1621523292
transform 1 0 39008 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_396
timestamp 1621523292
transform 1 0 37536 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_408
timestamp 1621523292
transform 1 0 38640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1621523292
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_424
timestamp 1621523292
transform 1 0 40112 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_436
timestamp 1621523292
transform 1 0 41216 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_420
timestamp 1621523292
transform 1 0 39744 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1621523292
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1621523292
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_448
timestamp 1621523292
transform 1 0 42320 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1621523292
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1621523292
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1621523292
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1621523292
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_465
timestamp 1621523292
transform 1 0 43884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1621523292
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1621523292
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1621523292
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_493
timestamp 1621523292
transform 1 0 46460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1621523292
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_498
timestamp 1621523292
transform 1 0 46920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_510
timestamp 1621523292
transform 1 0 48024 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1621523292
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_517
timestamp 1621523292
transform 1 0 48668 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_514
timestamp 1621523292
transform 1 0 48392 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1621523292
transform 1 0 48392 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1621523292
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_524
timestamp 1621523292
transform 1 0 49312 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_524
timestamp 1621523292
transform 1 0 49312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_520
timestamp 1621523292
transform 1 0 48944 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 49036 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1621523292
transform 1 0 49036 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_531
timestamp 1621523292
transform 1 0 49956 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_531
timestamp 1621523292
transform 1 0 49956 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1177_
timestamp 1621523292
transform 1 0 49680 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0909_
timestamp 1621523292
transform 1 0 49680 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_538
timestamp 1621523292
transform 1 0 50600 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_538
timestamp 1621523292
transform 1 0 50600 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0955_
timestamp 1621523292
transform 1 0 50324 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0837_
timestamp 1621523292
transform 1 0 50324 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_543
timestamp 1621523292
transform 1 0 51060 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1621523292
transform 1 0 50968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _0836_
timestamp 1621523292
transform 1 0 50968 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _0704_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52532 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0827_
timestamp 1621523292
transform 1 0 51888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0828_
timestamp 1621523292
transform 1 0 52532 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_33_549
timestamp 1621523292
transform 1 0 51612 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_557
timestamp 1621523292
transform 1 0 52348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_566
timestamp 1621523292
transform 1 0 53176 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_551
timestamp 1621523292
transform 1 0 51796 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_555
timestamp 1621523292
transform 1 0 52164 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_568
timestamp 1621523292
transform 1 0 53360 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_577
timestamp 1621523292
transform 1 0 54188 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_571
timestamp 1621523292
transform 1 0 53636 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1621523292
transform 1 0 53544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _0753_
timestamp 1621523292
transform 1 0 53728 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_581
timestamp 1621523292
transform 1 0 54556 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_585
timestamp 1621523292
transform 1 0 54924 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0745_
timestamp 1621523292
transform 1 0 54280 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _0703_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 54924 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1621523292
transform 1 0 55292 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_593
timestamp 1621523292
transform 1 0 55660 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_596
timestamp 1621523292
transform 1 0 55936 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_592
timestamp 1621523292
transform 1 0 55568 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1621523292
transform 1 0 56028 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_600
timestamp 1621523292
transform 1 0 56304 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_600
timestamp 1621523292
transform 1 0 56304 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1621523292
transform 1 0 56212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_608
timestamp 1621523292
transform 1 0 57040 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output218
timestamp 1621523292
transform 1 0 57132 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1283_
timestamp 1621523292
transform 1 0 57040 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1621523292
transform -1 0 58880 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1621523292
transform -1 0 58880 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output179
timestamp 1621523292
transform 1 0 57868 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_613
timestamp 1621523292
transform 1 0 57500 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_621
timestamp 1621523292
transform 1 0 58236 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_616
timestamp 1621523292
transform 1 0 57776 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_624
timestamp 1621523292
transform 1 0 58512 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1021_
timestamp 1621523292
transform 1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1229_
timestamp 1621523292
transform 1 0 1656 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1621523292
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1621523292
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1621523292
transform 1 0 2392 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1621523292
transform 1 0 3036 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1115_
timestamp 1621523292
transform 1 0 3404 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1116_
timestamp 1621523292
transform 1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_28
timestamp 1621523292
transform 1 0 3680 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_35
timestamp 1621523292
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1621523292
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_47
timestamp 1621523292
transform 1 0 5428 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_55
timestamp 1621523292
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1621523292
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1621523292
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1621523292
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1621523292
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1621523292
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1621523292
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1621523292
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1621523292
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1621523292
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1621523292
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1621523292
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1621523292
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1621523292
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1621523292
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1621523292
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1621523292
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1621523292
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_220
timestamp 1621523292
transform 1 0 21344 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1621523292
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1621523292
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1621523292
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1621523292
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1621523292
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1621523292
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1621523292
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_298
timestamp 1621523292
transform 1 0 28520 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_310
timestamp 1621523292
transform 1 0 29624 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_322
timestamp 1621523292
transform 1 0 30728 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1621523292
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_334
timestamp 1621523292
transform 1 0 31832 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1621523292
transform 1 0 32660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_355
timestamp 1621523292
transform 1 0 33764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1621523292
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1621523292
transform 1 0 35972 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_391
timestamp 1621523292
transform 1 0 37076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1621523292
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_400
timestamp 1621523292
transform 1 0 37904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_412
timestamp 1621523292
transform 1 0 39008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_424
timestamp 1621523292
transform 1 0 40112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1621523292
transform 1 0 41216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1621523292
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_448
timestamp 1621523292
transform 1 0 42320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_457
timestamp 1621523292
transform 1 0 43148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_469
timestamp 1621523292
transform 1 0 44252 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1621523292
transform 1 0 45356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_493
timestamp 1621523292
transform 1 0 46460 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1621523292
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1621523292
transform 1 0 47564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_514
timestamp 1621523292
transform 1 0 48392 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1621523292
transform 1 0 49864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1621523292
transform 1 0 50508 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_526
timestamp 1621523292
transform 1 0 49496 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_533
timestamp 1621523292
transform 1 0 50140 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _0754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52348 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_553
timestamp 1621523292
transform 1 0 51980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_565
timestamp 1621523292
transform 1 0 53084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0746_
timestamp 1621523292
transform 1 0 54188 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1621523292
transform 1 0 55108 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1621523292
transform 1 0 53544 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_569
timestamp 1621523292
transform 1 0 53452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_571
timestamp 1621523292
transform 1 0 53636 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_581
timestamp 1621523292
transform 1 0 54556 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_603
timestamp 1621523292
transform 1 0 56580 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_611
timestamp 1621523292
transform 1 0 57316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _1321_
timestamp 1621523292
transform 1 0 57500 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1621523292
transform -1 0 58880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1621523292
transform 1 0 58236 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1007_
timestamp 1621523292
transform 1 0 2484 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1621523292
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output303
timestamp 1621523292
transform 1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1621523292
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_11
timestamp 1621523292
transform 1 0 2116 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_21
timestamp 1621523292
transform 1 0 3036 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1621523292
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1621523292
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1621523292
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1621523292
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1621523292
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1621523292
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1621523292
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1621523292
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1621523292
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1621523292
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1621523292
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1621523292
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1621523292
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1621523292
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1621523292
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1621523292
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1621523292
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1621523292
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1621523292
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1621523292
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1621523292
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1621523292
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1621523292
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1621523292
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1621523292
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1621523292
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1621523292
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_282
timestamp 1621523292
transform 1 0 27048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_294
timestamp 1621523292
transform 1 0 28152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1621523292
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_306
timestamp 1621523292
transform 1 0 29256 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1621523292
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1621523292
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1621523292
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1621523292
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1621523292
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1621523292
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_372
timestamp 1621523292
transform 1 0 35328 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_384
timestamp 1621523292
transform 1 0 36432 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_396
timestamp 1621523292
transform 1 0 37536 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_408
timestamp 1621523292
transform 1 0 38640 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1621523292
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_420
timestamp 1621523292
transform 1 0 39744 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1621523292
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1621523292
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_453
timestamp 1621523292
transform 1 0 42780 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_465
timestamp 1621523292
transform 1 0 43884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1621523292
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1621523292
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1621523292
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1621523292
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 49036 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_510
timestamp 1621523292
transform 1 0 48024 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_518
timestamp 1621523292
transform 1 0 48760 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_524
timestamp 1621523292
transform 1 0 49312 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1178_
timestamp 1621523292
transform 1 0 50324 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1621523292
transform 1 0 50968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1621523292
transform 1 0 49680 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_531
timestamp 1621523292
transform 1 0 49956 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_538
timestamp 1621523292
transform 1 0 50600 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_543
timestamp 1621523292
transform 1 0 51060 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 1621523292
transform 1 0 52624 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0808_
timestamp 1621523292
transform 1 0 51428 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_551
timestamp 1621523292
transform 1 0 51796 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_559
timestamp 1621523292
transform 1 0 52532 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_563
timestamp 1621523292
transform 1 0 52900 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0624_
timestamp 1621523292
transform 1 0 54832 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0698_
timestamp 1621523292
transform 1 0 53820 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_36_571
timestamp 1621523292
transform 1 0 53636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_580
timestamp 1621523292
transform 1 0 54464 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_587
timestamp 1621523292
transform 1 0 55108 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0626_
timestamp 1621523292
transform 1 0 55476 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1621523292
transform 1 0 56212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output180
timestamp 1621523292
transform 1 0 56764 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_594
timestamp 1621523292
transform 1 0 55752 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_598
timestamp 1621523292
transform 1 0 56120 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_600
timestamp 1621523292
transform 1 0 56304 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_604
timestamp 1621523292
transform 1 0 56672 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_609
timestamp 1621523292
transform 1 0 57132 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1322_
timestamp 1621523292
transform 1 0 57500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1621523292
transform -1 0 58880 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_621
timestamp 1621523292
transform 1 0 58236 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1013_
timestamp 1621523292
transform 1 0 2668 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1230_
timestamp 1621523292
transform 1 0 1564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1621523292
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1621523292
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_13
timestamp 1621523292
transform 1 0 2300 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_20
timestamp 1621523292
transform 1 0 2944 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1018_
timestamp 1621523292
transform 1 0 3312 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1621523292
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1621523292
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1621523292
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_51
timestamp 1621523292
transform 1 0 5796 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1621523292
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1621523292
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1621523292
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1621523292
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1621523292
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1621523292
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1621523292
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1621523292
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1621523292
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1621523292
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1621523292
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1621523292
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1621523292
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1621523292
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1621523292
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1621523292
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1621523292
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_220
timestamp 1621523292
transform 1 0 21344 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1621523292
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1621523292
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1621523292
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_265
timestamp 1621523292
transform 1 0 25484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_277
timestamp 1621523292
transform 1 0 26588 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1621523292
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1621523292
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1621523292
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1621523292
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1621523292
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1621523292
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1621523292
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1621523292
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1621523292
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1621523292
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1621523292
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_391
timestamp 1621523292
transform 1 0 37076 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1621523292
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1621523292
transform 1 0 37904 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1621523292
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_424
timestamp 1621523292
transform 1 0 40112 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_436
timestamp 1621523292
transform 1 0 41216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1621523292
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_448
timestamp 1621523292
transform 1 0 42320 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1621523292
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1621523292
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_481
timestamp 1621523292
transform 1 0 45356 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_493
timestamp 1621523292
transform 1 0 46460 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1621523292
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1621523292
transform 1 0 47564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_514
timestamp 1621523292
transform 1 0 48392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0954_
timestamp 1621523292
transform 1 0 50784 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1071_
timestamp 1621523292
transform 1 0 50140 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_526
timestamp 1621523292
transform 1 0 49496 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_532
timestamp 1621523292
transform 1 0 50048 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_536
timestamp 1621523292
transform 1 0 50416 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_543
timestamp 1621523292
transform 1 0 51060 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 1621523292
transform 1 0 51428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0833_
timestamp 1621523292
transform 1 0 52072 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_550
timestamp 1621523292
transform 1 0 51704 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_562
timestamp 1621523292
transform 1 0 52808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1621523292
transform 1 0 54096 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1621523292
transform 1 0 54832 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1621523292
transform 1 0 53544 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_571
timestamp 1621523292
transform 1 0 53636 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_575
timestamp 1621523292
transform 1 0 54004 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_579
timestamp 1621523292
transform 1 0 54372 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_583
timestamp 1621523292
transform 1 0 54740 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1284_
timestamp 1621523292
transform 1 0 56948 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_600
timestamp 1621523292
transform 1 0 56304 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_606
timestamp 1621523292
transform 1 0 56856 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1621523292
transform -1 0 58880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_615
timestamp 1621523292
transform 1 0 57684 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1621523292
transform 1 0 58420 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1017_
timestamp 1621523292
transform 1 0 2484 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1621523292
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output304
timestamp 1621523292
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1621523292
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1621523292
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_18
timestamp 1621523292
transform 1 0 2760 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1117_
timestamp 1621523292
transform 1 0 3128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1621523292
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_25
timestamp 1621523292
transform 1 0 3404 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_30
timestamp 1621523292
transform 1 0 3864 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_42
timestamp 1621523292
transform 1 0 4968 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_54
timestamp 1621523292
transform 1 0 6072 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1621523292
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_66
timestamp 1621523292
transform 1 0 7176 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_78
timestamp 1621523292
transform 1 0 8280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1621523292
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1621523292
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1621523292
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1621523292
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1621523292
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1621523292
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1621523292
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1621523292
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1621523292
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1621523292
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1621523292
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1621523292
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_201
timestamp 1621523292
transform 1 0 19596 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_213
timestamp 1621523292
transform 1 0 20700 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_225
timestamp 1621523292
transform 1 0 21804 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_237
timestamp 1621523292
transform 1 0 22908 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1621523292
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_249
timestamp 1621523292
transform 1 0 24012 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1621523292
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1621523292
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_282
timestamp 1621523292
transform 1 0 27048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_294
timestamp 1621523292
transform 1 0 28152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1621523292
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_306
timestamp 1621523292
transform 1 0 29256 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1621523292
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1621523292
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1621523292
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1621523292
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1621523292
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1621523292
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1621523292
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1621523292
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_396
timestamp 1621523292
transform 1 0 37536 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_408
timestamp 1621523292
transform 1 0 38640 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1621523292
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_420
timestamp 1621523292
transform 1 0 39744 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1621523292
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1621523292
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1621523292
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1621523292
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1621523292
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1621523292
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1621523292
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_498
timestamp 1621523292
transform 1 0 46920 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_510
timestamp 1621523292
transform 1 0 48024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_522
timestamp 1621523292
transform 1 0 49128 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1072_
timestamp 1621523292
transform 1 0 50324 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1621523292
transform 1 0 50968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_534
timestamp 1621523292
transform 1 0 50232 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_538
timestamp 1621523292
transform 1 0 50600 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_543
timestamp 1621523292
transform 1 0 51060 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1621523292
transform 1 0 51520 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1621523292
transform 1 0 52164 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_38_547
timestamp 1621523292
transform 1 0 51428 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_551
timestamp 1621523292
transform 1 0 51796 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0752_
timestamp 1621523292
transform 1 0 54280 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_571
timestamp 1621523292
transform 1 0 53636 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_577
timestamp 1621523292
transform 1 0 54188 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_586
timestamp 1621523292
transform 1 0 55016 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1621523292
transform 1 0 55568 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1285_
timestamp 1621523292
transform 1 0 57132 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1621523292
transform 1 0 56212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_595
timestamp 1621523292
transform 1 0 55844 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_600
timestamp 1621523292
transform 1 0 56304 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_608
timestamp 1621523292
transform 1 0 57040 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1621523292
transform -1 0 58880 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_617
timestamp 1621523292
transform 1 0 57868 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1621523292
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1621523292
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1621523292
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1621523292
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1232_
timestamp 1621523292
transform 1 0 1656 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1231_
timestamp 1621523292
transform 1 0 1656 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_21
timestamp 1621523292
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_14
timestamp 1621523292
transform 1 0 2392 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1621523292
transform 1 0 2392 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1119_
timestamp 1621523292
transform 1 0 2760 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1118_
timestamp 1621523292
transform 1 0 2760 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_21
timestamp 1621523292
transform 1 0 3036 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1621523292
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_33
timestamp 1621523292
transform 1 0 4140 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1621523292
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1621523292
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1621523292
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_45
timestamp 1621523292
transform 1 0 5244 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1621523292
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1621523292
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1621523292
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1621523292
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1621523292
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1621523292
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1621523292
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1621523292
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1621523292
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1621523292
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1621523292
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1621523292
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1621523292
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1621523292
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1621523292
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1621523292
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1621523292
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1621523292
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1621523292
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1621523292
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1621523292
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1621523292
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1621523292
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1621523292
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1621523292
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1621523292
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1621523292
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1621523292
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1621523292
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1621523292
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1621523292
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1621523292
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1621523292
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1621523292
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1621523292
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1621523292
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_229
timestamp 1621523292
transform 1 0 22172 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_225
timestamp 1621523292
transform 1 0 21804 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1621523292
transform 1 0 22908 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1621523292
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_241
timestamp 1621523292
transform 1 0 23276 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_253
timestamp 1621523292
transform 1 0 24380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_249
timestamp 1621523292
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1621523292
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_265
timestamp 1621523292
transform 1 0 25484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_277
timestamp 1621523292
transform 1 0 26588 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1621523292
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1621523292
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1621523292
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_286
timestamp 1621523292
transform 1 0 27416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1621523292
transform 1 0 28520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_294
timestamp 1621523292
transform 1 0 28152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1621523292
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_310
timestamp 1621523292
transform 1 0 29624 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_322
timestamp 1621523292
transform 1 0 30728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_306
timestamp 1621523292
transform 1 0 29256 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1621523292
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1621523292
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1621523292
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_334
timestamp 1621523292
transform 1 0 31832 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1621523292
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1621523292
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1621523292
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1621523292
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1621523292
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1621523292
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1621523292
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1621523292
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1621523292
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_372
timestamp 1621523292
transform 1 0 35328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1621523292
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1621523292
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1621523292
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1621523292
transform 1 0 39008 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_396
timestamp 1621523292
transform 1 0 37536 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_408
timestamp 1621523292
transform 1 0 38640 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1621523292
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_424
timestamp 1621523292
transform 1 0 40112 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_436
timestamp 1621523292
transform 1 0 41216 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_420
timestamp 1621523292
transform 1 0 39744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_429
timestamp 1621523292
transform 1 0 40572 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1621523292
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_448
timestamp 1621523292
transform 1 0 42320 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1621523292
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_441
timestamp 1621523292
transform 1 0 41676 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_453
timestamp 1621523292
transform 1 0 42780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1621523292
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_465
timestamp 1621523292
transform 1 0 43884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1621523292
transform 1 0 44988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1621523292
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1621523292
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1621523292
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_486
timestamp 1621523292
transform 1 0 45816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_498
timestamp 1621523292
transform 1 0 46920 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1621523292
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1621523292
transform 1 0 49220 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1621523292
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_514
timestamp 1621523292
transform 1 0 48392 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_522
timestamp 1621523292
transform 1 0 49128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_510
timestamp 1621523292
transform 1 0 48024 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_522
timestamp 1621523292
transform 1 0 49128 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_526
timestamp 1621523292
transform 1 0 49496 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0953_
timestamp 1621523292
transform 1 0 49864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_538
timestamp 1621523292
transform 1 0 50600 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_534
timestamp 1621523292
transform 1 0 50232 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_540
timestamp 1621523292
transform 1 0 50784 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_533
timestamp 1621523292
transform 1 0 50140 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1179_
timestamp 1621523292
transform 1 0 50324 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0952_
timestamp 1621523292
transform 1 0 50508 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_543
timestamp 1621523292
transform 1 0 51060 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1621523292
transform 1 0 50968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1621523292
transform 1 0 51152 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_551
timestamp 1621523292
transform 1 0 51796 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_554
timestamp 1621523292
transform 1 0 52072 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_547
timestamp 1621523292
transform 1 0 51428 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0906_
timestamp 1621523292
transform 1 0 51796 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1621523292
transform 1 0 51888 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_555
timestamp 1621523292
transform 1 0 52164 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_561
timestamp 1621523292
transform 1 0 52716 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0832_
timestamp 1621523292
transform 1 0 52440 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0831_
timestamp 1621523292
transform 1 0 52532 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_40_566
timestamp 1621523292
transform 1 0 53176 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_573
timestamp 1621523292
transform 1 0 53820 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_571
timestamp 1621523292
transform 1 0 53636 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_569
timestamp 1621523292
transform 1 0 53452 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1621523292
transform 1 0 53544 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0830_
timestamp 1621523292
transform 1 0 54004 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0695_
timestamp 1621523292
transform 1 0 53544 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_584
timestamp 1621523292
transform 1 0 54832 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_581
timestamp 1621523292
transform 1 0 54556 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0696_
timestamp 1621523292
transform 1 0 54188 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0621_
timestamp 1621523292
transform 1 0 54924 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_588
timestamp 1621523292
transform 1 0 55200 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1621523292
transform 1 0 55200 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_591
timestamp 1621523292
transform 1 0 55476 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1621523292
transform 1 0 55936 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_604
timestamp 1621523292
transform 1 0 56672 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_600
timestamp 1621523292
transform 1 0 56304 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_607
timestamp 1621523292
transform 1 0 56948 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_599
timestamp 1621523292
transform 1 0 56212 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output220
timestamp 1621523292
transform 1 0 56764 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1621523292
transform 1 0 56212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_609
timestamp 1621523292
transform 1 0 57132 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output219
timestamp 1621523292
transform 1 0 57132 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1323_
timestamp 1621523292
transform 1 0 57500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1621523292
transform -1 0 58880 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1621523292
transform -1 0 58880 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output181
timestamp 1621523292
transform 1 0 57868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_613
timestamp 1621523292
transform 1 0 57500 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1621523292
transform 1 0 58236 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1621523292
transform 1 0 58236 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1621523292
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output305
timestamp 1621523292
transform 1 0 1748 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output306
timestamp 1621523292
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1621523292
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_11
timestamp 1621523292
transform 1 0 2116 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_19
timestamp 1621523292
transform 1 0 2852 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1016_
timestamp 1621523292
transform 1 0 3220 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_26
timestamp 1621523292
transform 1 0 3496 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1621523292
transform 1 0 4600 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1621523292
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1621523292
transform 1 0 5704 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_56
timestamp 1621523292
transform 1 0 6256 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1621523292
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1621523292
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1621523292
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1621523292
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1621523292
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1621523292
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1621523292
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1621523292
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1621523292
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1621523292
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1621523292
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1621523292
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1621523292
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1621523292
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1621523292
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1621523292
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1621523292
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1621523292
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1621523292
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_241
timestamp 1621523292
transform 1 0 23276 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_253
timestamp 1621523292
transform 1 0 24380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_265
timestamp 1621523292
transform 1 0 25484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_277
timestamp 1621523292
transform 1 0 26588 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1621523292
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1621523292
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_298
timestamp 1621523292
transform 1 0 28520 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_310
timestamp 1621523292
transform 1 0 29624 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_322
timestamp 1621523292
transform 1 0 30728 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1621523292
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_334
timestamp 1621523292
transform 1 0 31832 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1621523292
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_355
timestamp 1621523292
transform 1 0 33764 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1621523292
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1621523292
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_391
timestamp 1621523292
transform 1 0 37076 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1621523292
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_400
timestamp 1621523292
transform 1 0 37904 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_412
timestamp 1621523292
transform 1 0 39008 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_424
timestamp 1621523292
transform 1 0 40112 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_436
timestamp 1621523292
transform 1 0 41216 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1621523292
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_448
timestamp 1621523292
transform 1 0 42320 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_457
timestamp 1621523292
transform 1 0 43148 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_469
timestamp 1621523292
transform 1 0 44252 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_481
timestamp 1621523292
transform 1 0 45356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_493
timestamp 1621523292
transform 1 0 46460 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1621523292
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1621523292
transform 1 0 47564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_514
timestamp 1621523292
transform 1 0 48392 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0612_
timestamp 1621523292
transform 1 0 50784 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0945_
timestamp 1621523292
transform 1 0 50140 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1621523292
transform 1 0 49496 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_529
timestamp 1621523292
transform 1 0 49772 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_536
timestamp 1621523292
transform 1 0 50416 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_544
timestamp 1621523292
transform 1 0 51152 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1621523292
transform 1 0 51704 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_566
timestamp 1621523292
transform 1 0 53176 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1621523292
transform 1 0 54004 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1621523292
transform 1 0 54924 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1621523292
transform 1 0 53544 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_571
timestamp 1621523292
transform 1 0 53636 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_578
timestamp 1621523292
transform 1 0 54280 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_584
timestamp 1621523292
transform 1 0 54832 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0901_
timestamp 1621523292
transform 1 0 57224 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_601
timestamp 1621523292
transform 1 0 56396 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_609
timestamp 1621523292
transform 1 0 57132 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1621523292
transform -1 0 58880 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output182
timestamp 1621523292
transform 1 0 57868 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_613
timestamp 1621523292
transform 1 0 57500 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_621
timestamp 1621523292
transform 1 0 58236 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1621523292
transform 1 0 2944 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1233_
timestamp 1621523292
transform 1 0 1840 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1621523292
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1621523292
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_7
timestamp 1621523292
transform 1 0 1748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_16
timestamp 1621523292
transform 1 0 2576 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1621523292
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_23
timestamp 1621523292
transform 1 0 3220 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1621523292
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1621523292
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1621523292
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1621523292
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1621523292
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1621523292
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_87
timestamp 1621523292
transform 1 0 9108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_99
timestamp 1621523292
transform 1 0 10212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_111
timestamp 1621523292
transform 1 0 11316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_123
timestamp 1621523292
transform 1 0 12420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1621523292
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_135
timestamp 1621523292
transform 1 0 13524 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1621523292
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1621523292
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1621523292
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1621523292
transform 1 0 17664 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_192
timestamp 1621523292
transform 1 0 18768 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1621523292
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1621523292
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1621523292
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1621523292
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1621523292
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1621523292
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1621523292
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1621523292
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1621523292
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1621523292
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1621523292
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1621523292
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1621523292
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1621523292
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1621523292
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1621523292
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1621523292
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1621523292
transform 1 0 33396 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_363
timestamp 1621523292
transform 1 0 34500 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_372
timestamp 1621523292
transform 1 0 35328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_384
timestamp 1621523292
transform 1 0 36432 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_396
timestamp 1621523292
transform 1 0 37536 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_408
timestamp 1621523292
transform 1 0 38640 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1621523292
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_420
timestamp 1621523292
transform 1 0 39744 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_429
timestamp 1621523292
transform 1 0 40572 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_441
timestamp 1621523292
transform 1 0 41676 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_453
timestamp 1621523292
transform 1 0 42780 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_465
timestamp 1621523292
transform 1 0 43884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1621523292
transform 1 0 44988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1621523292
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_486
timestamp 1621523292
transform 1 0 45816 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_498
timestamp 1621523292
transform 1 0 46920 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1621523292
transform 1 0 48024 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_522
timestamp 1621523292
transform 1 0 49128 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1075_
timestamp 1621523292
transform 1 0 50324 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1180_
timestamp 1621523292
transform 1 0 49680 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1621523292
transform 1 0 50968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_531
timestamp 1621523292
transform 1 0 49956 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_538
timestamp 1621523292
transform 1 0 50600 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_543
timestamp 1621523292
transform 1 0 51060 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0903_
timestamp 1621523292
transform 1 0 52164 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0905_
timestamp 1621523292
transform 1 0 51520 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52808 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_42_547
timestamp 1621523292
transform 1 0 51428 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_551
timestamp 1621523292
transform 1 0 51796 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_558
timestamp 1621523292
transform 1 0 52440 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0617_
timestamp 1621523292
transform 1 0 55016 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_582
timestamp 1621523292
transform 1 0 54648 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_589
timestamp 1621523292
transform 1 0 55292 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1286_
timestamp 1621523292
transform 1 0 56764 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1621523292
transform 1 0 56212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_597
timestamp 1621523292
transform 1 0 56028 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_600
timestamp 1621523292
transform 1 0 56304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_604
timestamp 1621523292
transform 1 0 56672 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1621523292
transform -1 0 58880 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output221
timestamp 1621523292
transform 1 0 57868 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1621523292
transform 1 0 57500 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1621523292
transform 1 0 58236 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1014_
timestamp 1621523292
transform 1 0 2484 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1621523292
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output307
timestamp 1621523292
transform 1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1621523292
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_11
timestamp 1621523292
transform 1 0 2116 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_18
timestamp 1621523292
transform 1 0 2760 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1120_
timestamp 1621523292
transform 1 0 3128 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_25
timestamp 1621523292
transform 1 0 3404 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_37
timestamp 1621523292
transform 1 0 4508 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1621523292
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_49
timestamp 1621523292
transform 1 0 5612 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1621523292
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1621523292
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1621523292
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1621523292
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1621523292
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1621523292
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_115
timestamp 1621523292
transform 1 0 11684 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1621523292
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_139
timestamp 1621523292
transform 1 0 13892 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_151
timestamp 1621523292
transform 1 0 14996 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1621523292
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_163
timestamp 1621523292
transform 1 0 16100 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_172
timestamp 1621523292
transform 1 0 16928 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1621523292
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1621523292
transform 1 0 19136 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1621523292
transform 1 0 20240 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1621523292
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1621523292
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1621523292
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1621523292
transform 1 0 23276 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_253
timestamp 1621523292
transform 1 0 24380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_265
timestamp 1621523292
transform 1 0 25484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_277
timestamp 1621523292
transform 1 0 26588 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1621523292
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1621523292
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_298
timestamp 1621523292
transform 1 0 28520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_310
timestamp 1621523292
transform 1 0 29624 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_322
timestamp 1621523292
transform 1 0 30728 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1621523292
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_334
timestamp 1621523292
transform 1 0 31832 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_343
timestamp 1621523292
transform 1 0 32660 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_355
timestamp 1621523292
transform 1 0 33764 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1621523292
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1621523292
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_391
timestamp 1621523292
transform 1 0 37076 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1621523292
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_400
timestamp 1621523292
transform 1 0 37904 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_412
timestamp 1621523292
transform 1 0 39008 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_424
timestamp 1621523292
transform 1 0 40112 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_436
timestamp 1621523292
transform 1 0 41216 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1621523292
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_448
timestamp 1621523292
transform 1 0 42320 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1621523292
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1621523292
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_481
timestamp 1621523292
transform 1 0 45356 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_493
timestamp 1621523292
transform 1 0 46460 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1621523292
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1621523292
transform 1 0 49312 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1621523292
transform 1 0 47564 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_514
timestamp 1621523292
transform 1 0 48392 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_522
timestamp 1621523292
transform 1 0 49128 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _0615_
timestamp 1621523292
transform 1 0 49956 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1621523292
transform 1 0 50600 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_527
timestamp 1621523292
transform 1 0 49588 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_534
timestamp 1621523292
transform 1 0 50232 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1621523292
transform 1 0 52440 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_554
timestamp 1621523292
transform 1 0 52072 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_561
timestamp 1621523292
transform 1 0 52716 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0616_
timestamp 1621523292
transform 1 0 54280 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1621523292
transform 1 0 54924 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1621523292
transform 1 0 53544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_569
timestamp 1621523292
transform 1 0 53452 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_571
timestamp 1621523292
transform 1 0 53636 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_577
timestamp 1621523292
transform 1 0 54188 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_581
timestamp 1621523292
transform 1 0 54556 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0682_
timestamp 1621523292
transform 1 0 56764 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_601
timestamp 1621523292
transform 1 0 56396 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_608
timestamp 1621523292
transform 1 0 57040 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1324_
timestamp 1621523292
transform 1 0 57500 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1621523292
transform -1 0 58880 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_612
timestamp 1621523292
transform 1 0 57408 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_621
timestamp 1621523292
transform 1 0 58236 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1121_
timestamp 1621523292
transform 1 0 2760 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1234_
timestamp 1621523292
transform 1 0 1656 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1621523292
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1621523292
transform 1 0 1380 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_14
timestamp 1621523292
transform 1 0 2392 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_21
timestamp 1621523292
transform 1 0 3036 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1621523292
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_30
timestamp 1621523292
transform 1 0 3864 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_42
timestamp 1621523292
transform 1 0 4968 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_54
timestamp 1621523292
transform 1 0 6072 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1621523292
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_66
timestamp 1621523292
transform 1 0 7176 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_78
timestamp 1621523292
transform 1 0 8280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_87
timestamp 1621523292
transform 1 0 9108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_99
timestamp 1621523292
transform 1 0 10212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_111
timestamp 1621523292
transform 1 0 11316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_123
timestamp 1621523292
transform 1 0 12420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1621523292
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_135
timestamp 1621523292
transform 1 0 13524 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_144
timestamp 1621523292
transform 1 0 14352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_156
timestamp 1621523292
transform 1 0 15456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_168
timestamp 1621523292
transform 1 0 16560 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_180
timestamp 1621523292
transform 1 0 17664 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_192
timestamp 1621523292
transform 1 0 18768 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1621523292
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_201
timestamp 1621523292
transform 1 0 19596 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_213
timestamp 1621523292
transform 1 0 20700 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_225
timestamp 1621523292
transform 1 0 21804 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_237
timestamp 1621523292
transform 1 0 22908 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1621523292
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_249
timestamp 1621523292
transform 1 0 24012 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_258
timestamp 1621523292
transform 1 0 24840 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_270
timestamp 1621523292
transform 1 0 25944 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_282
timestamp 1621523292
transform 1 0 27048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1621523292
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1621523292
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_306
timestamp 1621523292
transform 1 0 29256 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_315
timestamp 1621523292
transform 1 0 30084 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_327
timestamp 1621523292
transform 1 0 31188 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_339
timestamp 1621523292
transform 1 0 32292 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1621523292
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_351
timestamp 1621523292
transform 1 0 33396 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_363
timestamp 1621523292
transform 1 0 34500 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_372
timestamp 1621523292
transform 1 0 35328 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_384
timestamp 1621523292
transform 1 0 36432 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_396
timestamp 1621523292
transform 1 0 37536 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_408
timestamp 1621523292
transform 1 0 38640 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1621523292
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_420
timestamp 1621523292
transform 1 0 39744 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_429
timestamp 1621523292
transform 1 0 40572 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_441
timestamp 1621523292
transform 1 0 41676 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_453
timestamp 1621523292
transform 1 0 42780 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_465
timestamp 1621523292
transform 1 0 43884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_477
timestamp 1621523292
transform 1 0 44988 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1621523292
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1621523292
transform 1 0 45816 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_498
timestamp 1621523292
transform 1 0 46920 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1181_
timestamp 1621523292
transform 1 0 49036 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_510
timestamp 1621523292
transform 1 0 48024 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_518
timestamp 1621523292
transform 1 0 48760 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_524
timestamp 1621523292
transform 1 0 49312 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0614_
timestamp 1621523292
transform 1 0 50324 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0950_
timestamp 1621523292
transform 1 0 49680 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1621523292
transform 1 0 50968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_531
timestamp 1621523292
transform 1 0 49956 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_538
timestamp 1621523292
transform 1 0 50600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_543
timestamp 1621523292
transform 1 0 51060 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0677_
timestamp 1621523292
transform 1 0 51428 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1621523292
transform 1 0 52900 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_44_554
timestamp 1621523292
transform 1 0 52072 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_562
timestamp 1621523292
transform 1 0 52808 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0683_
timestamp 1621523292
transform 1 0 54740 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_44_579
timestamp 1621523292
transform 1 0 54372 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1621523292
transform 1 0 56212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output222
timestamp 1621523292
transform 1 0 57132 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_590
timestamp 1621523292
transform 1 0 55384 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_598
timestamp 1621523292
transform 1 0 56120 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_600
timestamp 1621523292
transform 1 0 56304 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_608
timestamp 1621523292
transform 1 0 57040 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1621523292
transform -1 0 58880 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output183
timestamp 1621523292
transform 1 0 57868 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_613
timestamp 1621523292
transform 1 0 57500 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_621
timestamp 1621523292
transform 1 0 58236 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1621523292
transform 1 0 2484 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1621523292
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output308
timestamp 1621523292
transform 1 0 1748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1621523292
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_11
timestamp 1621523292
transform 1 0 2116 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1621523292
transform 1 0 2760 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1122_
timestamp 1621523292
transform 1 0 3128 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_25
timestamp 1621523292
transform 1 0 3404 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_37
timestamp 1621523292
transform 1 0 4508 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1621523292
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_49
timestamp 1621523292
transform 1 0 5612 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_58
timestamp 1621523292
transform 1 0 6440 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_70
timestamp 1621523292
transform 1 0 7544 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_82
timestamp 1621523292
transform 1 0 8648 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_94
timestamp 1621523292
transform 1 0 9752 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_106
timestamp 1621523292
transform 1 0 10856 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1621523292
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_115
timestamp 1621523292
transform 1 0 11684 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_127
timestamp 1621523292
transform 1 0 12788 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1621523292
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1621523292
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1621523292
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_163
timestamp 1621523292
transform 1 0 16100 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_172
timestamp 1621523292
transform 1 0 16928 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1621523292
transform 1 0 18032 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1621523292
transform 1 0 19136 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1621523292
transform 1 0 20240 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1621523292
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1621523292
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_229
timestamp 1621523292
transform 1 0 22172 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1621523292
transform 1 0 23276 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_253
timestamp 1621523292
transform 1 0 24380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_265
timestamp 1621523292
transform 1 0 25484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_277
timestamp 1621523292
transform 1 0 26588 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1621523292
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_286
timestamp 1621523292
transform 1 0 27416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_298
timestamp 1621523292
transform 1 0 28520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_310
timestamp 1621523292
transform 1 0 29624 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_322
timestamp 1621523292
transform 1 0 30728 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1621523292
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_334
timestamp 1621523292
transform 1 0 31832 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_343
timestamp 1621523292
transform 1 0 32660 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_355
timestamp 1621523292
transform 1 0 33764 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1621523292
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1621523292
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_391
timestamp 1621523292
transform 1 0 37076 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1621523292
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1621523292
transform 1 0 37904 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_412
timestamp 1621523292
transform 1 0 39008 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_424
timestamp 1621523292
transform 1 0 40112 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_436
timestamp 1621523292
transform 1 0 41216 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1621523292
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_448
timestamp 1621523292
transform 1 0 42320 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_457
timestamp 1621523292
transform 1 0 43148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_469
timestamp 1621523292
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1621523292
transform 1 0 45356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_493
timestamp 1621523292
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1621523292
transform 1 0 49220 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1621523292
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1621523292
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_514
timestamp 1621523292
transform 1 0 48392 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_522
timestamp 1621523292
transform 1 0 49128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _0820_
timestamp 1621523292
transform 1 0 51060 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_539
timestamp 1621523292
transform 1 0 50692 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _0823_
timestamp 1621523292
transform 1 0 52532 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_45_551
timestamp 1621523292
transform 1 0 51796 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_566
timestamp 1621523292
transform 1 0 53176 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0756_
timestamp 1621523292
transform 1 0 54740 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1621523292
transform 1 0 54004 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1621523292
transform 1 0 53544 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_571
timestamp 1621523292
transform 1 0 53636 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_578
timestamp 1621523292
transform 1 0 54280 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_582
timestamp 1621523292
transform 1 0 54648 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0679_
timestamp 1621523292
transform 1 0 56120 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1287_
timestamp 1621523292
transform 1 0 57132 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_590
timestamp 1621523292
transform 1 0 55384 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_601
timestamp 1621523292
transform 1 0 56396 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1621523292
transform -1 0 58880 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_617
timestamp 1621523292
transform 1 0 57868 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1621523292
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1621523292
transform 1 0 1380 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output309
timestamp 1621523292
transform 1 0 1748 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1621523292
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1621523292
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1235_
timestamp 1621523292
transform 1 0 1656 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_18
timestamp 1621523292
transform 1 0 2760 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_11
timestamp 1621523292
transform 1 0 2116 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1621523292
transform 1 0 2484 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_14
timestamp 1621523292
transform 1 0 2392 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1011_
timestamp 1621523292
transform 1 0 3128 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1123_
timestamp 1621523292
transform 1 0 3772 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1621523292
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_26
timestamp 1621523292
transform 1 0 3496 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_30
timestamp 1621523292
transform 1 0 3864 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_42
timestamp 1621523292
transform 1 0 4968 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_25
timestamp 1621523292
transform 1 0 3404 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_32
timestamp 1621523292
transform 1 0 4048 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1621523292
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_54
timestamp 1621523292
transform 1 0 6072 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_44
timestamp 1621523292
transform 1 0 5152 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_56
timestamp 1621523292
transform 1 0 6256 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_58
timestamp 1621523292
transform 1 0 6440 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1621523292
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_66
timestamp 1621523292
transform 1 0 7176 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_78
timestamp 1621523292
transform 1 0 8280 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1621523292
transform 1 0 9108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_70
timestamp 1621523292
transform 1 0 7544 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_82
timestamp 1621523292
transform 1 0 8648 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_99
timestamp 1621523292
transform 1 0 10212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_94
timestamp 1621523292
transform 1 0 9752 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_106
timestamp 1621523292
transform 1 0 10856 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1621523292
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_111
timestamp 1621523292
transform 1 0 11316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_123
timestamp 1621523292
transform 1 0 12420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_115
timestamp 1621523292
transform 1 0 11684 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_127
timestamp 1621523292
transform 1 0 12788 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1621523292
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_135
timestamp 1621523292
transform 1 0 13524 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_144
timestamp 1621523292
transform 1 0 14352 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_139
timestamp 1621523292
transform 1 0 13892 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_151
timestamp 1621523292
transform 1 0 14996 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1621523292
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_156
timestamp 1621523292
transform 1 0 15456 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_168
timestamp 1621523292
transform 1 0 16560 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_163
timestamp 1621523292
transform 1 0 16100 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_172
timestamp 1621523292
transform 1 0 16928 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1621523292
transform 1 0 17664 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_192
timestamp 1621523292
transform 1 0 18768 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1621523292
transform 1 0 18032 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1621523292
transform 1 0 19136 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1621523292
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_201
timestamp 1621523292
transform 1 0 19596 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_213
timestamp 1621523292
transform 1 0 20700 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1621523292
transform 1 0 20240 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1621523292
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1621523292
transform 1 0 21804 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1621523292
transform 1 0 22908 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1621523292
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1621523292
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1621523292
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_249
timestamp 1621523292
transform 1 0 24012 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_258
timestamp 1621523292
transform 1 0 24840 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_241
timestamp 1621523292
transform 1 0 23276 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_253
timestamp 1621523292
transform 1 0 24380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_270
timestamp 1621523292
transform 1 0 25944 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_282
timestamp 1621523292
transform 1 0 27048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_265
timestamp 1621523292
transform 1 0 25484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1621523292
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1621523292
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_294
timestamp 1621523292
transform 1 0 28152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_286
timestamp 1621523292
transform 1 0 27416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_298
timestamp 1621523292
transform 1 0 28520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1621523292
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1621523292
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_315
timestamp 1621523292
transform 1 0 30084 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_327
timestamp 1621523292
transform 1 0 31188 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_310
timestamp 1621523292
transform 1 0 29624 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_322
timestamp 1621523292
transform 1 0 30728 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1621523292
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_339
timestamp 1621523292
transform 1 0 32292 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_334
timestamp 1621523292
transform 1 0 31832 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_343
timestamp 1621523292
transform 1 0 32660 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1621523292
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_351
timestamp 1621523292
transform 1 0 33396 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_363
timestamp 1621523292
transform 1 0 34500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_355
timestamp 1621523292
transform 1 0 33764 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1621523292
transform 1 0 34868 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_372
timestamp 1621523292
transform 1 0 35328 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_384
timestamp 1621523292
transform 1 0 36432 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1621523292
transform 1 0 35972 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_391
timestamp 1621523292
transform 1 0 37076 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1621523292
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1621523292
transform 1 0 37536 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1621523292
transform 1 0 38640 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_400
timestamp 1621523292
transform 1 0 37904 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_412
timestamp 1621523292
transform 1 0 39008 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1621523292
transform 1 0 40480 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_420
timestamp 1621523292
transform 1 0 39744 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_429
timestamp 1621523292
transform 1 0 40572 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_424
timestamp 1621523292
transform 1 0 40112 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_436
timestamp 1621523292
transform 1 0 41216 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1621523292
transform 1 0 43056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_441
timestamp 1621523292
transform 1 0 41676 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_453
timestamp 1621523292
transform 1 0 42780 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_448
timestamp 1621523292
transform 1 0 42320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_457
timestamp 1621523292
transform 1 0 43148 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_465
timestamp 1621523292
transform 1 0 43884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1621523292
transform 1 0 44988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_469
timestamp 1621523292
transform 1 0 44252 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1621523292
transform 1 0 45724 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_486
timestamp 1621523292
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_498
timestamp 1621523292
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_481
timestamp 1621523292
transform 1 0 45356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_493
timestamp 1621523292
transform 1 0 46460 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1074_
timestamp 1621523292
transform 1 0 49036 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1621523292
transform 1 0 48760 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1621523292
transform 1 0 48300 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1621523292
transform 1 0 48392 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_510
timestamp 1621523292
transform 1 0 48024 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_517
timestamp 1621523292
transform 1 0 48668 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_524
timestamp 1621523292
transform 1 0 49312 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1621523292
transform 1 0 47564 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_514
timestamp 1621523292
transform 1 0 48392 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0613_
timestamp 1621523292
transform 1 0 50600 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1621523292
transform 1 0 50324 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0949_
timestamp 1621523292
transform 1 0 49680 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1621523292
transform 1 0 50968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_531
timestamp 1621523292
transform 1 0 49956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_538
timestamp 1621523292
transform 1 0 50600 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_543
timestamp 1621523292
transform 1 0 51060 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_534
timestamp 1621523292
transform 1 0 50232 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_541
timestamp 1621523292
transform 1 0 50876 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0815_
timestamp 1621523292
transform 1 0 52348 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0817_
timestamp 1621523292
transform 1 0 51428 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1621523292
transform 1 0 51612 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0825_
timestamp 1621523292
transform 1 0 52440 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_553
timestamp 1621523292
transform 1 0 51980 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_564
timestamp 1621523292
transform 1 0 52992 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_554
timestamp 1621523292
transform 1 0 52072 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_566
timestamp 1621523292
transform 1 0 53176 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_571
timestamp 1621523292
transform 1 0 53636 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_575
timestamp 1621523292
transform 1 0 54004 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_571
timestamp 1621523292
transform 1 0 53636 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1621523292
transform 1 0 53544 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0822_
timestamp 1621523292
transform 1 0 54004 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0681_
timestamp 1621523292
transform 1 0 53360 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0680_
timestamp 1621523292
transform 1 0 54096 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_47_581
timestamp 1621523292
transform 1 0 54556 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_583
timestamp 1621523292
transform 1 0 54740 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0757_
timestamp 1621523292
transform 1 0 55108 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1621523292
transform 1 0 55108 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_46_598
timestamp 1621523292
transform 1 0 56120 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_594
timestamp 1621523292
transform 1 0 55752 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_607
timestamp 1621523292
transform 1 0 56948 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_603
timestamp 1621523292
transform 1 0 56580 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_604
timestamp 1621523292
transform 1 0 56672 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_600
timestamp 1621523292
transform 1 0 56304 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output184
timestamp 1621523292
transform 1 0 56764 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1621523292
transform 1 0 56212 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_609
timestamp 1621523292
transform 1 0 57132 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1288_
timestamp 1621523292
transform 1 0 57040 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1325_
timestamp 1621523292
transform 1 0 57500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1621523292
transform -1 0 58880 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1621523292
transform -1 0 58880 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1621523292
transform 1 0 58236 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_616
timestamp 1621523292
transform 1 0 57776 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_624
timestamp 1621523292
transform 1 0 58512 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1236_
timestamp 1621523292
transform 1 0 1748 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1621523292
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1621523292
transform 1 0 1380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1621523292
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1621523292
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1621523292
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_30
timestamp 1621523292
transform 1 0 3864 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_42
timestamp 1621523292
transform 1 0 4968 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_54
timestamp 1621523292
transform 1 0 6072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1621523292
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_66
timestamp 1621523292
transform 1 0 7176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1621523292
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_87
timestamp 1621523292
transform 1 0 9108 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_99
timestamp 1621523292
transform 1 0 10212 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_111
timestamp 1621523292
transform 1 0 11316 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_123
timestamp 1621523292
transform 1 0 12420 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1621523292
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_135
timestamp 1621523292
transform 1 0 13524 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_144
timestamp 1621523292
transform 1 0 14352 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_156
timestamp 1621523292
transform 1 0 15456 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_168
timestamp 1621523292
transform 1 0 16560 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_180
timestamp 1621523292
transform 1 0 17664 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_192
timestamp 1621523292
transform 1 0 18768 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1621523292
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_201
timestamp 1621523292
transform 1 0 19596 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_213
timestamp 1621523292
transform 1 0 20700 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1621523292
transform 1 0 21804 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1621523292
transform 1 0 22908 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1621523292
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_249
timestamp 1621523292
transform 1 0 24012 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_258
timestamp 1621523292
transform 1 0 24840 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_270
timestamp 1621523292
transform 1 0 25944 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_282
timestamp 1621523292
transform 1 0 27048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_294
timestamp 1621523292
transform 1 0 28152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1621523292
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1621523292
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1621523292
transform 1 0 30084 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_327
timestamp 1621523292
transform 1 0 31188 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_339
timestamp 1621523292
transform 1 0 32292 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1621523292
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_351
timestamp 1621523292
transform 1 0 33396 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_363
timestamp 1621523292
transform 1 0 34500 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1621523292
transform 1 0 35328 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1621523292
transform 1 0 36432 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_396
timestamp 1621523292
transform 1 0 37536 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_408
timestamp 1621523292
transform 1 0 38640 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1621523292
transform 1 0 40480 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_420
timestamp 1621523292
transform 1 0 39744 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_429
timestamp 1621523292
transform 1 0 40572 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_441
timestamp 1621523292
transform 1 0 41676 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_453
timestamp 1621523292
transform 1 0 42780 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_465
timestamp 1621523292
transform 1 0 43884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1621523292
transform 1 0 44988 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1621523292
transform 1 0 45724 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1621523292
transform 1 0 47104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_486
timestamp 1621523292
transform 1 0 45816 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_498
timestamp 1621523292
transform 1 0 46920 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _1076_
timestamp 1621523292
transform 1 0 49036 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1621523292
transform 1 0 48392 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 47748 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_503
timestamp 1621523292
transform 1 0 47380 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_510
timestamp 1621523292
transform 1 0 48024 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_517
timestamp 1621523292
transform 1 0 48668 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_524
timestamp 1621523292
transform 1 0 49312 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0674_
timestamp 1621523292
transform 1 0 50324 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0678_
timestamp 1621523292
transform 1 0 49680 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1621523292
transform 1 0 50968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_531
timestamp 1621523292
transform 1 0 49956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_538
timestamp 1621523292
transform 1 0 50600 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_543
timestamp 1621523292
transform 1 0 51060 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0759_
timestamp 1621523292
transform 1 0 51704 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1621523292
transform 1 0 53268 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_549
timestamp 1621523292
transform 1 0 51612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_559
timestamp 1621523292
transform 1 0 52532 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1621523292
transform 1 0 55108 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_583
timestamp 1621523292
transform 1 0 54740 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1621523292
transform 1 0 56212 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output223
timestamp 1621523292
transform 1 0 56764 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_590
timestamp 1621523292
transform 1 0 55384 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_598
timestamp 1621523292
transform 1 0 56120 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_600
timestamp 1621523292
transform 1 0 56304 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_604
timestamp 1621523292
transform 1 0 56672 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_609
timestamp 1621523292
transform 1 0 57132 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1326_
timestamp 1621523292
transform 1 0 57500 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1621523292
transform -1 0 58880 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_621
timestamp 1621523292
transform 1 0 58236 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1237_
timestamp 1621523292
transform 1 0 1564 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1621523292
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1621523292
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_13
timestamp 1621523292
transform 1 0 2300 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_25
timestamp 1621523292
transform 1 0 3404 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_37
timestamp 1621523292
transform 1 0 4508 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1621523292
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_49
timestamp 1621523292
transform 1 0 5612 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_58
timestamp 1621523292
transform 1 0 6440 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_70
timestamp 1621523292
transform 1 0 7544 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_82
timestamp 1621523292
transform 1 0 8648 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_94
timestamp 1621523292
transform 1 0 9752 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1621523292
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1621523292
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_115
timestamp 1621523292
transform 1 0 11684 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_127
timestamp 1621523292
transform 1 0 12788 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_139
timestamp 1621523292
transform 1 0 13892 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_151
timestamp 1621523292
transform 1 0 14996 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1621523292
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_163
timestamp 1621523292
transform 1 0 16100 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_172
timestamp 1621523292
transform 1 0 16928 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1621523292
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1621523292
transform 1 0 19136 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1621523292
transform 1 0 20240 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1621523292
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_220
timestamp 1621523292
transform 1 0 21344 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_229
timestamp 1621523292
transform 1 0 22172 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_241
timestamp 1621523292
transform 1 0 23276 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_253
timestamp 1621523292
transform 1 0 24380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_265
timestamp 1621523292
transform 1 0 25484 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_277
timestamp 1621523292
transform 1 0 26588 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1621523292
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_286
timestamp 1621523292
transform 1 0 27416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_298
timestamp 1621523292
transform 1 0 28520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1621523292
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1621523292
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1621523292
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_334
timestamp 1621523292
transform 1 0 31832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_343
timestamp 1621523292
transform 1 0 32660 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1621523292
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1621523292
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1621523292
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_391
timestamp 1621523292
transform 1 0 37076 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1621523292
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_400
timestamp 1621523292
transform 1 0 37904 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_412
timestamp 1621523292
transform 1 0 39008 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_424
timestamp 1621523292
transform 1 0 40112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_436
timestamp 1621523292
transform 1 0 41216 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1621523292
transform 1 0 43056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_448
timestamp 1621523292
transform 1 0 42320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_457
timestamp 1621523292
transform 1 0 43148 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_469
timestamp 1621523292
transform 1 0 44252 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_481
timestamp 1621523292
transform 1 0 45356 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_493
timestamp 1621523292
transform 1 0 46460 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1182_
timestamp 1621523292
transform 1 0 48760 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1621523292
transform 1 0 48300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1621523292
transform 1 0 47656 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_505
timestamp 1621523292
transform 1 0 47564 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_509
timestamp 1621523292
transform 1 0 47932 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_514
timestamp 1621523292
transform 1 0 48392 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_521
timestamp 1621523292
transform 1 0 49036 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0675_
timestamp 1621523292
transform 1 0 50048 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0758_
timestamp 1621523292
transform 1 0 51244 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1077_
timestamp 1621523292
transform 1 0 49404 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_528
timestamp 1621523292
transform 1 0 49680 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_539
timestamp 1621523292
transform 1 0 50692 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _0684_
timestamp 1621523292
transform 1 0 52256 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_49_552
timestamp 1621523292
transform 1 0 51888 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_565
timestamp 1621523292
transform 1 0 53084 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0619_
timestamp 1621523292
transform 1 0 54924 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0812_
timestamp 1621523292
transform 1 0 54004 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1621523292
transform 1 0 53544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_569
timestamp 1621523292
transform 1 0 53452 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_571
timestamp 1621523292
transform 1 0 53636 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_578
timestamp 1621523292
transform 1 0 54280 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_584
timestamp 1621523292
transform 1 0 54832 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_588
timestamp 1621523292
transform 1 0 55200 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0688_
timestamp 1621523292
transform 1 0 56396 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0899_
timestamp 1621523292
transform 1 0 57224 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0902_
timestamp 1621523292
transform 1 0 55752 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_597
timestamp 1621523292
transform 1 0 56028 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_604
timestamp 1621523292
transform 1 0 56672 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1621523292
transform -1 0 58880 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output185
timestamp 1621523292
transform 1 0 57868 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_613
timestamp 1621523292
transform 1 0 57500 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_621
timestamp 1621523292
transform 1 0 58236 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1124_
timestamp 1621523292
transform 1 0 2484 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1621523292
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output311
timestamp 1621523292
transform 1 0 1748 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1621523292
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_11
timestamp 1621523292
transform 1 0 2116 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_18
timestamp 1621523292
transform 1 0 2760 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1621523292
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_26
timestamp 1621523292
transform 1 0 3496 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1621523292
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1621523292
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_54
timestamp 1621523292
transform 1 0 6072 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1621523292
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_66
timestamp 1621523292
transform 1 0 7176 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_78
timestamp 1621523292
transform 1 0 8280 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_87
timestamp 1621523292
transform 1 0 9108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_99
timestamp 1621523292
transform 1 0 10212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_111
timestamp 1621523292
transform 1 0 11316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1621523292
transform 1 0 12420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1621523292
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_135
timestamp 1621523292
transform 1 0 13524 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_144
timestamp 1621523292
transform 1 0 14352 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_156
timestamp 1621523292
transform 1 0 15456 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_168
timestamp 1621523292
transform 1 0 16560 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_180
timestamp 1621523292
transform 1 0 17664 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_192
timestamp 1621523292
transform 1 0 18768 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1621523292
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_201
timestamp 1621523292
transform 1 0 19596 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_213
timestamp 1621523292
transform 1 0 20700 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_225
timestamp 1621523292
transform 1 0 21804 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_237
timestamp 1621523292
transform 1 0 22908 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1621523292
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_249
timestamp 1621523292
transform 1 0 24012 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_258
timestamp 1621523292
transform 1 0 24840 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_270
timestamp 1621523292
transform 1 0 25944 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_282
timestamp 1621523292
transform 1 0 27048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_294
timestamp 1621523292
transform 1 0 28152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1621523292
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_306
timestamp 1621523292
transform 1 0 29256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1621523292
transform 1 0 30084 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_327
timestamp 1621523292
transform 1 0 31188 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_339
timestamp 1621523292
transform 1 0 32292 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1621523292
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_351
timestamp 1621523292
transform 1 0 33396 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_363
timestamp 1621523292
transform 1 0 34500 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_372
timestamp 1621523292
transform 1 0 35328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1621523292
transform 1 0 36432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_396
timestamp 1621523292
transform 1 0 37536 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_408
timestamp 1621523292
transform 1 0 38640 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1621523292
transform 1 0 40480 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_420
timestamp 1621523292
transform 1 0 39744 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_429
timestamp 1621523292
transform 1 0 40572 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_441
timestamp 1621523292
transform 1 0 41676 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_453
timestamp 1621523292
transform 1 0 42780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_465
timestamp 1621523292
transform 1 0 43884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1621523292
transform 1 0 44988 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1621523292
transform 1 0 45724 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_486
timestamp 1621523292
transform 1 0 45816 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_498
timestamp 1621523292
transform 1 0 46920 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _0819_
timestamp 1621523292
transform 1 0 49312 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0948_
timestamp 1621523292
transform 1 0 48668 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_510
timestamp 1621523292
transform 1 0 48024 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_516
timestamp 1621523292
transform 1 0 48576 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_520
timestamp 1621523292
transform 1 0 48944 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _0818_
timestamp 1621523292
transform 1 0 49956 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1621523292
transform 1 0 50968 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_527
timestamp 1621523292
transform 1 0 49588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_538
timestamp 1621523292
transform 1 0 50600 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_543
timestamp 1621523292
transform 1 0 51060 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0611_
timestamp 1621523292
transform 1 0 51428 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1621523292
transform 1 0 53176 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0800_
timestamp 1621523292
transform 1 0 52164 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_50_550
timestamp 1621523292
transform 1 0 51704 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_554
timestamp 1621523292
transform 1 0 52072 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_562
timestamp 1621523292
transform 1 0 52808 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1621523292
transform 1 0 54280 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_569
timestamp 1621523292
transform 1 0 53452 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_577
timestamp 1621523292
transform 1 0 54188 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1289_
timestamp 1621523292
transform 1 0 56856 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1621523292
transform 1 0 56212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_594
timestamp 1621523292
transform 1 0 55752 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_598
timestamp 1621523292
transform 1 0 56120 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_600
timestamp 1621523292
transform 1 0 56304 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1621523292
transform 1 0 57960 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1621523292
transform -1 0 58880 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_614
timestamp 1621523292
transform 1 0 57592 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1621523292
transform 1 0 58236 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1621523292
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output312
timestamp 1621523292
transform 1 0 1748 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_3
timestamp 1621523292
transform 1 0 1380 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_11
timestamp 1621523292
transform 1 0 2116 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_23
timestamp 1621523292
transform 1 0 3220 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_35
timestamp 1621523292
transform 1 0 4324 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1621523292
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_47
timestamp 1621523292
transform 1 0 5428 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_55
timestamp 1621523292
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1621523292
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1621523292
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_82
timestamp 1621523292
transform 1 0 8648 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_94
timestamp 1621523292
transform 1 0 9752 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_106
timestamp 1621523292
transform 1 0 10856 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1621523292
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_115
timestamp 1621523292
transform 1 0 11684 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_127
timestamp 1621523292
transform 1 0 12788 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_139
timestamp 1621523292
transform 1 0 13892 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_151
timestamp 1621523292
transform 1 0 14996 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1621523292
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_163
timestamp 1621523292
transform 1 0 16100 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_172
timestamp 1621523292
transform 1 0 16928 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1621523292
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1621523292
transform 1 0 19136 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1621523292
transform 1 0 20240 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1621523292
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_220
timestamp 1621523292
transform 1 0 21344 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_229
timestamp 1621523292
transform 1 0 22172 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_241
timestamp 1621523292
transform 1 0 23276 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_253
timestamp 1621523292
transform 1 0 24380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_265
timestamp 1621523292
transform 1 0 25484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_277
timestamp 1621523292
transform 1 0 26588 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1621523292
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_286
timestamp 1621523292
transform 1 0 27416 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_298
timestamp 1621523292
transform 1 0 28520 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1621523292
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1621523292
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1621523292
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_334
timestamp 1621523292
transform 1 0 31832 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1621523292
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1621523292
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1621523292
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1621523292
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_391
timestamp 1621523292
transform 1 0 37076 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1621523292
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_400
timestamp 1621523292
transform 1 0 37904 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_412
timestamp 1621523292
transform 1 0 39008 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_424
timestamp 1621523292
transform 1 0 40112 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_436
timestamp 1621523292
transform 1 0 41216 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1621523292
transform 1 0 43056 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_448
timestamp 1621523292
transform 1 0 42320 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_457
timestamp 1621523292
transform 1 0 43148 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_469
timestamp 1621523292
transform 1 0 44252 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_481
timestamp 1621523292
transform 1 0 45356 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_493
timestamp 1621523292
transform 1 0 46460 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1621523292
transform 1 0 48300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1621523292
transform 1 0 48852 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1621523292
transform 1 0 47564 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_514
timestamp 1621523292
transform 1 0 48392 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_518
timestamp 1621523292
transform 1 0 48760 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_522
timestamp 1621523292
transform 1 0 49128 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1621523292
transform 1 0 49496 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_542
timestamp 1621523292
transform 1 0 50968 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1621523292
transform 1 0 51888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0760_
timestamp 1621523292
transform 1 0 52532 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_51_550
timestamp 1621523292
transform 1 0 51704 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_555
timestamp 1621523292
transform 1 0 52164 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_566
timestamp 1621523292
transform 1 0 53176 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0609_
timestamp 1621523292
transform 1 0 55016 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0811_
timestamp 1621523292
transform 1 0 54004 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1621523292
transform 1 0 53544 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_571
timestamp 1621523292
transform 1 0 53636 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_582
timestamp 1621523292
transform 1 0 54648 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_589
timestamp 1621523292
transform 1 0 55292 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0610_
timestamp 1621523292
transform 1 0 55660 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1621523292
transform 1 0 56488 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_596
timestamp 1621523292
transform 1 0 55936 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_51_606
timestamp 1621523292
transform 1 0 56856 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _1327_
timestamp 1621523292
transform 1 0 57500 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1621523292
transform -1 0 58880 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_612
timestamp 1621523292
transform 1 0 57408 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_621
timestamp 1621523292
transform 1 0 58236 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1621523292
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1621523292
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1621523292
transform 1 0 1380 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1621523292
transform 1 0 1380 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_6
timestamp 1621523292
transform 1 0 1656 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_18
timestamp 1621523292
transform 1 0 2760 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_6
timestamp 1621523292
transform 1 0 1656 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_18
timestamp 1621523292
transform 1 0 2760 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1621523292
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_26
timestamp 1621523292
transform 1 0 3496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1621523292
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1621523292
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_30
timestamp 1621523292
transform 1 0 3864 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_42
timestamp 1621523292
transform 1 0 4968 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1621523292
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1621523292
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_54
timestamp 1621523292
transform 1 0 6072 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1621523292
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1621523292
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1621523292
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1621523292
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1621523292
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1621523292
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1621523292
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_99
timestamp 1621523292
transform 1 0 10212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1621523292
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1621523292
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1621523292
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_111
timestamp 1621523292
transform 1 0 11316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_123
timestamp 1621523292
transform 1 0 12420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_115
timestamp 1621523292
transform 1 0 11684 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_127
timestamp 1621523292
transform 1 0 12788 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1621523292
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_135
timestamp 1621523292
transform 1 0 13524 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_144
timestamp 1621523292
transform 1 0 14352 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_139
timestamp 1621523292
transform 1 0 13892 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_151
timestamp 1621523292
transform 1 0 14996 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1621523292
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_156
timestamp 1621523292
transform 1 0 15456 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_168
timestamp 1621523292
transform 1 0 16560 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_163
timestamp 1621523292
transform 1 0 16100 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_172
timestamp 1621523292
transform 1 0 16928 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_180
timestamp 1621523292
transform 1 0 17664 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_192
timestamp 1621523292
transform 1 0 18768 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1621523292
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1621523292
transform 1 0 19136 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1621523292
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_201
timestamp 1621523292
transform 1 0 19596 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_213
timestamp 1621523292
transform 1 0 20700 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_208
timestamp 1621523292
transform 1 0 20240 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1621523292
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_225
timestamp 1621523292
transform 1 0 21804 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_237
timestamp 1621523292
transform 1 0 22908 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_220
timestamp 1621523292
transform 1 0 21344 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_229
timestamp 1621523292
transform 1 0 22172 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1621523292
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_249
timestamp 1621523292
transform 1 0 24012 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_258
timestamp 1621523292
transform 1 0 24840 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_241
timestamp 1621523292
transform 1 0 23276 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_253
timestamp 1621523292
transform 1 0 24380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1621523292
transform 1 0 25944 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_282
timestamp 1621523292
transform 1 0 27048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_265
timestamp 1621523292
transform 1 0 25484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1621523292
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1621523292
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_294
timestamp 1621523292
transform 1 0 28152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_286
timestamp 1621523292
transform 1 0 27416 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_298
timestamp 1621523292
transform 1 0 28520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1621523292
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_306
timestamp 1621523292
transform 1 0 29256 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1621523292
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1621523292
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_310
timestamp 1621523292
transform 1 0 29624 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_322
timestamp 1621523292
transform 1 0 30728 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1621523292
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1621523292
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_334
timestamp 1621523292
transform 1 0 31832 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1621523292
transform 1 0 32660 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1621523292
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1621523292
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1621523292
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1621523292
transform 1 0 33764 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1621523292
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1621523292
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1621523292
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1621523292
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1621523292
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1621523292
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_396
timestamp 1621523292
transform 1 0 37536 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_408
timestamp 1621523292
transform 1 0 38640 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_400
timestamp 1621523292
transform 1 0 37904 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1621523292
transform 1 0 39008 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1621523292
transform 1 0 40480 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_420
timestamp 1621523292
transform 1 0 39744 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1621523292
transform 1 0 40572 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_424
timestamp 1621523292
transform 1 0 40112 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1621523292
transform 1 0 41216 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1621523292
transform 1 0 43056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1621523292
transform 1 0 41676 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_453
timestamp 1621523292
transform 1 0 42780 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_448
timestamp 1621523292
transform 1 0 42320 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_457
timestamp 1621523292
transform 1 0 43148 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_465
timestamp 1621523292
transform 1 0 43884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_477
timestamp 1621523292
transform 1 0 44988 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_469
timestamp 1621523292
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1621523292
transform 1 0 45724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_486
timestamp 1621523292
transform 1 0 45816 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_498
timestamp 1621523292
transform 1 0 46920 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_481
timestamp 1621523292
transform 1 0 45356 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_493
timestamp 1621523292
transform 1 0 46460 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1621523292
transform 1 0 48300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1621523292
transform 1 0 49312 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_510
timestamp 1621523292
transform 1 0 48024 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_522
timestamp 1621523292
transform 1 0 49128 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1621523292
transform 1 0 47564 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_514
timestamp 1621523292
transform 1 0 48392 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_522
timestamp 1621523292
transform 1 0 49128 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_527
timestamp 1621523292
transform 1 0 49588 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1621523292
transform 1 0 49680 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_531
timestamp 1621523292
transform 1 0 49956 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1621523292
transform 1 0 49956 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_534
timestamp 1621523292
transform 1 0 50232 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_538
timestamp 1621523292
transform 1 0 50600 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1183_
timestamp 1621523292
transform 1 0 50600 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1078_
timestamp 1621523292
transform 1 0 50324 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_541
timestamp 1621523292
transform 1 0 50876 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_543
timestamp 1621523292
transform 1 0 51060 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1621523292
transform 1 0 50968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0806_
timestamp 1621523292
transform 1 0 51244 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_549
timestamp 1621523292
transform 1 0 51612 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_551
timestamp 1621523292
transform 1 0 51796 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_547
timestamp 1621523292
transform 1 0 51428 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0947_
timestamp 1621523292
transform 1 0 51520 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_559
timestamp 1621523292
transform 1 0 52532 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_555
timestamp 1621523292
transform 1 0 52164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_563
timestamp 1621523292
transform 1 0 52900 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0946_
timestamp 1621523292
transform 1 0 52900 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0813_
timestamp 1621523292
transform 1 0 52164 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0809_
timestamp 1621523292
transform 1 0 52256 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_566
timestamp 1621523292
transform 1 0 53176 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_567
timestamp 1621523292
transform 1 0 53268 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_571
timestamp 1621523292
transform 1 0 53636 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_574
timestamp 1621523292
transform 1 0 53912 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1621523292
transform 1 0 53544 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _0810_
timestamp 1621523292
transform 1 0 53360 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0689_
timestamp 1621523292
transform 1 0 54280 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_585
timestamp 1621523292
transform 1 0 54924 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_585
timestamp 1621523292
transform 1 0 54924 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0762_
timestamp 1621523292
transform 1 0 54372 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0608_
timestamp 1621523292
transform 1 0 55292 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1621523292
transform 1 0 55292 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1621523292
transform 1 0 56212 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output224
timestamp 1621523292
transform 1 0 57132 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_592
timestamp 1621523292
transform 1 0 55568 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_598
timestamp 1621523292
transform 1 0 56120 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_600
timestamp 1621523292
transform 1 0 56304 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_608
timestamp 1621523292
transform 1 0 57040 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_605
timestamp 1621523292
transform 1 0 56764 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_611
timestamp 1621523292
transform 1 0 57316 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1290_
timestamp 1621523292
transform 1 0 57408 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1621523292
transform -1 0 58880 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1621523292
transform -1 0 58880 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output186
timestamp 1621523292
transform 1 0 57868 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1621523292
transform 1 0 57500 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1621523292
transform 1 0 58236 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_620
timestamp 1621523292
transform 1 0 58144 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_624
timestamp 1621523292
transform 1 0 58512 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1621523292
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1621523292
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1621523292
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1621523292
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_27
timestamp 1621523292
transform 1 0 3588 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1621523292
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1621523292
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1621523292
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1621523292
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1621523292
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1621523292
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1621523292
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1621523292
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1621523292
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_123
timestamp 1621523292
transform 1 0 12420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1621523292
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_135
timestamp 1621523292
transform 1 0 13524 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_144
timestamp 1621523292
transform 1 0 14352 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_156
timestamp 1621523292
transform 1 0 15456 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_168
timestamp 1621523292
transform 1 0 16560 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_180
timestamp 1621523292
transform 1 0 17664 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_192
timestamp 1621523292
transform 1 0 18768 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1621523292
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_201
timestamp 1621523292
transform 1 0 19596 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_213
timestamp 1621523292
transform 1 0 20700 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_225
timestamp 1621523292
transform 1 0 21804 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_237
timestamp 1621523292
transform 1 0 22908 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1621523292
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_249
timestamp 1621523292
transform 1 0 24012 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_258
timestamp 1621523292
transform 1 0 24840 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_270
timestamp 1621523292
transform 1 0 25944 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_282
timestamp 1621523292
transform 1 0 27048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_294
timestamp 1621523292
transform 1 0 28152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1621523292
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_306
timestamp 1621523292
transform 1 0 29256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1621523292
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_327
timestamp 1621523292
transform 1 0 31188 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_339
timestamp 1621523292
transform 1 0 32292 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1621523292
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_351
timestamp 1621523292
transform 1 0 33396 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_363
timestamp 1621523292
transform 1 0 34500 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_372
timestamp 1621523292
transform 1 0 35328 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_384
timestamp 1621523292
transform 1 0 36432 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_396
timestamp 1621523292
transform 1 0 37536 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_408
timestamp 1621523292
transform 1 0 38640 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1621523292
transform 1 0 40480 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_420
timestamp 1621523292
transform 1 0 39744 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1621523292
transform 1 0 40572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_441
timestamp 1621523292
transform 1 0 41676 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_453
timestamp 1621523292
transform 1 0 42780 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_465
timestamp 1621523292
transform 1 0 43884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_477
timestamp 1621523292
transform 1 0 44988 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1621523292
transform 1 0 45724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_486
timestamp 1621523292
transform 1 0 45816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_498
timestamp 1621523292
transform 1 0 46920 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_510
timestamp 1621523292
transform 1 0 48024 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_522
timestamp 1621523292
transform 1 0 49128 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _1184_
timestamp 1621523292
transform 1 0 50324 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1621523292
transform 1 0 50968 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1621523292
transform 1 0 49680 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_531
timestamp 1621523292
transform 1 0 49956 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_538
timestamp 1621523292
transform 1 0 50600 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_543
timestamp 1621523292
transform 1 0 51060 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0801_
timestamp 1621523292
transform 1 0 51704 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1621523292
transform 1 0 52716 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_54_549
timestamp 1621523292
transform 1 0 51612 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_557
timestamp 1621523292
transform 1 0 52348 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0761_
timestamp 1621523292
transform 1 0 54832 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_54_577
timestamp 1621523292
transform 1 0 54188 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_583
timestamp 1621523292
transform 1 0 54740 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1621523292
transform 1 0 56212 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output226
timestamp 1621523292
transform 1 0 57132 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_591
timestamp 1621523292
transform 1 0 55476 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_600
timestamp 1621523292
transform 1 0 56304 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_608
timestamp 1621523292
transform 1 0 57040 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1621523292
transform -1 0 58880 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output188
timestamp 1621523292
transform 1 0 57868 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1621523292
transform 1 0 57500 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_621
timestamp 1621523292
transform 1 0 58236 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1621523292
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1621523292
transform 1 0 1380 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_6
timestamp 1621523292
transform 1 0 1656 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_18
timestamp 1621523292
transform 1 0 2760 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_30
timestamp 1621523292
transform 1 0 3864 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_42
timestamp 1621523292
transform 1 0 4968 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1621523292
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_54
timestamp 1621523292
transform 1 0 6072 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1621523292
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1621523292
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1621523292
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1621523292
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1621523292
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1621523292
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1621523292
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1621523292
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_139
timestamp 1621523292
transform 1 0 13892 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_151
timestamp 1621523292
transform 1 0 14996 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1621523292
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_163
timestamp 1621523292
transform 1 0 16100 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_172
timestamp 1621523292
transform 1 0 16928 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1621523292
transform 1 0 18032 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1621523292
transform 1 0 19136 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1621523292
transform 1 0 20240 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1621523292
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_220
timestamp 1621523292
transform 1 0 21344 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_229
timestamp 1621523292
transform 1 0 22172 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_241
timestamp 1621523292
transform 1 0 23276 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_253
timestamp 1621523292
transform 1 0 24380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_265
timestamp 1621523292
transform 1 0 25484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_277
timestamp 1621523292
transform 1 0 26588 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1621523292
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1621523292
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1621523292
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1621523292
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1621523292
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1621523292
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_334
timestamp 1621523292
transform 1 0 31832 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1621523292
transform 1 0 32660 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1621523292
transform 1 0 33764 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1621523292
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1621523292
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_391
timestamp 1621523292
transform 1 0 37076 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1621523292
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_400
timestamp 1621523292
transform 1 0 37904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_412
timestamp 1621523292
transform 1 0 39008 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_424
timestamp 1621523292
transform 1 0 40112 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_436
timestamp 1621523292
transform 1 0 41216 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1621523292
transform 1 0 43056 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_448
timestamp 1621523292
transform 1 0 42320 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_457
timestamp 1621523292
transform 1 0 43148 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_469
timestamp 1621523292
transform 1 0 44252 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_481
timestamp 1621523292
transform 1 0 45356 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_493
timestamp 1621523292
transform 1 0 46460 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1621523292
transform 1 0 48300 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1621523292
transform 1 0 47564 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_514
timestamp 1621523292
transform 1 0 48392 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0802_
timestamp 1621523292
transform 1 0 50876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_526
timestamp 1621523292
transform 1 0 49496 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_538
timestamp 1621523292
transform 1 0 50600 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_544
timestamp 1621523292
transform 1 0 51152 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1621523292
transform 1 0 52900 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0807_
timestamp 1621523292
transform 1 0 51520 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_556
timestamp 1621523292
transform 1 0 52256 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_562
timestamp 1621523292
transform 1 0 52808 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_566
timestamp 1621523292
transform 1 0 53176 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0766_
timestamp 1621523292
transform 1 0 54004 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1621523292
transform 1 0 55292 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1621523292
transform 1 0 53544 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_571
timestamp 1621523292
transform 1 0 53636 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_582
timestamp 1621523292
transform 1 0 54648 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_588
timestamp 1621523292
transform 1 0 55200 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_605
timestamp 1621523292
transform 1 0 56764 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1328_
timestamp 1621523292
transform 1 0 57500 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1621523292
transform -1 0 58880 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1621523292
transform 1 0 58236 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1621523292
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1621523292
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1621523292
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1621523292
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1621523292
transform 1 0 3588 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1621523292
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1621523292
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1621523292
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1621523292
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1621523292
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1621523292
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1621523292
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1621523292
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1621523292
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1621523292
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1621523292
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1621523292
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1621523292
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1621523292
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1621523292
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1621523292
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1621523292
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1621523292
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_201
timestamp 1621523292
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_213
timestamp 1621523292
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_225
timestamp 1621523292
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1621523292
transform 1 0 22908 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1621523292
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_249
timestamp 1621523292
transform 1 0 24012 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_258
timestamp 1621523292
transform 1 0 24840 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_270
timestamp 1621523292
transform 1 0 25944 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_282
timestamp 1621523292
transform 1 0 27048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_294
timestamp 1621523292
transform 1 0 28152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1621523292
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_306
timestamp 1621523292
transform 1 0 29256 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1621523292
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_327
timestamp 1621523292
transform 1 0 31188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_339
timestamp 1621523292
transform 1 0 32292 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1621523292
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_351
timestamp 1621523292
transform 1 0 33396 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_363
timestamp 1621523292
transform 1 0 34500 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1621523292
transform 1 0 35328 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1621523292
transform 1 0 36432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_396
timestamp 1621523292
transform 1 0 37536 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_408
timestamp 1621523292
transform 1 0 38640 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1621523292
transform 1 0 40480 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_420
timestamp 1621523292
transform 1 0 39744 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1621523292
transform 1 0 40572 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_441
timestamp 1621523292
transform 1 0 41676 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_453
timestamp 1621523292
transform 1 0 42780 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_465
timestamp 1621523292
transform 1 0 43884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_477
timestamp 1621523292
transform 1 0 44988 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1621523292
transform 1 0 45724 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_486
timestamp 1621523292
transform 1 0 45816 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_498
timestamp 1621523292
transform 1 0 46920 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_510
timestamp 1621523292
transform 1 0 48024 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_522
timestamp 1621523292
transform 1 0 49128 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0900_
timestamp 1621523292
transform 1 0 50324 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1621523292
transform 1 0 50968 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1621523292
transform 1 0 49680 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_531
timestamp 1621523292
transform 1 0 49956 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_538
timestamp 1621523292
transform 1 0 50600 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_543
timestamp 1621523292
transform 1 0 51060 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0694_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 53268 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1621523292
transform 1 0 51428 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_56_563
timestamp 1621523292
transform 1 0 52900 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0607_
timestamp 1621523292
transform 1 0 54280 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0687_
timestamp 1621523292
transform 1 0 54924 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_56_574
timestamp 1621523292
transform 1 0 53912 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_581
timestamp 1621523292
transform 1 0 54556 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1291_
timestamp 1621523292
transform 1 0 57132 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1621523292
transform 1 0 56212 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_592
timestamp 1621523292
transform 1 0 55568 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_598
timestamp 1621523292
transform 1 0 56120 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_600
timestamp 1621523292
transform 1 0 56304 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_608
timestamp 1621523292
transform 1 0 57040 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1621523292
transform -1 0 58880 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_617
timestamp 1621523292
transform 1 0 57868 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1621523292
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1621523292
transform 1 0 1380 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_6
timestamp 1621523292
transform 1 0 1656 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_18
timestamp 1621523292
transform 1 0 2760 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1621523292
transform 1 0 3864 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1621523292
transform 1 0 4968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1621523292
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_54
timestamp 1621523292
transform 1 0 6072 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1621523292
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1621523292
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1621523292
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1621523292
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1621523292
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1621523292
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1621523292
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1621523292
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1621523292
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1621523292
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1621523292
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1621523292
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1621523292
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1621523292
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1621523292
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1621523292
transform 1 0 20240 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1621523292
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_220
timestamp 1621523292
transform 1 0 21344 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1621523292
transform 1 0 22172 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1621523292
transform 1 0 23276 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_253
timestamp 1621523292
transform 1 0 24380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_265
timestamp 1621523292
transform 1 0 25484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_277
timestamp 1621523292
transform 1 0 26588 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1621523292
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1621523292
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1621523292
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1621523292
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1621523292
transform 1 0 30728 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1621523292
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_334
timestamp 1621523292
transform 1 0 31832 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1621523292
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_355
timestamp 1621523292
transform 1 0 33764 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1621523292
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1621523292
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_391
timestamp 1621523292
transform 1 0 37076 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1621523292
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_400
timestamp 1621523292
transform 1 0 37904 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_412
timestamp 1621523292
transform 1 0 39008 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_424
timestamp 1621523292
transform 1 0 40112 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_436
timestamp 1621523292
transform 1 0 41216 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1621523292
transform 1 0 43056 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_448
timestamp 1621523292
transform 1 0 42320 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_457
timestamp 1621523292
transform 1 0 43148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_469
timestamp 1621523292
transform 1 0 44252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_481
timestamp 1621523292
transform 1 0 45356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_493
timestamp 1621523292
transform 1 0 46460 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1621523292
transform 1 0 48300 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1621523292
transform 1 0 47564 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_514
timestamp 1621523292
transform 1 0 48392 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _0634_
timestamp 1621523292
transform 1 0 50876 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1080_
timestamp 1621523292
transform 1 0 50232 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1185_
timestamp 1621523292
transform 1 0 49588 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_526
timestamp 1621523292
transform 1 0 49496 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_530
timestamp 1621523292
transform 1 0 49864 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_537
timestamp 1621523292
transform 1 0 50508 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_545
timestamp 1621523292
transform 1 0 51244 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0605_
timestamp 1621523292
transform 1 0 51888 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0764_
timestamp 1621523292
transform 1 0 52532 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_57_551
timestamp 1621523292
transform 1 0 51796 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_555
timestamp 1621523292
transform 1 0 52164 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_566
timestamp 1621523292
transform 1 0 53176 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0763_
timestamp 1621523292
transform 1 0 54004 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0765_
timestamp 1621523292
transform 1 0 55016 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1621523292
transform 1 0 53544 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_571
timestamp 1621523292
transform 1 0 53636 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_582
timestamp 1621523292
transform 1 0 54648 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0606_
timestamp 1621523292
transform 1 0 56028 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output227
timestamp 1621523292
transform 1 0 57132 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_593
timestamp 1621523292
transform 1 0 55660 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_600
timestamp 1621523292
transform 1 0 56304 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_608
timestamp 1621523292
transform 1 0 57040 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1621523292
transform -1 0 58880 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output189
timestamp 1621523292
transform 1 0 57868 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_613
timestamp 1621523292
transform 1 0 57500 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1621523292
transform 1 0 58236 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1621523292
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1621523292
transform 1 0 1380 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_6
timestamp 1621523292
transform 1 0 1656 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_18
timestamp 1621523292
transform 1 0 2760 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1621523292
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_26
timestamp 1621523292
transform 1 0 3496 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1621523292
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1621523292
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1621523292
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1621523292
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1621523292
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1621523292
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_87
timestamp 1621523292
transform 1 0 9108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_99
timestamp 1621523292
transform 1 0 10212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_111
timestamp 1621523292
transform 1 0 11316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1621523292
transform 1 0 12420 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1621523292
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1621523292
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1621523292
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1621523292
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1621523292
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1621523292
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1621523292
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1621523292
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1621523292
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_213
timestamp 1621523292
transform 1 0 20700 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_225
timestamp 1621523292
transform 1 0 21804 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_237
timestamp 1621523292
transform 1 0 22908 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1621523292
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_249
timestamp 1621523292
transform 1 0 24012 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1621523292
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1621523292
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1621523292
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1621523292
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1621523292
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1621523292
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_315
timestamp 1621523292
transform 1 0 30084 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_327
timestamp 1621523292
transform 1 0 31188 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_339
timestamp 1621523292
transform 1 0 32292 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1621523292
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_351
timestamp 1621523292
transform 1 0 33396 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_363
timestamp 1621523292
transform 1 0 34500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_372
timestamp 1621523292
transform 1 0 35328 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_384
timestamp 1621523292
transform 1 0 36432 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_396
timestamp 1621523292
transform 1 0 37536 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_408
timestamp 1621523292
transform 1 0 38640 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1621523292
transform 1 0 40480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_420
timestamp 1621523292
transform 1 0 39744 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_429
timestamp 1621523292
transform 1 0 40572 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_441
timestamp 1621523292
transform 1 0 41676 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_453
timestamp 1621523292
transform 1 0 42780 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_465
timestamp 1621523292
transform 1 0 43884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_477
timestamp 1621523292
transform 1 0 44988 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1621523292
transform 1 0 45724 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1621523292
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1621523292
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_510
timestamp 1621523292
transform 1 0 48024 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_522
timestamp 1621523292
transform 1 0 49128 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 1621523292
transform 1 0 50324 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1621523292
transform 1 0 50968 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1621523292
transform 1 0 49680 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_531
timestamp 1621523292
transform 1 0 49956 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_538
timestamp 1621523292
transform 1 0 50600 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_543
timestamp 1621523292
transform 1 0 51060 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0693_
timestamp 1621523292
transform 1 0 52808 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0803_
timestamp 1621523292
transform 1 0 51888 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_551
timestamp 1621523292
transform 1 0 51796 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_558
timestamp 1621523292
transform 1 0 52440 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1621523292
transform 1 0 54372 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_58_569
timestamp 1621523292
transform 1 0 53452 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_577
timestamp 1621523292
transform 1 0 54188 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1621523292
transform 1 0 56672 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1621523292
transform 1 0 56212 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_595
timestamp 1621523292
transform 1 0 55844 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_600
timestamp 1621523292
transform 1 0 56304 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_608
timestamp 1621523292
transform 1 0 57040 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1329_
timestamp 1621523292
transform 1 0 57500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1621523292
transform -1 0 58880 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_58_612
timestamp 1621523292
transform 1 0 57408 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_621
timestamp 1621523292
transform 1 0 58236 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1621523292
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1621523292
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1621523292
transform 1 0 1380 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1621523292
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1621523292
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_6
timestamp 1621523292
transform 1 0 1656 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_18
timestamp 1621523292
transform 1 0 2760 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1621523292
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1621523292
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1621523292
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_26
timestamp 1621523292
transform 1 0 3496 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1621523292
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1621523292
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1621523292
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_51
timestamp 1621523292
transform 1 0 5796 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1621523292
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1621523292
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1621523292
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1621523292
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1621523292
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1621523292
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1621523292
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1621523292
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1621523292
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1621523292
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1621523292
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1621523292
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1621523292
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1621523292
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1621523292
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1621523292
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1621523292
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1621523292
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1621523292
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1621523292
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1621523292
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1621523292
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1621523292
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1621523292
transform 1 0 16928 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1621523292
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1621523292
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1621523292
transform 1 0 18032 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1621523292
transform 1 0 19136 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1621523292
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1621523292
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1621523292
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_208
timestamp 1621523292
transform 1 0 20240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_201
timestamp 1621523292
transform 1 0 19596 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_213
timestamp 1621523292
transform 1 0 20700 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1621523292
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_220
timestamp 1621523292
transform 1 0 21344 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_229
timestamp 1621523292
transform 1 0 22172 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_225
timestamp 1621523292
transform 1 0 21804 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_237
timestamp 1621523292
transform 1 0 22908 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1621523292
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_241
timestamp 1621523292
transform 1 0 23276 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_253
timestamp 1621523292
transform 1 0 24380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_249
timestamp 1621523292
transform 1 0 24012 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1621523292
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1621523292
transform 1 0 25484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_277
timestamp 1621523292
transform 1 0 26588 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1621523292
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1621523292
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1621523292
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1621523292
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1621523292
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1621523292
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1621523292
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_310
timestamp 1621523292
transform 1 0 29624 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_322
timestamp 1621523292
transform 1 0 30728 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1621523292
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_315
timestamp 1621523292
transform 1 0 30084 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_327
timestamp 1621523292
transform 1 0 31188 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1621523292
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_334
timestamp 1621523292
transform 1 0 31832 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_343
timestamp 1621523292
transform 1 0 32660 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_339
timestamp 1621523292
transform 1 0 32292 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1621523292
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_355
timestamp 1621523292
transform 1 0 33764 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1621523292
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_351
timestamp 1621523292
transform 1 0 33396 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_363
timestamp 1621523292
transform 1 0 34500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1621523292
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_391
timestamp 1621523292
transform 1 0 37076 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1621523292
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1621523292
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1621523292
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_400
timestamp 1621523292
transform 1 0 37904 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_412
timestamp 1621523292
transform 1 0 39008 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_396
timestamp 1621523292
transform 1 0 37536 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_408
timestamp 1621523292
transform 1 0 38640 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1621523292
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_424
timestamp 1621523292
transform 1 0 40112 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_436
timestamp 1621523292
transform 1 0 41216 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_420
timestamp 1621523292
transform 1 0 39744 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_429
timestamp 1621523292
transform 1 0 40572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1621523292
transform 1 0 43056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_448
timestamp 1621523292
transform 1 0 42320 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1621523292
transform 1 0 43148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_441
timestamp 1621523292
transform 1 0 41676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_453
timestamp 1621523292
transform 1 0 42780 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1621523292
transform 1 0 44252 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_465
timestamp 1621523292
transform 1 0 43884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_477
timestamp 1621523292
transform 1 0 44988 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1621523292
transform 1 0 45724 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_481
timestamp 1621523292
transform 1 0 45356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_493
timestamp 1621523292
transform 1 0 46460 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_486
timestamp 1621523292
transform 1 0 45816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_498
timestamp 1621523292
transform 1 0 46920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1621523292
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1621523292
transform 1 0 47564 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_514
timestamp 1621523292
transform 1 0 48392 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_510
timestamp 1621523292
transform 1 0 48024 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_522
timestamp 1621523292
transform 1 0 49128 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_531
timestamp 1621523292
transform 1 0 49956 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_529
timestamp 1621523292
transform 1 0 49772 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1186_
timestamp 1621523292
transform 1 0 49496 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1621523292
transform 1 0 49680 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_538
timestamp 1621523292
transform 1 0 50600 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_537
timestamp 1621523292
transform 1 0 50508 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0943_
timestamp 1621523292
transform 1 0 50324 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0589_
timestamp 1621523292
transform 1 0 50140 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0588_
timestamp 1621523292
transform 1 0 50876 0 1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_60_543
timestamp 1621523292
transform 1 0 51060 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1621523292
transform 1 0 50968 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _0782_
timestamp 1621523292
transform 1 0 52716 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _0804_
timestamp 1621523292
transform 1 0 51704 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1621523292
transform 1 0 51796 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_59_546
timestamp 1621523292
transform 1 0 51336 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_557
timestamp 1621523292
transform 1 0 52348 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_565
timestamp 1621523292
transform 1 0 53084 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_567
timestamp 1621523292
transform 1 0 53268 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_574
timestamp 1621523292
transform 1 0 53912 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_571
timestamp 1621523292
transform 1 0 53636 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_569
timestamp 1621523292
transform 1 0 53452 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1621523292
transform 1 0 53544 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0691_
timestamp 1621523292
transform 1 0 54004 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0603_
timestamp 1621523292
transform 1 0 53636 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_589
timestamp 1621523292
transform 1 0 55292 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_582
timestamp 1621523292
transform 1 0 54648 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0604_
timestamp 1621523292
transform 1 0 55016 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1621523292
transform 1 0 54280 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_598
timestamp 1621523292
transform 1 0 56120 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_594
timestamp 1621523292
transform 1 0 55752 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_597
timestamp 1621523292
transform 1 0 56028 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output228
timestamp 1621523292
transform 1 0 56120 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_604
timestamp 1621523292
transform 1 0 56672 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_600
timestamp 1621523292
transform 1 0 56304 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_602
timestamp 1621523292
transform 1 0 56488 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output190
timestamp 1621523292
transform 1 0 56764 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1621523292
transform 1 0 56212 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1292_
timestamp 1621523292
transform 1 0 56856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_609
timestamp 1621523292
transform 1 0 57132 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1621523292
transform 1 0 57960 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1330_
timestamp 1621523292
transform 1 0 57500 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1621523292
transform -1 0 58880 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1621523292
transform -1 0 58880 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_614
timestamp 1621523292
transform 1 0 57592 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_621
timestamp 1621523292
transform 1 0 58236 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1621523292
transform 1 0 58236 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1621523292
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1621523292
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1621523292
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1621523292
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1621523292
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1621523292
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_51
timestamp 1621523292
transform 1 0 5796 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1621523292
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1621523292
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1621523292
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1621523292
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1621523292
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1621523292
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1621523292
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1621523292
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1621523292
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1621523292
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1621523292
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1621523292
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_172
timestamp 1621523292
transform 1 0 16928 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1621523292
transform 1 0 18032 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1621523292
transform 1 0 19136 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1621523292
transform 1 0 20240 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1621523292
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_220
timestamp 1621523292
transform 1 0 21344 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1621523292
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1621523292
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1621523292
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1621523292
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1621523292
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1621523292
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1621523292
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1621523292
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1621523292
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_322
timestamp 1621523292
transform 1 0 30728 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1621523292
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_334
timestamp 1621523292
transform 1 0 31832 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_343
timestamp 1621523292
transform 1 0 32660 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_355
timestamp 1621523292
transform 1 0 33764 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1621523292
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1621523292
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_391
timestamp 1621523292
transform 1 0 37076 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1621523292
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_400
timestamp 1621523292
transform 1 0 37904 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_412
timestamp 1621523292
transform 1 0 39008 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_424
timestamp 1621523292
transform 1 0 40112 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_436
timestamp 1621523292
transform 1 0 41216 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1621523292
transform 1 0 43056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_448
timestamp 1621523292
transform 1 0 42320 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_457
timestamp 1621523292
transform 1 0 43148 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_469
timestamp 1621523292
transform 1 0 44252 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_481
timestamp 1621523292
transform 1 0 45356 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_493
timestamp 1621523292
transform 1 0 46460 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1621523292
transform 1 0 48300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1621523292
transform 1 0 47564 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_514
timestamp 1621523292
transform 1 0 48392 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1621523292
transform 1 0 50968 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0942_
timestamp 1621523292
transform 1 0 50324 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1621523292
transform 1 0 49680 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_526
timestamp 1621523292
transform 1 0 49496 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_531
timestamp 1621523292
transform 1 0 49956 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_538
timestamp 1621523292
transform 1 0 50600 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_545
timestamp 1621523292
transform 1 0 51244 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0805_
timestamp 1621523292
transform 1 0 51704 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0897_
timestamp 1621523292
transform 1 0 52900 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_549
timestamp 1621523292
transform 1 0 51612 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_553
timestamp 1621523292
transform 1 0 51980 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_561
timestamp 1621523292
transform 1 0 52716 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_566
timestamp 1621523292
transform 1 0 53176 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0590_
timestamp 1621523292
transform 1 0 54372 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0601_
timestamp 1621523292
transform 1 0 55108 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1621523292
transform 1 0 53544 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_571
timestamp 1621523292
transform 1 0 53636 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_583
timestamp 1621523292
transform 1 0 54740 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1621523292
transform 1 0 56120 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1293_
timestamp 1621523292
transform 1 0 56856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_591
timestamp 1621523292
transform 1 0 55476 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_597
timestamp 1621523292
transform 1 0 56028 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_602
timestamp 1621523292
transform 1 0 56488 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0895_
timestamp 1621523292
transform 1 0 57960 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1621523292
transform -1 0 58880 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_614
timestamp 1621523292
transform 1 0 57592 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_621
timestamp 1621523292
transform 1 0 58236 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1621523292
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1621523292
transform 1 0 1380 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_6
timestamp 1621523292
transform 1 0 1656 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 1621523292
transform 1 0 2760 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1621523292
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_26
timestamp 1621523292
transform 1 0 3496 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1621523292
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1621523292
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1621523292
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1621523292
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1621523292
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_78
timestamp 1621523292
transform 1 0 8280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1621523292
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1621523292
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1621523292
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1621523292
transform 1 0 12420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1621523292
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1621523292
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1621523292
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_156
timestamp 1621523292
transform 1 0 15456 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_168
timestamp 1621523292
transform 1 0 16560 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_180
timestamp 1621523292
transform 1 0 17664 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_192
timestamp 1621523292
transform 1 0 18768 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1621523292
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1621523292
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1621523292
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1621523292
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1621523292
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1621523292
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1621523292
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1621523292
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1621523292
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_282
timestamp 1621523292
transform 1 0 27048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_294
timestamp 1621523292
transform 1 0 28152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1621523292
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_306
timestamp 1621523292
transform 1 0 29256 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_315
timestamp 1621523292
transform 1 0 30084 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_327
timestamp 1621523292
transform 1 0 31188 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_339
timestamp 1621523292
transform 1 0 32292 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1621523292
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_351
timestamp 1621523292
transform 1 0 33396 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_363
timestamp 1621523292
transform 1 0 34500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1621523292
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1621523292
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_396
timestamp 1621523292
transform 1 0 37536 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_408
timestamp 1621523292
transform 1 0 38640 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1621523292
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_420
timestamp 1621523292
transform 1 0 39744 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_429
timestamp 1621523292
transform 1 0 40572 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_441
timestamp 1621523292
transform 1 0 41676 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_453
timestamp 1621523292
transform 1 0 42780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_465
timestamp 1621523292
transform 1 0 43884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1621523292
transform 1 0 44988 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1621523292
transform 1 0 45724 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1621523292
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_498
timestamp 1621523292
transform 1 0 46920 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_510
timestamp 1621523292
transform 1 0 48024 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_522
timestamp 1621523292
transform 1 0 49128 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1187_
timestamp 1621523292
transform 1 0 50324 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1621523292
transform 1 0 50968 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_534
timestamp 1621523292
transform 1 0 50232 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_538
timestamp 1621523292
transform 1 0 50600 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_543
timestamp 1621523292
transform 1 0 51060 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0779_
timestamp 1621523292
transform 1 0 51428 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0796_
timestamp 1621523292
transform 1 0 52440 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_551
timestamp 1621523292
transform 1 0 51796 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_557
timestamp 1621523292
transform 1 0 52348 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_564
timestamp 1621523292
transform 1 0 52992 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0602_
timestamp 1621523292
transform 1 0 54556 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0667_
timestamp 1621523292
transform 1 0 53544 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_62_577
timestamp 1621523292
transform 1 0 54188 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_584
timestamp 1621523292
transform 1 0 54832 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1621523292
transform 1 0 55568 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1621523292
transform 1 0 56212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output229
timestamp 1621523292
transform 1 0 56764 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_595
timestamp 1621523292
transform 1 0 55844 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_600
timestamp 1621523292
transform 1 0 56304 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_604
timestamp 1621523292
transform 1 0 56672 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_609
timestamp 1621523292
transform 1 0 57132 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1331_
timestamp 1621523292
transform 1 0 57500 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1621523292
transform -1 0 58880 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1621523292
transform 1 0 58236 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1621523292
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1621523292
transform 1 0 1380 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_6
timestamp 1621523292
transform 1 0 1656 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_18
timestamp 1621523292
transform 1 0 2760 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1621523292
transform 1 0 3864 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1621523292
transform 1 0 4968 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1621523292
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_54
timestamp 1621523292
transform 1 0 6072 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1621523292
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1621523292
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1621523292
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1621523292
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1621523292
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1621523292
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1621523292
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1621523292
transform 1 0 12788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_139
timestamp 1621523292
transform 1 0 13892 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_151
timestamp 1621523292
transform 1 0 14996 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1621523292
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_163
timestamp 1621523292
transform 1 0 16100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_172
timestamp 1621523292
transform 1 0 16928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1621523292
transform 1 0 18032 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1621523292
transform 1 0 19136 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1621523292
transform 1 0 20240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1621523292
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_220
timestamp 1621523292
transform 1 0 21344 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1621523292
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1621523292
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1621523292
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1621523292
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1621523292
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1621523292
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_286
timestamp 1621523292
transform 1 0 27416 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_298
timestamp 1621523292
transform 1 0 28520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_310
timestamp 1621523292
transform 1 0 29624 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_322
timestamp 1621523292
transform 1 0 30728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1621523292
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_334
timestamp 1621523292
transform 1 0 31832 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1621523292
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_355
timestamp 1621523292
transform 1 0 33764 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1621523292
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1621523292
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_391
timestamp 1621523292
transform 1 0 37076 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1621523292
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1621523292
transform 1 0 37904 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1621523292
transform 1 0 39008 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1621523292
transform 1 0 40112 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_436
timestamp 1621523292
transform 1 0 41216 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1621523292
transform 1 0 43056 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_448
timestamp 1621523292
transform 1 0 42320 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_457
timestamp 1621523292
transform 1 0 43148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_469
timestamp 1621523292
transform 1 0 44252 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_481
timestamp 1621523292
transform 1 0 45356 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_493
timestamp 1621523292
transform 1 0 46460 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1621523292
transform 1 0 48300 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1621523292
transform 1 0 47564 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_514
timestamp 1621523292
transform 1 0 48392 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1621523292
transform 1 0 50048 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_63_526
timestamp 1621523292
transform 1 0 49496 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0799_
timestamp 1621523292
transform 1 0 52256 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_548
timestamp 1621523292
transform 1 0 51520 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_564
timestamp 1621523292
transform 1 0 52992 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0600_
timestamp 1621523292
transform 1 0 54004 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1621523292
transform 1 0 54740 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1621523292
transform 1 0 53544 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_571
timestamp 1621523292
transform 1 0 53636 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_578
timestamp 1621523292
transform 1 0 54280 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_582
timestamp 1621523292
transform 1 0 54648 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1621523292
transform 1 0 56580 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0896_
timestamp 1621523292
transform 1 0 57224 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_599
timestamp 1621523292
transform 1 0 56212 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_606
timestamp 1621523292
transform 1 0 56856 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1621523292
transform -1 0 58880 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output191
timestamp 1621523292
transform 1 0 57868 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_613
timestamp 1621523292
transform 1 0 57500 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_621
timestamp 1621523292
transform 1 0 58236 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1621523292
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1621523292
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1621523292
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1621523292
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_27
timestamp 1621523292
transform 1 0 3588 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1621523292
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1621523292
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1621523292
transform 1 0 6072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1621523292
transform 1 0 9016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_66
timestamp 1621523292
transform 1 0 7176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_78
timestamp 1621523292
transform 1 0 8280 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_87
timestamp 1621523292
transform 1 0 9108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_99
timestamp 1621523292
transform 1 0 10212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_111
timestamp 1621523292
transform 1 0 11316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_123
timestamp 1621523292
transform 1 0 12420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1621523292
transform 1 0 14260 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_135
timestamp 1621523292
transform 1 0 13524 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_144
timestamp 1621523292
transform 1 0 14352 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_156
timestamp 1621523292
transform 1 0 15456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_168
timestamp 1621523292
transform 1 0 16560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_180
timestamp 1621523292
transform 1 0 17664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_192
timestamp 1621523292
transform 1 0 18768 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1621523292
transform 1 0 19504 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_201
timestamp 1621523292
transform 1 0 19596 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_213
timestamp 1621523292
transform 1 0 20700 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1621523292
transform 1 0 21804 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_237
timestamp 1621523292
transform 1 0 22908 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1621523292
transform 1 0 24748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_249
timestamp 1621523292
transform 1 0 24012 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_258
timestamp 1621523292
transform 1 0 24840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_270
timestamp 1621523292
transform 1 0 25944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_282
timestamp 1621523292
transform 1 0 27048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_294
timestamp 1621523292
transform 1 0 28152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1621523292
transform 1 0 29992 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_306
timestamp 1621523292
transform 1 0 29256 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_315
timestamp 1621523292
transform 1 0 30084 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_327
timestamp 1621523292
transform 1 0 31188 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_339
timestamp 1621523292
transform 1 0 32292 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1621523292
transform 1 0 35236 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_351
timestamp 1621523292
transform 1 0 33396 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_363
timestamp 1621523292
transform 1 0 34500 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_372
timestamp 1621523292
transform 1 0 35328 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1621523292
transform 1 0 36432 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_396
timestamp 1621523292
transform 1 0 37536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_408
timestamp 1621523292
transform 1 0 38640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1621523292
transform 1 0 40480 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_420
timestamp 1621523292
transform 1 0 39744 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_429
timestamp 1621523292
transform 1 0 40572 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_441
timestamp 1621523292
transform 1 0 41676 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_453
timestamp 1621523292
transform 1 0 42780 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_465
timestamp 1621523292
transform 1 0 43884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_477
timestamp 1621523292
transform 1 0 44988 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1621523292
transform 1 0 45724 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_486
timestamp 1621523292
transform 1 0 45816 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_498
timestamp 1621523292
transform 1 0 46920 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1621523292
transform 1 0 49036 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_510
timestamp 1621523292
transform 1 0 48024 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_518
timestamp 1621523292
transform 1 0 48760 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_524
timestamp 1621523292
transform 1 0 49312 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0941_
timestamp 1621523292
transform 1 0 50324 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1083_
timestamp 1621523292
transform 1 0 49680 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1621523292
transform 1 0 50968 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_531
timestamp 1621523292
transform 1 0 49956 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_538
timestamp 1621523292
transform 1 0 50600 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_543
timestamp 1621523292
transform 1 0 51060 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0795_
timestamp 1621523292
transform 1 0 51888 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1621523292
transform 1 0 52532 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_64_551
timestamp 1621523292
transform 1 0 51796 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_555
timestamp 1621523292
transform 1 0 52164 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0767_
timestamp 1621523292
transform 1 0 54372 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_64_575
timestamp 1621523292
transform 1 0 54004 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_586
timestamp 1621523292
transform 1 0 55016 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0599_
timestamp 1621523292
transform 1 0 55384 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1294_
timestamp 1621523292
transform 1 0 57040 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1621523292
transform 1 0 56212 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_593
timestamp 1621523292
transform 1 0 55660 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_600
timestamp 1621523292
transform 1 0 56304 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1621523292
transform -1 0 58880 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_616
timestamp 1621523292
transform 1 0 57776 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_624
timestamp 1621523292
transform 1 0 58512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1621523292
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1621523292
transform 1 0 1380 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_6
timestamp 1621523292
transform 1 0 1656 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_18
timestamp 1621523292
transform 1 0 2760 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_30
timestamp 1621523292
transform 1 0 3864 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_42
timestamp 1621523292
transform 1 0 4968 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1621523292
transform 1 0 6348 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_54
timestamp 1621523292
transform 1 0 6072 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_58
timestamp 1621523292
transform 1 0 6440 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_70
timestamp 1621523292
transform 1 0 7544 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_82
timestamp 1621523292
transform 1 0 8648 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_94
timestamp 1621523292
transform 1 0 9752 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_106
timestamp 1621523292
transform 1 0 10856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1621523292
transform 1 0 11592 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_115
timestamp 1621523292
transform 1 0 11684 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_127
timestamp 1621523292
transform 1 0 12788 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_139
timestamp 1621523292
transform 1 0 13892 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_151
timestamp 1621523292
transform 1 0 14996 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1621523292
transform 1 0 16836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_163
timestamp 1621523292
transform 1 0 16100 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_172
timestamp 1621523292
transform 1 0 16928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1621523292
transform 1 0 18032 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1621523292
transform 1 0 19136 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1621523292
transform 1 0 20240 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1621523292
transform 1 0 22080 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_220
timestamp 1621523292
transform 1 0 21344 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_229
timestamp 1621523292
transform 1 0 22172 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_241
timestamp 1621523292
transform 1 0 23276 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_253
timestamp 1621523292
transform 1 0 24380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_265
timestamp 1621523292
transform 1 0 25484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_277
timestamp 1621523292
transform 1 0 26588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1621523292
transform 1 0 27324 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_286
timestamp 1621523292
transform 1 0 27416 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_298
timestamp 1621523292
transform 1 0 28520 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_310
timestamp 1621523292
transform 1 0 29624 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1621523292
transform 1 0 30728 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1621523292
transform 1 0 32568 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_334
timestamp 1621523292
transform 1 0 31832 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_343
timestamp 1621523292
transform 1 0 32660 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_355
timestamp 1621523292
transform 1 0 33764 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1621523292
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1621523292
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_391
timestamp 1621523292
transform 1 0 37076 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1621523292
transform 1 0 37812 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_400
timestamp 1621523292
transform 1 0 37904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_412
timestamp 1621523292
transform 1 0 39008 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_424
timestamp 1621523292
transform 1 0 40112 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_436
timestamp 1621523292
transform 1 0 41216 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1621523292
transform 1 0 43056 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_448
timestamp 1621523292
transform 1 0 42320 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_457
timestamp 1621523292
transform 1 0 43148 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_469
timestamp 1621523292
transform 1 0 44252 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_481
timestamp 1621523292
transform 1 0 45356 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_493
timestamp 1621523292
transform 1 0 46460 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1621523292
transform 1 0 48300 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1621523292
transform 1 0 47564 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_514
timestamp 1621523292
transform 1 0 48392 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_522
timestamp 1621523292
transform 1 0 49128 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0798_
timestamp 1621523292
transform 1 0 50048 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1188_
timestamp 1621523292
transform 1 0 49404 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1621523292
transform 1 0 50692 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_528
timestamp 1621523292
transform 1 0 49680 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_535
timestamp 1621523292
transform 1 0 50324 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1621523292
transform 1 0 52900 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_555
timestamp 1621523292
transform 1 0 52164 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_566
timestamp 1621523292
transform 1 0 53176 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _0768_
timestamp 1621523292
transform 1 0 54004 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1621523292
transform 1 0 55016 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1621523292
transform 1 0 53544 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_571
timestamp 1621523292
transform 1 0 53636 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_582
timestamp 1621523292
transform 1 0 54648 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1621523292
transform 1 0 56856 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_602
timestamp 1621523292
transform 1 0 56488 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_609
timestamp 1621523292
transform 1 0 57132 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1332_
timestamp 1621523292
transform 1 0 57500 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1621523292
transform -1 0 58880 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1621523292
transform 1 0 58236 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1621523292
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1621523292
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1621523292
transform 1 0 1380 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1621523292
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1621523292
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_6
timestamp 1621523292
transform 1 0 1656 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_18
timestamp 1621523292
transform 1 0 2760 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1621523292
transform 1 0 3772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_27
timestamp 1621523292
transform 1 0 3588 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_30
timestamp 1621523292
transform 1 0 3864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_42
timestamp 1621523292
transform 1 0 4968 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1621523292
transform 1 0 3864 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1621523292
transform 1 0 4968 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1621523292
transform 1 0 6348 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_54
timestamp 1621523292
transform 1 0 6072 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_54
timestamp 1621523292
transform 1 0 6072 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_58
timestamp 1621523292
transform 1 0 6440 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1621523292
transform 1 0 9016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_66
timestamp 1621523292
transform 1 0 7176 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_78
timestamp 1621523292
transform 1 0 8280 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_87
timestamp 1621523292
transform 1 0 9108 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_70
timestamp 1621523292
transform 1 0 7544 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_82
timestamp 1621523292
transform 1 0 8648 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_99
timestamp 1621523292
transform 1 0 10212 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_94
timestamp 1621523292
transform 1 0 9752 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_106
timestamp 1621523292
transform 1 0 10856 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1621523292
transform 1 0 11592 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_111
timestamp 1621523292
transform 1 0 11316 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_123
timestamp 1621523292
transform 1 0 12420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_115
timestamp 1621523292
transform 1 0 11684 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_127
timestamp 1621523292
transform 1 0 12788 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1621523292
transform 1 0 14260 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_135
timestamp 1621523292
transform 1 0 13524 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_144
timestamp 1621523292
transform 1 0 14352 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_139
timestamp 1621523292
transform 1 0 13892 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_151
timestamp 1621523292
transform 1 0 14996 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1621523292
transform 1 0 16836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_156
timestamp 1621523292
transform 1 0 15456 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_168
timestamp 1621523292
transform 1 0 16560 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_163
timestamp 1621523292
transform 1 0 16100 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_172
timestamp 1621523292
transform 1 0 16928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_180
timestamp 1621523292
transform 1 0 17664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_192
timestamp 1621523292
transform 1 0 18768 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1621523292
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1621523292
transform 1 0 19136 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1621523292
transform 1 0 19504 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_201
timestamp 1621523292
transform 1 0 19596 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_213
timestamp 1621523292
transform 1 0 20700 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_208
timestamp 1621523292
transform 1 0 20240 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1621523292
transform 1 0 22080 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_225
timestamp 1621523292
transform 1 0 21804 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_237
timestamp 1621523292
transform 1 0 22908 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_220
timestamp 1621523292
transform 1 0 21344 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_229
timestamp 1621523292
transform 1 0 22172 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1621523292
transform 1 0 24748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_249
timestamp 1621523292
transform 1 0 24012 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_258
timestamp 1621523292
transform 1 0 24840 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_241
timestamp 1621523292
transform 1 0 23276 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_253
timestamp 1621523292
transform 1 0 24380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_270
timestamp 1621523292
transform 1 0 25944 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_282
timestamp 1621523292
transform 1 0 27048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_265
timestamp 1621523292
transform 1 0 25484 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_277
timestamp 1621523292
transform 1 0 26588 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1621523292
transform 1 0 27324 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_294
timestamp 1621523292
transform 1 0 28152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_286
timestamp 1621523292
transform 1 0 27416 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_298
timestamp 1621523292
transform 1 0 28520 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1621523292
transform 1 0 29992 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_306
timestamp 1621523292
transform 1 0 29256 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_315
timestamp 1621523292
transform 1 0 30084 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_327
timestamp 1621523292
transform 1 0 31188 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_310
timestamp 1621523292
transform 1 0 29624 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_322
timestamp 1621523292
transform 1 0 30728 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1621523292
transform 1 0 32568 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_339
timestamp 1621523292
transform 1 0 32292 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_334
timestamp 1621523292
transform 1 0 31832 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_343
timestamp 1621523292
transform 1 0 32660 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1621523292
transform 1 0 35236 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_351
timestamp 1621523292
transform 1 0 33396 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_363
timestamp 1621523292
transform 1 0 34500 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_355
timestamp 1621523292
transform 1 0 33764 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1621523292
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_372
timestamp 1621523292
transform 1 0 35328 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_384
timestamp 1621523292
transform 1 0 36432 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1621523292
transform 1 0 35972 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_391
timestamp 1621523292
transform 1 0 37076 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1621523292
transform 1 0 37812 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_396
timestamp 1621523292
transform 1 0 37536 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_408
timestamp 1621523292
transform 1 0 38640 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_400
timestamp 1621523292
transform 1 0 37904 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_412
timestamp 1621523292
transform 1 0 39008 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1621523292
transform 1 0 40480 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_420
timestamp 1621523292
transform 1 0 39744 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_429
timestamp 1621523292
transform 1 0 40572 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_424
timestamp 1621523292
transform 1 0 40112 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_436
timestamp 1621523292
transform 1 0 41216 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1621523292
transform 1 0 43056 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_441
timestamp 1621523292
transform 1 0 41676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_453
timestamp 1621523292
transform 1 0 42780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_448
timestamp 1621523292
transform 1 0 42320 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_457
timestamp 1621523292
transform 1 0 43148 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_465
timestamp 1621523292
transform 1 0 43884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_477
timestamp 1621523292
transform 1 0 44988 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_469
timestamp 1621523292
transform 1 0 44252 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1621523292
transform 1 0 45724 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_486
timestamp 1621523292
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_498
timestamp 1621523292
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_481
timestamp 1621523292
transform 1 0 45356 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_493
timestamp 1621523292
transform 1 0 46460 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1621523292
transform 1 0 48300 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_510
timestamp 1621523292
transform 1 0 48024 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_522
timestamp 1621523292
transform 1 0 49128 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1621523292
transform 1 0 47564 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_514
timestamp 1621523292
transform 1 0 48392 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0940_
timestamp 1621523292
transform 1 0 51244 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1621523292
transform 1 0 50324 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1621523292
transform 1 0 50968 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1621523292
transform 1 0 50600 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_534
timestamp 1621523292
transform 1 0 50232 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_538
timestamp 1621523292
transform 1 0 50600 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_543
timestamp 1621523292
transform 1 0 51060 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_526
timestamp 1621523292
transform 1 0 49496 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_541
timestamp 1621523292
transform 1 0 50876 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0771_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52716 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0789_
timestamp 1621523292
transform 1 0 52532 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2oi_1  _0797_
timestamp 1621523292
transform 1 0 51428 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0938_
timestamp 1621523292
transform 1 0 51888 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_554
timestamp 1621523292
transform 1 0 52072 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_560
timestamp 1621523292
transform 1 0 52624 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_548
timestamp 1621523292
transform 1 0 51520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_555
timestamp 1621523292
transform 1 0 52164 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_566
timestamp 1621523292
transform 1 0 53176 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_571
timestamp 1621523292
transform 1 0 53636 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_569
timestamp 1621523292
transform 1 0 53452 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1621523292
transform 1 0 53544 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0673_
timestamp 1621523292
transform 1 0 54004 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_578
timestamp 1621523292
transform 1 0 54280 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_585
timestamp 1621523292
transform 1 0 54924 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_577
timestamp 1621523292
transform 1 0 54188 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0671_
timestamp 1621523292
transform 1 0 54832 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0665_
timestamp 1621523292
transform 1 0 54280 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0598_
timestamp 1621523292
transform 1 0 55292 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_599
timestamp 1621523292
transform 1 0 56212 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_591
timestamp 1621523292
transform 1 0 55476 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_600
timestamp 1621523292
transform 1 0 56304 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_598
timestamp 1621523292
transform 1 0 56120 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_592
timestamp 1621523292
transform 1 0 55568 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1621523292
transform 1 0 56212 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_611
timestamp 1621523292
transform 1 0 57316 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_608
timestamp 1621523292
transform 1 0 57040 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 56396 0 1 38624
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0894_
timestamp 1621523292
transform 1 0 57224 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1621523292
transform -1 0 58880 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1621523292
transform -1 0 58880 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output192
timestamp 1621523292
transform 1 0 57868 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output230
timestamp 1621523292
transform 1 0 57868 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_613
timestamp 1621523292
transform 1 0 57500 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_621
timestamp 1621523292
transform 1 0 58236 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1621523292
transform 1 0 58236 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1621523292
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1621523292
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1621523292
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1621523292
transform 1 0 3772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_27
timestamp 1621523292
transform 1 0 3588 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_30
timestamp 1621523292
transform 1 0 3864 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_42
timestamp 1621523292
transform 1 0 4968 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_54
timestamp 1621523292
transform 1 0 6072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1621523292
transform 1 0 9016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_66
timestamp 1621523292
transform 1 0 7176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_78
timestamp 1621523292
transform 1 0 8280 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_87
timestamp 1621523292
transform 1 0 9108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_99
timestamp 1621523292
transform 1 0 10212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_111
timestamp 1621523292
transform 1 0 11316 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_123
timestamp 1621523292
transform 1 0 12420 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1621523292
transform 1 0 14260 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_135
timestamp 1621523292
transform 1 0 13524 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_144
timestamp 1621523292
transform 1 0 14352 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_156
timestamp 1621523292
transform 1 0 15456 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_168
timestamp 1621523292
transform 1 0 16560 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_180
timestamp 1621523292
transform 1 0 17664 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_192
timestamp 1621523292
transform 1 0 18768 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1621523292
transform 1 0 19504 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_201
timestamp 1621523292
transform 1 0 19596 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_213
timestamp 1621523292
transform 1 0 20700 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_225
timestamp 1621523292
transform 1 0 21804 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_237
timestamp 1621523292
transform 1 0 22908 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1621523292
transform 1 0 24748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_249
timestamp 1621523292
transform 1 0 24012 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_258
timestamp 1621523292
transform 1 0 24840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_270
timestamp 1621523292
transform 1 0 25944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_282
timestamp 1621523292
transform 1 0 27048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_294
timestamp 1621523292
transform 1 0 28152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1621523292
transform 1 0 29992 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_306
timestamp 1621523292
transform 1 0 29256 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_315
timestamp 1621523292
transform 1 0 30084 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_327
timestamp 1621523292
transform 1 0 31188 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_339
timestamp 1621523292
transform 1 0 32292 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1621523292
transform 1 0 35236 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_351
timestamp 1621523292
transform 1 0 33396 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_363
timestamp 1621523292
transform 1 0 34500 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1621523292
transform 1 0 35328 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1621523292
transform 1 0 36432 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_396
timestamp 1621523292
transform 1 0 37536 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_408
timestamp 1621523292
transform 1 0 38640 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1621523292
transform 1 0 40480 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_420
timestamp 1621523292
transform 1 0 39744 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_429
timestamp 1621523292
transform 1 0 40572 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_441
timestamp 1621523292
transform 1 0 41676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_453
timestamp 1621523292
transform 1 0 42780 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_465
timestamp 1621523292
transform 1 0 43884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_477
timestamp 1621523292
transform 1 0 44988 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1621523292
transform 1 0 45724 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_486
timestamp 1621523292
transform 1 0 45816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_498
timestamp 1621523292
transform 1 0 46920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_510
timestamp 1621523292
transform 1 0 48024 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_522
timestamp 1621523292
transform 1 0 49128 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1189_
timestamp 1621523292
transform 1 0 50324 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1621523292
transform 1 0 50968 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_534
timestamp 1621523292
transform 1 0 50232 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_538
timestamp 1621523292
transform 1 0 50600 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_543
timestamp 1621523292
transform 1 0 51060 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1621523292
transform 1 0 51612 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0794_
timestamp 1621523292
transform 1 0 52256 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_552
timestamp 1621523292
transform 1 0 51888 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_564
timestamp 1621523292
transform 1 0 52992 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1621523292
transform 1 0 53728 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_588
timestamp 1621523292
transform 1 0 55200 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0596_
timestamp 1621523292
transform 1 0 55568 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1621523292
transform 1 0 56212 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output231
timestamp 1621523292
transform 1 0 56672 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_595
timestamp 1621523292
transform 1 0 55844 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_600
timestamp 1621523292
transform 1 0 56304 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_608
timestamp 1621523292
transform 1 0 57040 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1295_
timestamp 1621523292
transform 1 0 57408 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1621523292
transform -1 0 58880 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_620
timestamp 1621523292
transform 1 0 58144 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_624
timestamp 1621523292
transform 1 0 58512 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1621523292
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1621523292
transform 1 0 1380 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_6
timestamp 1621523292
transform 1 0 1656 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_18
timestamp 1621523292
transform 1 0 2760 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1621523292
transform 1 0 3864 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1621523292
transform 1 0 4968 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1621523292
transform 1 0 6348 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_54
timestamp 1621523292
transform 1 0 6072 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_58
timestamp 1621523292
transform 1 0 6440 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_70
timestamp 1621523292
transform 1 0 7544 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_82
timestamp 1621523292
transform 1 0 8648 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_94
timestamp 1621523292
transform 1 0 9752 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_106
timestamp 1621523292
transform 1 0 10856 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1621523292
transform 1 0 11592 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_115
timestamp 1621523292
transform 1 0 11684 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_127
timestamp 1621523292
transform 1 0 12788 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_139
timestamp 1621523292
transform 1 0 13892 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_151
timestamp 1621523292
transform 1 0 14996 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1621523292
transform 1 0 16836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_163
timestamp 1621523292
transform 1 0 16100 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_172
timestamp 1621523292
transform 1 0 16928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1621523292
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1621523292
transform 1 0 19136 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1621523292
transform 1 0 20240 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1621523292
transform 1 0 22080 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_220
timestamp 1621523292
transform 1 0 21344 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_229
timestamp 1621523292
transform 1 0 22172 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_241
timestamp 1621523292
transform 1 0 23276 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_253
timestamp 1621523292
transform 1 0 24380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_265
timestamp 1621523292
transform 1 0 25484 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_277
timestamp 1621523292
transform 1 0 26588 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1621523292
transform 1 0 27324 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_286
timestamp 1621523292
transform 1 0 27416 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_298
timestamp 1621523292
transform 1 0 28520 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_310
timestamp 1621523292
transform 1 0 29624 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_322
timestamp 1621523292
transform 1 0 30728 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1621523292
transform 1 0 32568 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_334
timestamp 1621523292
transform 1 0 31832 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_343
timestamp 1621523292
transform 1 0 32660 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_355
timestamp 1621523292
transform 1 0 33764 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1621523292
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1621523292
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_391
timestamp 1621523292
transform 1 0 37076 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1621523292
transform 1 0 37812 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_400
timestamp 1621523292
transform 1 0 37904 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_412
timestamp 1621523292
transform 1 0 39008 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_424
timestamp 1621523292
transform 1 0 40112 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_436
timestamp 1621523292
transform 1 0 41216 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1621523292
transform 1 0 43056 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_448
timestamp 1621523292
transform 1 0 42320 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_457
timestamp 1621523292
transform 1 0 43148 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_469
timestamp 1621523292
transform 1 0 44252 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_481
timestamp 1621523292
transform 1 0 45356 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_493
timestamp 1621523292
transform 1 0 46460 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1621523292
transform 1 0 48300 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1621523292
transform 1 0 47564 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_514
timestamp 1621523292
transform 1 0 48392 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0939_
timestamp 1621523292
transform 1 0 50876 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1621523292
transform 1 0 50232 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_526
timestamp 1621523292
transform 1 0 49496 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_537
timestamp 1621523292
transform 1 0 50508 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_544
timestamp 1621523292
transform 1 0 51152 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0672_
timestamp 1621523292
transform 1 0 51520 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0791_
timestamp 1621523292
transform 1 0 52164 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_551
timestamp 1621523292
transform 1 0 51796 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_561
timestamp 1621523292
transform 1 0 52716 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0769_
timestamp 1621523292
transform 1 0 54004 0 1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1621523292
transform 1 0 55292 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1621523292
transform 1 0 53544 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_569
timestamp 1621523292
transform 1 0 53452 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_571
timestamp 1621523292
transform 1 0 53636 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_582
timestamp 1621523292
transform 1 0 54648 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_588
timestamp 1621523292
transform 1 0 55200 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1296_
timestamp 1621523292
transform 1 0 57132 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_605
timestamp 1621523292
transform 1 0 56764 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1621523292
transform -1 0 58880 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1621523292
transform 1 0 57868 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1621523292
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1621523292
transform 1 0 1380 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_6
timestamp 1621523292
transform 1 0 1656 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_18
timestamp 1621523292
transform 1 0 2760 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1621523292
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_26
timestamp 1621523292
transform 1 0 3496 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_30
timestamp 1621523292
transform 1 0 3864 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_42
timestamp 1621523292
transform 1 0 4968 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_54
timestamp 1621523292
transform 1 0 6072 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1621523292
transform 1 0 9016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_66
timestamp 1621523292
transform 1 0 7176 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_78
timestamp 1621523292
transform 1 0 8280 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_87
timestamp 1621523292
transform 1 0 9108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_99
timestamp 1621523292
transform 1 0 10212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_111
timestamp 1621523292
transform 1 0 11316 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_123
timestamp 1621523292
transform 1 0 12420 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1621523292
transform 1 0 14260 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_135
timestamp 1621523292
transform 1 0 13524 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_144
timestamp 1621523292
transform 1 0 14352 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_156
timestamp 1621523292
transform 1 0 15456 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_168
timestamp 1621523292
transform 1 0 16560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_180
timestamp 1621523292
transform 1 0 17664 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_192
timestamp 1621523292
transform 1 0 18768 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1621523292
transform 1 0 19504 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_201
timestamp 1621523292
transform 1 0 19596 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_213
timestamp 1621523292
transform 1 0 20700 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_225
timestamp 1621523292
transform 1 0 21804 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_237
timestamp 1621523292
transform 1 0 22908 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1621523292
transform 1 0 24748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_249
timestamp 1621523292
transform 1 0 24012 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_258
timestamp 1621523292
transform 1 0 24840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_270
timestamp 1621523292
transform 1 0 25944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_282
timestamp 1621523292
transform 1 0 27048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_294
timestamp 1621523292
transform 1 0 28152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1621523292
transform 1 0 29992 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_306
timestamp 1621523292
transform 1 0 29256 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_315
timestamp 1621523292
transform 1 0 30084 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_327
timestamp 1621523292
transform 1 0 31188 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_339
timestamp 1621523292
transform 1 0 32292 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1621523292
transform 1 0 35236 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_351
timestamp 1621523292
transform 1 0 33396 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_363
timestamp 1621523292
transform 1 0 34500 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_372
timestamp 1621523292
transform 1 0 35328 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_384
timestamp 1621523292
transform 1 0 36432 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_396
timestamp 1621523292
transform 1 0 37536 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_408
timestamp 1621523292
transform 1 0 38640 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1621523292
transform 1 0 40480 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_420
timestamp 1621523292
transform 1 0 39744 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_429
timestamp 1621523292
transform 1 0 40572 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_441
timestamp 1621523292
transform 1 0 41676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_453
timestamp 1621523292
transform 1 0 42780 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_465
timestamp 1621523292
transform 1 0 43884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_477
timestamp 1621523292
transform 1 0 44988 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1621523292
transform 1 0 45724 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_486
timestamp 1621523292
transform 1 0 45816 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_498
timestamp 1621523292
transform 1 0 46920 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_510
timestamp 1621523292
transform 1 0 48024 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_522
timestamp 1621523292
transform 1 0 49128 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1621523292
transform 1 0 50324 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1621523292
transform 1 0 50968 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1621523292
transform 1 0 49680 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_531
timestamp 1621523292
transform 1 0 49956 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_538
timestamp 1621523292
transform 1 0 50600 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_543
timestamp 1621523292
transform 1 0 51060 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_2  _0770_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 52992 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2oi_1  _0792_
timestamp 1621523292
transform 1 0 51428 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_70_554
timestamp 1621523292
transform 1 0 52072 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_562
timestamp 1621523292
transform 1 0 52808 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _0597_
timestamp 1621523292
transform 1 0 55108 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0893_
timestamp 1621523292
transform 1 0 54464 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_576
timestamp 1621523292
transform 1 0 54096 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_583
timestamp 1621523292
transform 1 0 54740 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0670_
timestamp 1621523292
transform 1 0 56672 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1621523292
transform 1 0 56212 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_590
timestamp 1621523292
transform 1 0 55384 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_598
timestamp 1621523292
transform 1 0 56120 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_600
timestamp 1621523292
transform 1 0 56304 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_607
timestamp 1621523292
transform 1 0 56948 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _1333_
timestamp 1621523292
transform 1 0 57500 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1621523292
transform -1 0 58880 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1621523292
transform 1 0 58236 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1621523292
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1621523292
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1621523292
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1621523292
transform 1 0 3588 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1621523292
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1621523292
transform 1 0 6348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_51
timestamp 1621523292
transform 1 0 5796 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_58
timestamp 1621523292
transform 1 0 6440 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_70
timestamp 1621523292
transform 1 0 7544 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_82
timestamp 1621523292
transform 1 0 8648 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_94
timestamp 1621523292
transform 1 0 9752 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_106
timestamp 1621523292
transform 1 0 10856 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1621523292
transform 1 0 11592 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_115
timestamp 1621523292
transform 1 0 11684 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_127
timestamp 1621523292
transform 1 0 12788 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_139
timestamp 1621523292
transform 1 0 13892 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_151
timestamp 1621523292
transform 1 0 14996 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1621523292
transform 1 0 16836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_163
timestamp 1621523292
transform 1 0 16100 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_172
timestamp 1621523292
transform 1 0 16928 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1621523292
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_196
timestamp 1621523292
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_208
timestamp 1621523292
transform 1 0 20240 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1621523292
transform 1 0 22080 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_220
timestamp 1621523292
transform 1 0 21344 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_229
timestamp 1621523292
transform 1 0 22172 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_241
timestamp 1621523292
transform 1 0 23276 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_253
timestamp 1621523292
transform 1 0 24380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_265
timestamp 1621523292
transform 1 0 25484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_277
timestamp 1621523292
transform 1 0 26588 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1621523292
transform 1 0 27324 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_286
timestamp 1621523292
transform 1 0 27416 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_298
timestamp 1621523292
transform 1 0 28520 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_310
timestamp 1621523292
transform 1 0 29624 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_322
timestamp 1621523292
transform 1 0 30728 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1621523292
transform 1 0 32568 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_334
timestamp 1621523292
transform 1 0 31832 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_343
timestamp 1621523292
transform 1 0 32660 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_355
timestamp 1621523292
transform 1 0 33764 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1621523292
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1621523292
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_391
timestamp 1621523292
transform 1 0 37076 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1621523292
transform 1 0 37812 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_400
timestamp 1621523292
transform 1 0 37904 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_412
timestamp 1621523292
transform 1 0 39008 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_424
timestamp 1621523292
transform 1 0 40112 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_436
timestamp 1621523292
transform 1 0 41216 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1621523292
transform 1 0 43056 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_448
timestamp 1621523292
transform 1 0 42320 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_457
timestamp 1621523292
transform 1 0 43148 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_469
timestamp 1621523292
transform 1 0 44252 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_481
timestamp 1621523292
transform 1 0 45356 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_493
timestamp 1621523292
transform 1 0 46460 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1621523292
transform 1 0 48300 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1621523292
transform 1 0 47564 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_514
timestamp 1621523292
transform 1 0 48392 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1190_
timestamp 1621523292
transform 1 0 50692 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_526
timestamp 1621523292
transform 1 0 49496 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_538
timestamp 1621523292
transform 1 0 50600 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_542
timestamp 1621523292
transform 1 0 50968 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1621523292
transform 1 0 51336 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_562
timestamp 1621523292
transform 1 0 52808 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1621523292
transform 1 0 54556 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1621523292
transform 1 0 53544 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_571
timestamp 1621523292
transform 1 0 53636 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_579
timestamp 1621523292
transform 1 0 54372 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1621523292
transform 1 0 56396 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output232
timestamp 1621523292
transform 1 0 57132 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_597
timestamp 1621523292
transform 1 0 56028 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_604
timestamp 1621523292
transform 1 0 56672 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_608
timestamp 1621523292
transform 1 0 57040 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1621523292
transform -1 0 58880 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output193
timestamp 1621523292
transform 1 0 57868 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_613
timestamp 1621523292
transform 1 0 57500 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_621
timestamp 1621523292
transform 1 0 58236 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1621523292
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1621523292
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1621523292
transform 1 0 1380 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_6
timestamp 1621523292
transform 1 0 1656 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp 1621523292
transform 1 0 2760 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1621523292
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1621523292
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1621523292
transform 1 0 3772 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_26
timestamp 1621523292
transform 1 0 3496 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_30
timestamp 1621523292
transform 1 0 3864 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_42
timestamp 1621523292
transform 1 0 4968 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1621523292
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1621523292
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1621523292
transform 1 0 6348 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_54
timestamp 1621523292
transform 1 0 6072 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_51
timestamp 1621523292
transform 1 0 5796 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_58
timestamp 1621523292
transform 1 0 6440 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1621523292
transform 1 0 9016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_66
timestamp 1621523292
transform 1 0 7176 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_78
timestamp 1621523292
transform 1 0 8280 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_87
timestamp 1621523292
transform 1 0 9108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_70
timestamp 1621523292
transform 1 0 7544 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_82
timestamp 1621523292
transform 1 0 8648 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_99
timestamp 1621523292
transform 1 0 10212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_94
timestamp 1621523292
transform 1 0 9752 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_106
timestamp 1621523292
transform 1 0 10856 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1621523292
transform 1 0 11592 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_111
timestamp 1621523292
transform 1 0 11316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_123
timestamp 1621523292
transform 1 0 12420 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_115
timestamp 1621523292
transform 1 0 11684 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_127
timestamp 1621523292
transform 1 0 12788 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1621523292
transform 1 0 14260 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_135
timestamp 1621523292
transform 1 0 13524 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_144
timestamp 1621523292
transform 1 0 14352 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_139
timestamp 1621523292
transform 1 0 13892 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_151
timestamp 1621523292
transform 1 0 14996 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1621523292
transform 1 0 16836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_156
timestamp 1621523292
transform 1 0 15456 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_168
timestamp 1621523292
transform 1 0 16560 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_163
timestamp 1621523292
transform 1 0 16100 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_172
timestamp 1621523292
transform 1 0 16928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_180
timestamp 1621523292
transform 1 0 17664 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_192
timestamp 1621523292
transform 1 0 18768 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_184
timestamp 1621523292
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_196
timestamp 1621523292
transform 1 0 19136 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1621523292
transform 1 0 19504 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_201
timestamp 1621523292
transform 1 0 19596 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_213
timestamp 1621523292
transform 1 0 20700 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_208
timestamp 1621523292
transform 1 0 20240 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1621523292
transform 1 0 22080 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_225
timestamp 1621523292
transform 1 0 21804 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_237
timestamp 1621523292
transform 1 0 22908 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_220
timestamp 1621523292
transform 1 0 21344 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_229
timestamp 1621523292
transform 1 0 22172 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1621523292
transform 1 0 24748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_249
timestamp 1621523292
transform 1 0 24012 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_258
timestamp 1621523292
transform 1 0 24840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_241
timestamp 1621523292
transform 1 0 23276 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_253
timestamp 1621523292
transform 1 0 24380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_270
timestamp 1621523292
transform 1 0 25944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_282
timestamp 1621523292
transform 1 0 27048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_265
timestamp 1621523292
transform 1 0 25484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_277
timestamp 1621523292
transform 1 0 26588 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1621523292
transform 1 0 27324 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_294
timestamp 1621523292
transform 1 0 28152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_286
timestamp 1621523292
transform 1 0 27416 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_298
timestamp 1621523292
transform 1 0 28520 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1621523292
transform 1 0 29992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_306
timestamp 1621523292
transform 1 0 29256 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_315
timestamp 1621523292
transform 1 0 30084 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_327
timestamp 1621523292
transform 1 0 31188 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_310
timestamp 1621523292
transform 1 0 29624 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_322
timestamp 1621523292
transform 1 0 30728 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1621523292
transform 1 0 32568 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_339
timestamp 1621523292
transform 1 0 32292 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_334
timestamp 1621523292
transform 1 0 31832 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_343
timestamp 1621523292
transform 1 0 32660 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1621523292
transform 1 0 35236 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_351
timestamp 1621523292
transform 1 0 33396 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_363
timestamp 1621523292
transform 1 0 34500 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_355
timestamp 1621523292
transform 1 0 33764 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1621523292
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_372
timestamp 1621523292
transform 1 0 35328 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_384
timestamp 1621523292
transform 1 0 36432 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1621523292
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_391
timestamp 1621523292
transform 1 0 37076 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1621523292
transform 1 0 37812 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_396
timestamp 1621523292
transform 1 0 37536 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_408
timestamp 1621523292
transform 1 0 38640 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_400
timestamp 1621523292
transform 1 0 37904 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_412
timestamp 1621523292
transform 1 0 39008 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1621523292
transform 1 0 40480 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_420
timestamp 1621523292
transform 1 0 39744 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_429
timestamp 1621523292
transform 1 0 40572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_424
timestamp 1621523292
transform 1 0 40112 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_436
timestamp 1621523292
transform 1 0 41216 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1621523292
transform 1 0 43056 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_441
timestamp 1621523292
transform 1 0 41676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_453
timestamp 1621523292
transform 1 0 42780 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_448
timestamp 1621523292
transform 1 0 42320 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_457
timestamp 1621523292
transform 1 0 43148 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_465
timestamp 1621523292
transform 1 0 43884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_477
timestamp 1621523292
transform 1 0 44988 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_469
timestamp 1621523292
transform 1 0 44252 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1621523292
transform 1 0 45724 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_486
timestamp 1621523292
transform 1 0 45816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_498
timestamp 1621523292
transform 1 0 46920 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_481
timestamp 1621523292
transform 1 0 45356 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_493
timestamp 1621523292
transform 1 0 46460 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1621523292
transform 1 0 48300 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_510
timestamp 1621523292
transform 1 0 48024 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_522
timestamp 1621523292
transform 1 0 49128 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1621523292
transform 1 0 47564 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_73_514
timestamp 1621523292
transform 1 0 48392 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_522
timestamp 1621523292
transform 1 0 49128 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_528
timestamp 1621523292
transform 1 0 49680 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1621523292
transform 1 0 49404 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0780_
timestamp 1621523292
transform 1 0 50048 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_538
timestamp 1621523292
transform 1 0 50600 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_538
timestamp 1621523292
transform 1 0 50600 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_534
timestamp 1621523292
transform 1 0 50232 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1087_
timestamp 1621523292
transform 1 0 50324 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_543
timestamp 1621523292
transform 1 0 51060 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1621523292
transform 1 0 50968 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _0781_
timestamp 1621523292
transform 1 0 50968 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_550
timestamp 1621523292
transform 1 0 51704 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_550
timestamp 1621523292
transform 1 0 51704 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1621523292
transform 1 0 52072 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1621523292
transform 1 0 51428 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_557
timestamp 1621523292
transform 1 0 52348 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_562
timestamp 1621523292
transform 1 0 52808 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_558
timestamp 1621523292
transform 1 0 52440 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0937_
timestamp 1621523292
transform 1 0 52532 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0783_
timestamp 1621523292
transform 1 0 52716 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_564
timestamp 1621523292
transform 1 0 52992 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0669_
timestamp 1621523292
transform 1 0 53176 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0594_
timestamp 1621523292
transform 1 0 54188 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0595_
timestamp 1621523292
transform 1 0 54832 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1621523292
transform 1 0 54004 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1621523292
transform 1 0 53544 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_573
timestamp 1621523292
transform 1 0 53820 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_580
timestamp 1621523292
transform 1 0 54464 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_587
timestamp 1621523292
transform 1 0 55108 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_571
timestamp 1621523292
transform 1 0 53636 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_598
timestamp 1621523292
transform 1 0 56120 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_591
timestamp 1621523292
transform 1 0 55476 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_595
timestamp 1621523292
transform 1 0 55844 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_591
timestamp 1621523292
transform 1 0 55476 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1621523292
transform 1 0 55568 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0593_
timestamp 1621523292
transform 1 0 55844 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_604
timestamp 1621523292
transform 1 0 56672 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_600
timestamp 1621523292
transform 1 0 56304 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1621523292
transform 1 0 56212 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1297_
timestamp 1621523292
transform 1 0 56764 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0889_
timestamp 1621523292
transform 1 0 56856 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_609
timestamp 1621523292
transform 1 0 57132 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1334_
timestamp 1621523292
transform 1 0 57500 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1621523292
transform -1 0 58880 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1621523292
transform -1 0 58880 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output194
timestamp 1621523292
transform 1 0 57868 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1621523292
transform 1 0 58236 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_613
timestamp 1621523292
transform 1 0 57500 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_621
timestamp 1621523292
transform 1 0 58236 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1621523292
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1621523292
transform 1 0 1380 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_6
timestamp 1621523292
transform 1 0 1656 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_18
timestamp 1621523292
transform 1 0 2760 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1621523292
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_26
timestamp 1621523292
transform 1 0 3496 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_30
timestamp 1621523292
transform 1 0 3864 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_42
timestamp 1621523292
transform 1 0 4968 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_54
timestamp 1621523292
transform 1 0 6072 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1621523292
transform 1 0 9016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_66
timestamp 1621523292
transform 1 0 7176 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_78
timestamp 1621523292
transform 1 0 8280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_87
timestamp 1621523292
transform 1 0 9108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_99
timestamp 1621523292
transform 1 0 10212 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_111
timestamp 1621523292
transform 1 0 11316 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_123
timestamp 1621523292
transform 1 0 12420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1621523292
transform 1 0 14260 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_135
timestamp 1621523292
transform 1 0 13524 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_144
timestamp 1621523292
transform 1 0 14352 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_156
timestamp 1621523292
transform 1 0 15456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_168
timestamp 1621523292
transform 1 0 16560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_180
timestamp 1621523292
transform 1 0 17664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_192
timestamp 1621523292
transform 1 0 18768 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1621523292
transform 1 0 19504 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_201
timestamp 1621523292
transform 1 0 19596 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_213
timestamp 1621523292
transform 1 0 20700 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_225
timestamp 1621523292
transform 1 0 21804 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_237
timestamp 1621523292
transform 1 0 22908 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1621523292
transform 1 0 24748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_249
timestamp 1621523292
transform 1 0 24012 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_258
timestamp 1621523292
transform 1 0 24840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_270
timestamp 1621523292
transform 1 0 25944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_282
timestamp 1621523292
transform 1 0 27048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_294
timestamp 1621523292
transform 1 0 28152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1621523292
transform 1 0 29992 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_306
timestamp 1621523292
transform 1 0 29256 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_315
timestamp 1621523292
transform 1 0 30084 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_327
timestamp 1621523292
transform 1 0 31188 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_339
timestamp 1621523292
transform 1 0 32292 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1621523292
transform 1 0 35236 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_351
timestamp 1621523292
transform 1 0 33396 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_363
timestamp 1621523292
transform 1 0 34500 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_372
timestamp 1621523292
transform 1 0 35328 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_384
timestamp 1621523292
transform 1 0 36432 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_396
timestamp 1621523292
transform 1 0 37536 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_408
timestamp 1621523292
transform 1 0 38640 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1621523292
transform 1 0 40480 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_420
timestamp 1621523292
transform 1 0 39744 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_429
timestamp 1621523292
transform 1 0 40572 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_441
timestamp 1621523292
transform 1 0 41676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_453
timestamp 1621523292
transform 1 0 42780 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_465
timestamp 1621523292
transform 1 0 43884 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_477
timestamp 1621523292
transform 1 0 44988 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1621523292
transform 1 0 45724 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_486
timestamp 1621523292
transform 1 0 45816 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_498
timestamp 1621523292
transform 1 0 46920 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1621523292
transform 1 0 48944 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_74_510
timestamp 1621523292
transform 1 0 48024 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_518
timestamp 1621523292
transform 1 0 48760 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1621523292
transform 1 0 50968 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_536
timestamp 1621523292
transform 1 0 50416 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_543
timestamp 1621523292
transform 1 0 51060 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0659_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 51428 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0787_
timestamp 1621523292
transform 1 0 52624 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_551
timestamp 1621523292
transform 1 0 51796 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_559
timestamp 1621523292
transform 1 0 52532 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _0663_
timestamp 1621523292
transform 1 0 54464 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1621523292
transform 1 0 53728 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_568
timestamp 1621523292
transform 1 0 53360 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_575
timestamp 1621523292
transform 1 0 54004 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_579
timestamp 1621523292
transform 1 0 54372 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_587
timestamp 1621523292
transform 1 0 55108 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0592_
timestamp 1621523292
transform 1 0 55476 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1621523292
transform 1 0 56212 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output233
timestamp 1621523292
transform 1 0 56764 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_594
timestamp 1621523292
transform 1 0 55752 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_598
timestamp 1621523292
transform 1 0 56120 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_600
timestamp 1621523292
transform 1 0 56304 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_604
timestamp 1621523292
transform 1 0 56672 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_609
timestamp 1621523292
transform 1 0 57132 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1335_
timestamp 1621523292
transform 1 0 57500 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1621523292
transform -1 0 58880 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_621
timestamp 1621523292
transform 1 0 58236 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1621523292
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1621523292
transform 1 0 1380 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_6
timestamp 1621523292
transform 1 0 1656 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_18
timestamp 1621523292
transform 1 0 2760 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_30
timestamp 1621523292
transform 1 0 3864 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_42
timestamp 1621523292
transform 1 0 4968 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1621523292
transform 1 0 6348 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_54
timestamp 1621523292
transform 1 0 6072 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_58
timestamp 1621523292
transform 1 0 6440 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_70
timestamp 1621523292
transform 1 0 7544 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_82
timestamp 1621523292
transform 1 0 8648 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_94
timestamp 1621523292
transform 1 0 9752 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_106
timestamp 1621523292
transform 1 0 10856 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1621523292
transform 1 0 11592 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_115
timestamp 1621523292
transform 1 0 11684 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_127
timestamp 1621523292
transform 1 0 12788 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_139
timestamp 1621523292
transform 1 0 13892 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_151
timestamp 1621523292
transform 1 0 14996 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1621523292
transform 1 0 16836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_163
timestamp 1621523292
transform 1 0 16100 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_172
timestamp 1621523292
transform 1 0 16928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1621523292
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1621523292
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_208
timestamp 1621523292
transform 1 0 20240 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1621523292
transform 1 0 22080 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_220
timestamp 1621523292
transform 1 0 21344 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_229
timestamp 1621523292
transform 1 0 22172 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_241
timestamp 1621523292
transform 1 0 23276 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_253
timestamp 1621523292
transform 1 0 24380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_265
timestamp 1621523292
transform 1 0 25484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_277
timestamp 1621523292
transform 1 0 26588 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1621523292
transform 1 0 27324 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_286
timestamp 1621523292
transform 1 0 27416 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_298
timestamp 1621523292
transform 1 0 28520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_310
timestamp 1621523292
transform 1 0 29624 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_322
timestamp 1621523292
transform 1 0 30728 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1621523292
transform 1 0 32568 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_334
timestamp 1621523292
transform 1 0 31832 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_343
timestamp 1621523292
transform 1 0 32660 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_355
timestamp 1621523292
transform 1 0 33764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1621523292
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1621523292
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_391
timestamp 1621523292
transform 1 0 37076 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1621523292
transform 1 0 37812 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_400
timestamp 1621523292
transform 1 0 37904 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_412
timestamp 1621523292
transform 1 0 39008 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_424
timestamp 1621523292
transform 1 0 40112 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_436
timestamp 1621523292
transform 1 0 41216 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1621523292
transform 1 0 43056 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_448
timestamp 1621523292
transform 1 0 42320 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_457
timestamp 1621523292
transform 1 0 43148 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_469
timestamp 1621523292
transform 1 0 44252 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_481
timestamp 1621523292
transform 1 0 45356 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_493
timestamp 1621523292
transform 1 0 46460 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1621523292
transform 1 0 48300 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1621523292
transform 1 0 47564 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_514
timestamp 1621523292
transform 1 0 48392 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0656_
timestamp 1621523292
transform 1 0 50416 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1621523292
transform 1 0 51060 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_526
timestamp 1621523292
transform 1 0 49496 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_534
timestamp 1621523292
transform 1 0 50232 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_539
timestamp 1621523292
transform 1 0 50692 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0775_
timestamp 1621523292
transform 1 0 52532 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__conb_1  _1191_
timestamp 1621523292
transform 1 0 51888 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_546
timestamp 1621523292
transform 1 0 51336 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_75_555
timestamp 1621523292
transform 1 0 52164 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_566
timestamp 1621523292
transform 1 0 53176 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0784_
timestamp 1621523292
transform 1 0 54004 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1621523292
transform 1 0 55016 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1621523292
transform 1 0 53544 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_571
timestamp 1621523292
transform 1 0 53636 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_581
timestamp 1621523292
transform 1 0 54556 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_585
timestamp 1621523292
transform 1 0 54924 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0662_
timestamp 1621523292
transform 1 0 56856 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_602
timestamp 1621523292
transform 1 0 56488 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_609
timestamp 1621523292
transform 1 0 57132 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1621523292
transform -1 0 58880 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output195
timestamp 1621523292
transform 1 0 57868 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1621523292
transform 1 0 58236 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1621523292
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1621523292
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1621523292
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1621523292
transform 1 0 3772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_27
timestamp 1621523292
transform 1 0 3588 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_30
timestamp 1621523292
transform 1 0 3864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1621523292
transform 1 0 4968 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1621523292
transform 1 0 6072 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1621523292
transform 1 0 9016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1621523292
transform 1 0 7176 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_78
timestamp 1621523292
transform 1 0 8280 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_87
timestamp 1621523292
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_99
timestamp 1621523292
transform 1 0 10212 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_111
timestamp 1621523292
transform 1 0 11316 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_123
timestamp 1621523292
transform 1 0 12420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1621523292
transform 1 0 14260 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_135
timestamp 1621523292
transform 1 0 13524 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_144
timestamp 1621523292
transform 1 0 14352 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1621523292
transform 1 0 15456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1621523292
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_180
timestamp 1621523292
transform 1 0 17664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_192
timestamp 1621523292
transform 1 0 18768 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1621523292
transform 1 0 19504 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_201
timestamp 1621523292
transform 1 0 19596 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_213
timestamp 1621523292
transform 1 0 20700 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_225
timestamp 1621523292
transform 1 0 21804 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_237
timestamp 1621523292
transform 1 0 22908 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1621523292
transform 1 0 24748 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_249
timestamp 1621523292
transform 1 0 24012 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_258
timestamp 1621523292
transform 1 0 24840 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_270
timestamp 1621523292
transform 1 0 25944 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_282
timestamp 1621523292
transform 1 0 27048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_294
timestamp 1621523292
transform 1 0 28152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1621523292
transform 1 0 29992 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_306
timestamp 1621523292
transform 1 0 29256 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_315
timestamp 1621523292
transform 1 0 30084 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_327
timestamp 1621523292
transform 1 0 31188 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_339
timestamp 1621523292
transform 1 0 32292 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1621523292
transform 1 0 35236 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_351
timestamp 1621523292
transform 1 0 33396 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_363
timestamp 1621523292
transform 1 0 34500 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_372
timestamp 1621523292
transform 1 0 35328 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_384
timestamp 1621523292
transform 1 0 36432 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_396
timestamp 1621523292
transform 1 0 37536 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_408
timestamp 1621523292
transform 1 0 38640 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1621523292
transform 1 0 40480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_420
timestamp 1621523292
transform 1 0 39744 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_429
timestamp 1621523292
transform 1 0 40572 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_441
timestamp 1621523292
transform 1 0 41676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_453
timestamp 1621523292
transform 1 0 42780 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_465
timestamp 1621523292
transform 1 0 43884 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_477
timestamp 1621523292
transform 1 0 44988 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1621523292
transform 1 0 45724 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_486
timestamp 1621523292
transform 1 0 45816 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_498
timestamp 1621523292
transform 1 0 46920 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_510
timestamp 1621523292
transform 1 0 48024 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_522
timestamp 1621523292
transform 1 0 49128 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1621523292
transform 1 0 50324 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1621523292
transform 1 0 50968 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_534
timestamp 1621523292
transform 1 0 50232 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_538
timestamp 1621523292
transform 1 0 50600 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_543
timestamp 1621523292
transform 1 0 51060 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0657_
timestamp 1621523292
transform 1 0 51428 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _0785_
timestamp 1621523292
transform 1 0 52164 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1621523292
transform 1 0 53268 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_550
timestamp 1621523292
transform 1 0 51704 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_554
timestamp 1621523292
transform 1 0 52072 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_562
timestamp 1621523292
transform 1 0 52808 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_566
timestamp 1621523292
transform 1 0 53176 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0591_
timestamp 1621523292
transform 1 0 55016 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0773_
timestamp 1621523292
transform 1 0 53912 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_570
timestamp 1621523292
transform 1 0 53544 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_582
timestamp 1621523292
transform 1 0 54648 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_589
timestamp 1621523292
transform 1 0 55292 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1298_
timestamp 1621523292
transform 1 0 56856 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1621523292
transform 1 0 56212 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_597
timestamp 1621523292
transform 1 0 56028 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_600
timestamp 1621523292
transform 1 0 56304 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0890_
timestamp 1621523292
transform 1 0 57960 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1621523292
transform -1 0 58880 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_614
timestamp 1621523292
transform 1 0 57592 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_621
timestamp 1621523292
transform 1 0 58236 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1621523292
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1621523292
transform 1 0 1380 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_6
timestamp 1621523292
transform 1 0 1656 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_18
timestamp 1621523292
transform 1 0 2760 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_30
timestamp 1621523292
transform 1 0 3864 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1621523292
transform 1 0 4968 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1621523292
transform 1 0 6348 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_54
timestamp 1621523292
transform 1 0 6072 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_58
timestamp 1621523292
transform 1 0 6440 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_70
timestamp 1621523292
transform 1 0 7544 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_82
timestamp 1621523292
transform 1 0 8648 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_94
timestamp 1621523292
transform 1 0 9752 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_106
timestamp 1621523292
transform 1 0 10856 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1621523292
transform 1 0 11592 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_115
timestamp 1621523292
transform 1 0 11684 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_127
timestamp 1621523292
transform 1 0 12788 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_139
timestamp 1621523292
transform 1 0 13892 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_151
timestamp 1621523292
transform 1 0 14996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1621523292
transform 1 0 16836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_163
timestamp 1621523292
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_172
timestamp 1621523292
transform 1 0 16928 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1621523292
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1621523292
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1621523292
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1621523292
transform 1 0 22080 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_220
timestamp 1621523292
transform 1 0 21344 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_229
timestamp 1621523292
transform 1 0 22172 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_241
timestamp 1621523292
transform 1 0 23276 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_253
timestamp 1621523292
transform 1 0 24380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_265
timestamp 1621523292
transform 1 0 25484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_277
timestamp 1621523292
transform 1 0 26588 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1621523292
transform 1 0 27324 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_286
timestamp 1621523292
transform 1 0 27416 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_298
timestamp 1621523292
transform 1 0 28520 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_310
timestamp 1621523292
transform 1 0 29624 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_322
timestamp 1621523292
transform 1 0 30728 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1621523292
transform 1 0 32568 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_334
timestamp 1621523292
transform 1 0 31832 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_343
timestamp 1621523292
transform 1 0 32660 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_355
timestamp 1621523292
transform 1 0 33764 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1621523292
transform 1 0 34868 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_379
timestamp 1621523292
transform 1 0 35972 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_391
timestamp 1621523292
transform 1 0 37076 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1621523292
transform 1 0 37812 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_400
timestamp 1621523292
transform 1 0 37904 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_412
timestamp 1621523292
transform 1 0 39008 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_424
timestamp 1621523292
transform 1 0 40112 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_436
timestamp 1621523292
transform 1 0 41216 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1621523292
transform 1 0 43056 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_448
timestamp 1621523292
transform 1 0 42320 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_457
timestamp 1621523292
transform 1 0 43148 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_469
timestamp 1621523292
transform 1 0 44252 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_481
timestamp 1621523292
transform 1 0 45356 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_493
timestamp 1621523292
transform 1 0 46460 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1621523292
transform 1 0 48300 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1621523292
transform 1 0 47564 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_514
timestamp 1621523292
transform 1 0 48392 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1621523292
transform 1 0 50140 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_77_526
timestamp 1621523292
transform 1 0 49496 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_532
timestamp 1621523292
transform 1 0 50048 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1621523292
transform 1 0 51980 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1089_
timestamp 1621523292
transform 1 0 52900 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_549
timestamp 1621523292
transform 1 0 51612 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_556
timestamp 1621523292
transform 1 0 52256 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_562
timestamp 1621523292
transform 1 0 52808 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_566
timestamp 1621523292
transform 1 0 53176 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1621523292
transform 1 0 54464 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1621523292
transform 1 0 53544 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_571
timestamp 1621523292
transform 1 0 53636 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_579
timestamp 1621523292
transform 1 0 54372 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output234
timestamp 1621523292
transform 1 0 56764 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_596
timestamp 1621523292
transform 1 0 55936 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_604
timestamp 1621523292
transform 1 0 56672 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_609
timestamp 1621523292
transform 1 0 57132 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1336_
timestamp 1621523292
transform 1 0 57500 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1621523292
transform -1 0 58880 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1621523292
transform 1 0 58236 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1621523292
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_3
timestamp 1621523292
transform 1 0 1380 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1621523292
transform 1 0 2484 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1621523292
transform 1 0 3772 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_27
timestamp 1621523292
transform 1 0 3588 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_30
timestamp 1621523292
transform 1 0 3864 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_42
timestamp 1621523292
transform 1 0 4968 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_54
timestamp 1621523292
transform 1 0 6072 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1621523292
transform 1 0 9016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_66
timestamp 1621523292
transform 1 0 7176 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_78
timestamp 1621523292
transform 1 0 8280 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_87
timestamp 1621523292
transform 1 0 9108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_99
timestamp 1621523292
transform 1 0 10212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_111
timestamp 1621523292
transform 1 0 11316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_123
timestamp 1621523292
transform 1 0 12420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1621523292
transform 1 0 14260 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_135
timestamp 1621523292
transform 1 0 13524 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_144
timestamp 1621523292
transform 1 0 14352 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_156
timestamp 1621523292
transform 1 0 15456 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_168
timestamp 1621523292
transform 1 0 16560 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_180
timestamp 1621523292
transform 1 0 17664 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_192
timestamp 1621523292
transform 1 0 18768 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1621523292
transform 1 0 19504 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_201
timestamp 1621523292
transform 1 0 19596 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_213
timestamp 1621523292
transform 1 0 20700 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_225
timestamp 1621523292
transform 1 0 21804 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_237
timestamp 1621523292
transform 1 0 22908 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1621523292
transform 1 0 24748 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_249
timestamp 1621523292
transform 1 0 24012 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_258
timestamp 1621523292
transform 1 0 24840 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_270
timestamp 1621523292
transform 1 0 25944 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_282
timestamp 1621523292
transform 1 0 27048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_294
timestamp 1621523292
transform 1 0 28152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1621523292
transform 1 0 29992 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_306
timestamp 1621523292
transform 1 0 29256 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_315
timestamp 1621523292
transform 1 0 30084 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_327
timestamp 1621523292
transform 1 0 31188 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_339
timestamp 1621523292
transform 1 0 32292 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1621523292
transform 1 0 35236 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_351
timestamp 1621523292
transform 1 0 33396 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_363
timestamp 1621523292
transform 1 0 34500 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_372
timestamp 1621523292
transform 1 0 35328 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_384
timestamp 1621523292
transform 1 0 36432 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_396
timestamp 1621523292
transform 1 0 37536 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_408
timestamp 1621523292
transform 1 0 38640 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1621523292
transform 1 0 40480 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_420
timestamp 1621523292
transform 1 0 39744 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_429
timestamp 1621523292
transform 1 0 40572 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_441
timestamp 1621523292
transform 1 0 41676 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_453
timestamp 1621523292
transform 1 0 42780 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_465
timestamp 1621523292
transform 1 0 43884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1621523292
transform 1 0 44988 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1621523292
transform 1 0 45724 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_486
timestamp 1621523292
transform 1 0 45816 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_498
timestamp 1621523292
transform 1 0 46920 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_510
timestamp 1621523292
transform 1 0 48024 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_522
timestamp 1621523292
transform 1 0 49128 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1621523292
transform 1 0 50968 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_534
timestamp 1621523292
transform 1 0 50232 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_543
timestamp 1621523292
transform 1 0 51060 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1621523292
transform 1 0 51980 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_78_551
timestamp 1621523292
transform 1 0 51796 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0587_
timestamp 1621523292
transform 1 0 54832 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0661_
timestamp 1621523292
transform 1 0 53820 0 -1 45152
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_78_569
timestamp 1621523292
transform 1 0 53452 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_580
timestamp 1621523292
transform 1 0 54464 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_587
timestamp 1621523292
transform 1 0 55108 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0772_
timestamp 1621523292
transform 1 0 55568 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1299_
timestamp 1621523292
transform 1 0 56672 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1621523292
transform 1 0 56212 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_591
timestamp 1621523292
transform 1 0 55476 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_595
timestamp 1621523292
transform 1 0 55844 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_600
timestamp 1621523292
transform 1 0 56304 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1621523292
transform -1 0 58880 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output196
timestamp 1621523292
transform 1 0 57868 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_612
timestamp 1621523292
transform 1 0 57408 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_616
timestamp 1621523292
transform 1 0 57776 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_621
timestamp 1621523292
transform 1 0 58236 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1621523292
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1621523292
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1621523292
transform 1 0 1380 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_6
timestamp 1621523292
transform 1 0 1656 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_18
timestamp 1621523292
transform 1 0 2760 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1621523292
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1621523292
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1621523292
transform 1 0 3772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1621523292
transform 1 0 3864 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1621523292
transform 1 0 4968 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_27
timestamp 1621523292
transform 1 0 3588 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_30
timestamp 1621523292
transform 1 0 3864 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_42
timestamp 1621523292
transform 1 0 4968 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1621523292
transform 1 0 6348 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_54
timestamp 1621523292
transform 1 0 6072 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_58
timestamp 1621523292
transform 1 0 6440 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_54
timestamp 1621523292
transform 1 0 6072 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1621523292
transform 1 0 9016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_70
timestamp 1621523292
transform 1 0 7544 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_82
timestamp 1621523292
transform 1 0 8648 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_66
timestamp 1621523292
transform 1 0 7176 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_78
timestamp 1621523292
transform 1 0 8280 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_87
timestamp 1621523292
transform 1 0 9108 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_94
timestamp 1621523292
transform 1 0 9752 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_106
timestamp 1621523292
transform 1 0 10856 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_99
timestamp 1621523292
transform 1 0 10212 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1621523292
transform 1 0 11592 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_115
timestamp 1621523292
transform 1 0 11684 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_127
timestamp 1621523292
transform 1 0 12788 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_111
timestamp 1621523292
transform 1 0 11316 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1621523292
transform 1 0 12420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1621523292
transform 1 0 14260 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_139
timestamp 1621523292
transform 1 0 13892 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_151
timestamp 1621523292
transform 1 0 14996 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_135
timestamp 1621523292
transform 1 0 13524 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_144
timestamp 1621523292
transform 1 0 14352 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1621523292
transform 1 0 16836 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_163
timestamp 1621523292
transform 1 0 16100 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_172
timestamp 1621523292
transform 1 0 16928 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_156
timestamp 1621523292
transform 1 0 15456 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_168
timestamp 1621523292
transform 1 0 16560 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1621523292
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1621523292
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_180
timestamp 1621523292
transform 1 0 17664 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_192
timestamp 1621523292
transform 1 0 18768 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1621523292
transform 1 0 19504 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1621523292
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_201
timestamp 1621523292
transform 1 0 19596 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_213
timestamp 1621523292
transform 1 0 20700 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1621523292
transform 1 0 22080 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_220
timestamp 1621523292
transform 1 0 21344 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_229
timestamp 1621523292
transform 1 0 22172 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_225
timestamp 1621523292
transform 1 0 21804 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_237
timestamp 1621523292
transform 1 0 22908 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1621523292
transform 1 0 24748 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_241
timestamp 1621523292
transform 1 0 23276 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_253
timestamp 1621523292
transform 1 0 24380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_249
timestamp 1621523292
transform 1 0 24012 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_258
timestamp 1621523292
transform 1 0 24840 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_265
timestamp 1621523292
transform 1 0 25484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_277
timestamp 1621523292
transform 1 0 26588 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_270
timestamp 1621523292
transform 1 0 25944 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_282
timestamp 1621523292
transform 1 0 27048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1621523292
transform 1 0 27324 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_286
timestamp 1621523292
transform 1 0 27416 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_298
timestamp 1621523292
transform 1 0 28520 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_294
timestamp 1621523292
transform 1 0 28152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1621523292
transform 1 0 29992 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_310
timestamp 1621523292
transform 1 0 29624 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_322
timestamp 1621523292
transform 1 0 30728 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_306
timestamp 1621523292
transform 1 0 29256 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_315
timestamp 1621523292
transform 1 0 30084 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_327
timestamp 1621523292
transform 1 0 31188 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1621523292
transform 1 0 32568 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_334
timestamp 1621523292
transform 1 0 31832 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_343
timestamp 1621523292
transform 1 0 32660 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_339
timestamp 1621523292
transform 1 0 32292 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1621523292
transform 1 0 35236 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_355
timestamp 1621523292
transform 1 0 33764 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1621523292
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_351
timestamp 1621523292
transform 1 0 33396 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_363
timestamp 1621523292
transform 1 0 34500 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1621523292
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_391
timestamp 1621523292
transform 1 0 37076 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_372
timestamp 1621523292
transform 1 0 35328 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_384
timestamp 1621523292
transform 1 0 36432 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1621523292
transform 1 0 37812 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_400
timestamp 1621523292
transform 1 0 37904 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_412
timestamp 1621523292
transform 1 0 39008 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_396
timestamp 1621523292
transform 1 0 37536 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_408
timestamp 1621523292
transform 1 0 38640 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1621523292
transform 1 0 40480 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_424
timestamp 1621523292
transform 1 0 40112 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_436
timestamp 1621523292
transform 1 0 41216 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_420
timestamp 1621523292
transform 1 0 39744 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_429
timestamp 1621523292
transform 1 0 40572 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1621523292
transform 1 0 43056 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_448
timestamp 1621523292
transform 1 0 42320 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_457
timestamp 1621523292
transform 1 0 43148 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_441
timestamp 1621523292
transform 1 0 41676 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_453
timestamp 1621523292
transform 1 0 42780 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_469
timestamp 1621523292
transform 1 0 44252 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_465
timestamp 1621523292
transform 1 0 43884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_477
timestamp 1621523292
transform 1 0 44988 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1621523292
transform 1 0 45724 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_481
timestamp 1621523292
transform 1 0 45356 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_493
timestamp 1621523292
transform 1 0 46460 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_486
timestamp 1621523292
transform 1 0 45816 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_498
timestamp 1621523292
transform 1 0 46920 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1621523292
transform 1 0 48300 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1621523292
transform 1 0 47564 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_514
timestamp 1621523292
transform 1 0 48392 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_510
timestamp 1621523292
transform 1 0 48024 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_522
timestamp 1621523292
transform 1 0 49128 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1621523292
transform 1 0 50968 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_526
timestamp 1621523292
transform 1 0 49496 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_538
timestamp 1621523292
transform 1 0 50600 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_534
timestamp 1621523292
transform 1 0 50232 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_543
timestamp 1621523292
transform 1 0 51060 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_550
timestamp 1621523292
transform 1 0 51704 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_562
timestamp 1621523292
transform 1 0 52808 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_555
timestamp 1621523292
transform 1 0 52164 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_567
timestamp 1621523292
transform 1 0 53268 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_574
timestamp 1621523292
transform 1 0 53912 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_571
timestamp 1621523292
transform 1 0 53636 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1621523292
transform 1 0 53636 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1621523292
transform 1 0 53544 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_581
timestamp 1621523292
transform 1 0 54556 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_578
timestamp 1621523292
transform 1 0 54280 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _1192_
timestamp 1621523292
transform 1 0 54280 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0660_
timestamp 1621523292
transform 1 0 54004 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_588
timestamp 1621523292
transform 1 0 55200 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_587
timestamp 1621523292
transform 1 0 55108 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1090_
timestamp 1621523292
transform 1 0 54924 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1621523292
transform 1 0 54832 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_595
timestamp 1621523292
transform 1 0 55844 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_594
timestamp 1621523292
transform 1 0 55752 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0935_
timestamp 1621523292
transform 1 0 55476 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0925_
timestamp 1621523292
transform 1 0 55568 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0891_
timestamp 1621523292
transform 1 0 56120 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_80_600
timestamp 1621523292
transform 1 0 56304 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_601
timestamp 1621523292
transform 1 0 56396 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output235
timestamp 1621523292
transform 1 0 56764 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1621523292
transform 1 0 56212 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_608
timestamp 1621523292
transform 1 0 57040 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_609
timestamp 1621523292
transform 1 0 57132 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0920_
timestamp 1621523292
transform 1 0 57224 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0883_
timestamp 1621523292
transform 1 0 57960 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1337_
timestamp 1621523292
transform 1 0 57500 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1621523292
transform -1 0 58880 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1621523292
transform -1 0 58880 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_621
timestamp 1621523292
transform 1 0 58236 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_614
timestamp 1621523292
transform 1 0 57592 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1621523292
transform 1 0 58236 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1621523292
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1621523292
transform 1 0 1380 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_6
timestamp 1621523292
transform 1 0 1656 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_18
timestamp 1621523292
transform 1 0 2760 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1621523292
transform 1 0 3864 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1621523292
transform 1 0 4968 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1621523292
transform 1 0 6348 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_54
timestamp 1621523292
transform 1 0 6072 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_58
timestamp 1621523292
transform 1 0 6440 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_70
timestamp 1621523292
transform 1 0 7544 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_82
timestamp 1621523292
transform 1 0 8648 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_94
timestamp 1621523292
transform 1 0 9752 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_106
timestamp 1621523292
transform 1 0 10856 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1621523292
transform 1 0 11592 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_115
timestamp 1621523292
transform 1 0 11684 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_127
timestamp 1621523292
transform 1 0 12788 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_139
timestamp 1621523292
transform 1 0 13892 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_151
timestamp 1621523292
transform 1 0 14996 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1621523292
transform 1 0 16836 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_163
timestamp 1621523292
transform 1 0 16100 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_172
timestamp 1621523292
transform 1 0 16928 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1621523292
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1621523292
transform 1 0 19136 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_208
timestamp 1621523292
transform 1 0 20240 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1621523292
transform 1 0 22080 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_220
timestamp 1621523292
transform 1 0 21344 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_229
timestamp 1621523292
transform 1 0 22172 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_241
timestamp 1621523292
transform 1 0 23276 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_253
timestamp 1621523292
transform 1 0 24380 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_265
timestamp 1621523292
transform 1 0 25484 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_277
timestamp 1621523292
transform 1 0 26588 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1621523292
transform 1 0 27324 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_286
timestamp 1621523292
transform 1 0 27416 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_298
timestamp 1621523292
transform 1 0 28520 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_310
timestamp 1621523292
transform 1 0 29624 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_322
timestamp 1621523292
transform 1 0 30728 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1621523292
transform 1 0 32568 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_334
timestamp 1621523292
transform 1 0 31832 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_343
timestamp 1621523292
transform 1 0 32660 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_355
timestamp 1621523292
transform 1 0 33764 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1621523292
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1621523292
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_391
timestamp 1621523292
transform 1 0 37076 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1621523292
transform 1 0 37812 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_400
timestamp 1621523292
transform 1 0 37904 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_412
timestamp 1621523292
transform 1 0 39008 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_424
timestamp 1621523292
transform 1 0 40112 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_436
timestamp 1621523292
transform 1 0 41216 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1621523292
transform 1 0 43056 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_448
timestamp 1621523292
transform 1 0 42320 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_457
timestamp 1621523292
transform 1 0 43148 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_469
timestamp 1621523292
transform 1 0 44252 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_481
timestamp 1621523292
transform 1 0 45356 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_493
timestamp 1621523292
transform 1 0 46460 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1621523292
transform 1 0 48300 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1621523292
transform 1 0 47564 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_514
timestamp 1621523292
transform 1 0 48392 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_526
timestamp 1621523292
transform 1 0 49496 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_538
timestamp 1621523292
transform 1 0 50600 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_550
timestamp 1621523292
transform 1 0 51704 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_562
timestamp 1621523292
transform 1 0 52808 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1163_
timestamp 1621523292
transform 1 0 55016 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1621523292
transform 1 0 53544 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1621523292
transform 1 0 54372 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_571
timestamp 1621523292
transform 1 0 53636 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_582
timestamp 1621523292
transform 1 0 54648 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_589
timestamp 1621523292
transform 1 0 55292 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0934_
timestamp 1621523292
transform 1 0 55660 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1300_
timestamp 1621523292
transform 1 0 56304 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_596
timestamp 1621523292
transform 1 0 55936 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_608
timestamp 1621523292
transform 1 0 57040 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _1307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 57408 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1621523292
transform -1 0 58880 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_621
timestamp 1621523292
transform 1 0 58236 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1621523292
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1621523292
transform 1 0 1380 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_6
timestamp 1621523292
transform 1 0 1656 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_18
timestamp 1621523292
transform 1 0 2760 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1621523292
transform 1 0 3772 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_26
timestamp 1621523292
transform 1 0 3496 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_30
timestamp 1621523292
transform 1 0 3864 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_42
timestamp 1621523292
transform 1 0 4968 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_54
timestamp 1621523292
transform 1 0 6072 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1621523292
transform 1 0 9016 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_66
timestamp 1621523292
transform 1 0 7176 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_78
timestamp 1621523292
transform 1 0 8280 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_87
timestamp 1621523292
transform 1 0 9108 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_99
timestamp 1621523292
transform 1 0 10212 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_111
timestamp 1621523292
transform 1 0 11316 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_123
timestamp 1621523292
transform 1 0 12420 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1621523292
transform 1 0 14260 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_135
timestamp 1621523292
transform 1 0 13524 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_144
timestamp 1621523292
transform 1 0 14352 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_156
timestamp 1621523292
transform 1 0 15456 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_168
timestamp 1621523292
transform 1 0 16560 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_180
timestamp 1621523292
transform 1 0 17664 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_192
timestamp 1621523292
transform 1 0 18768 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1621523292
transform 1 0 19504 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_201
timestamp 1621523292
transform 1 0 19596 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_213
timestamp 1621523292
transform 1 0 20700 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_225
timestamp 1621523292
transform 1 0 21804 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_237
timestamp 1621523292
transform 1 0 22908 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1621523292
transform 1 0 24748 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_249
timestamp 1621523292
transform 1 0 24012 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_258
timestamp 1621523292
transform 1 0 24840 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_270
timestamp 1621523292
transform 1 0 25944 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_282
timestamp 1621523292
transform 1 0 27048 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_294
timestamp 1621523292
transform 1 0 28152 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1621523292
transform 1 0 29992 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_306
timestamp 1621523292
transform 1 0 29256 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_315
timestamp 1621523292
transform 1 0 30084 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_327
timestamp 1621523292
transform 1 0 31188 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_339
timestamp 1621523292
transform 1 0 32292 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1621523292
transform 1 0 35236 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_351
timestamp 1621523292
transform 1 0 33396 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_363
timestamp 1621523292
transform 1 0 34500 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_372
timestamp 1621523292
transform 1 0 35328 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_384
timestamp 1621523292
transform 1 0 36432 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_396
timestamp 1621523292
transform 1 0 37536 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_408
timestamp 1621523292
transform 1 0 38640 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1621523292
transform 1 0 40480 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_420
timestamp 1621523292
transform 1 0 39744 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1621523292
transform 1 0 40572 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_441
timestamp 1621523292
transform 1 0 41676 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_453
timestamp 1621523292
transform 1 0 42780 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_465
timestamp 1621523292
transform 1 0 43884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_477
timestamp 1621523292
transform 1 0 44988 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1621523292
transform 1 0 45724 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_486
timestamp 1621523292
transform 1 0 45816 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_498
timestamp 1621523292
transform 1 0 46920 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_510
timestamp 1621523292
transform 1 0 48024 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_522
timestamp 1621523292
transform 1 0 49128 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1621523292
transform 1 0 50968 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_534
timestamp 1621523292
transform 1 0 50232 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_543
timestamp 1621523292
transform 1 0 51060 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_555
timestamp 1621523292
transform 1 0 52164 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_567
timestamp 1621523292
transform 1 0 53268 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1193_
timestamp 1621523292
transform 1 0 54924 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1621523292
transform 1 0 54280 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_82_575
timestamp 1621523292
transform 1 0 54004 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_581
timestamp 1621523292
transform 1 0 54556 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_588
timestamp 1621523292
transform 1 0 55200 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1621523292
transform 1 0 55568 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1621523292
transform 1 0 56212 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output237
timestamp 1621523292
transform 1 0 57132 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_595
timestamp 1621523292
transform 1 0 55844 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_600
timestamp 1621523292
transform 1 0 56304 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_608
timestamp 1621523292
transform 1 0 57040 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1621523292
transform -1 0 58880 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output197
timestamp 1621523292
transform 1 0 57868 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1621523292
transform 1 0 57500 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1621523292
transform 1 0 58236 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1621523292
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1621523292
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1621523292
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1621523292
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1621523292
transform 1 0 4692 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1621523292
transform 1 0 6348 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_51
timestamp 1621523292
transform 1 0 5796 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_58
timestamp 1621523292
transform 1 0 6440 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_70
timestamp 1621523292
transform 1 0 7544 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_82
timestamp 1621523292
transform 1 0 8648 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_94
timestamp 1621523292
transform 1 0 9752 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_106
timestamp 1621523292
transform 1 0 10856 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1621523292
transform 1 0 11592 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_115
timestamp 1621523292
transform 1 0 11684 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_127
timestamp 1621523292
transform 1 0 12788 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_139
timestamp 1621523292
transform 1 0 13892 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_151
timestamp 1621523292
transform 1 0 14996 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1621523292
transform 1 0 16836 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_163
timestamp 1621523292
transform 1 0 16100 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_172
timestamp 1621523292
transform 1 0 16928 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_184
timestamp 1621523292
transform 1 0 18032 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_196
timestamp 1621523292
transform 1 0 19136 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_208
timestamp 1621523292
transform 1 0 20240 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1621523292
transform 1 0 22080 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_220
timestamp 1621523292
transform 1 0 21344 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_229
timestamp 1621523292
transform 1 0 22172 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_241
timestamp 1621523292
transform 1 0 23276 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_253
timestamp 1621523292
transform 1 0 24380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_265
timestamp 1621523292
transform 1 0 25484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_277
timestamp 1621523292
transform 1 0 26588 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1621523292
transform 1 0 27324 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_286
timestamp 1621523292
transform 1 0 27416 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_298
timestamp 1621523292
transform 1 0 28520 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_310
timestamp 1621523292
transform 1 0 29624 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_322
timestamp 1621523292
transform 1 0 30728 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1621523292
transform 1 0 32568 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_334
timestamp 1621523292
transform 1 0 31832 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_343
timestamp 1621523292
transform 1 0 32660 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_355
timestamp 1621523292
transform 1 0 33764 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_367
timestamp 1621523292
transform 1 0 34868 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_379
timestamp 1621523292
transform 1 0 35972 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_391
timestamp 1621523292
transform 1 0 37076 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1621523292
transform 1 0 37812 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_400
timestamp 1621523292
transform 1 0 37904 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_412
timestamp 1621523292
transform 1 0 39008 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_424
timestamp 1621523292
transform 1 0 40112 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_436
timestamp 1621523292
transform 1 0 41216 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1621523292
transform 1 0 43056 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_448
timestamp 1621523292
transform 1 0 42320 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_457
timestamp 1621523292
transform 1 0 43148 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_469
timestamp 1621523292
transform 1 0 44252 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_481
timestamp 1621523292
transform 1 0 45356 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_493
timestamp 1621523292
transform 1 0 46460 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1621523292
transform 1 0 48300 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_505
timestamp 1621523292
transform 1 0 47564 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_514
timestamp 1621523292
transform 1 0 48392 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_526
timestamp 1621523292
transform 1 0 49496 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_538
timestamp 1621523292
transform 1 0 50600 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_550
timestamp 1621523292
transform 1 0 51704 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_562
timestamp 1621523292
transform 1 0 52808 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1621523292
transform 1 0 53544 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_571
timestamp 1621523292
transform 1 0 53636 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_583
timestamp 1621523292
transform 1 0 54740 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1621523292
transform 1 0 56120 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0933_
timestamp 1621523292
transform 1 0 55476 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output199
timestamp 1621523292
transform 1 0 56764 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_594
timestamp 1621523292
transform 1 0 55752 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_601
timestamp 1621523292
transform 1 0 56396 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_609
timestamp 1621523292
transform 1 0 57132 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1338_
timestamp 1621523292
transform 1 0 57500 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1621523292
transform -1 0 58880 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_621
timestamp 1621523292
transform 1 0 58236 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1621523292
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1621523292
transform 1 0 1380 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_6
timestamp 1621523292
transform 1 0 1656 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1621523292
transform 1 0 2760 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1621523292
transform 1 0 3772 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_26
timestamp 1621523292
transform 1 0 3496 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_30
timestamp 1621523292
transform 1 0 3864 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_42
timestamp 1621523292
transform 1 0 4968 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_54
timestamp 1621523292
transform 1 0 6072 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1621523292
transform 1 0 9016 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_66
timestamp 1621523292
transform 1 0 7176 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_78
timestamp 1621523292
transform 1 0 8280 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_87
timestamp 1621523292
transform 1 0 9108 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_99
timestamp 1621523292
transform 1 0 10212 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_111
timestamp 1621523292
transform 1 0 11316 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_123
timestamp 1621523292
transform 1 0 12420 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1621523292
transform 1 0 14260 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_135
timestamp 1621523292
transform 1 0 13524 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_144
timestamp 1621523292
transform 1 0 14352 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_156
timestamp 1621523292
transform 1 0 15456 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_168
timestamp 1621523292
transform 1 0 16560 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_180
timestamp 1621523292
transform 1 0 17664 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_192
timestamp 1621523292
transform 1 0 18768 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1621523292
transform 1 0 19504 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_201
timestamp 1621523292
transform 1 0 19596 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_213
timestamp 1621523292
transform 1 0 20700 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_225
timestamp 1621523292
transform 1 0 21804 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_237
timestamp 1621523292
transform 1 0 22908 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1621523292
transform 1 0 24748 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_249
timestamp 1621523292
transform 1 0 24012 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_258
timestamp 1621523292
transform 1 0 24840 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_270
timestamp 1621523292
transform 1 0 25944 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_282
timestamp 1621523292
transform 1 0 27048 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_294
timestamp 1621523292
transform 1 0 28152 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1621523292
transform 1 0 29992 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_306
timestamp 1621523292
transform 1 0 29256 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_315
timestamp 1621523292
transform 1 0 30084 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_327
timestamp 1621523292
transform 1 0 31188 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_339
timestamp 1621523292
transform 1 0 32292 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1621523292
transform 1 0 35236 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_351
timestamp 1621523292
transform 1 0 33396 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_363
timestamp 1621523292
transform 1 0 34500 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_372
timestamp 1621523292
transform 1 0 35328 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_384
timestamp 1621523292
transform 1 0 36432 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_396
timestamp 1621523292
transform 1 0 37536 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_408
timestamp 1621523292
transform 1 0 38640 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1621523292
transform 1 0 40480 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_420
timestamp 1621523292
transform 1 0 39744 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_429
timestamp 1621523292
transform 1 0 40572 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_441
timestamp 1621523292
transform 1 0 41676 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_453
timestamp 1621523292
transform 1 0 42780 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_465
timestamp 1621523292
transform 1 0 43884 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_477
timestamp 1621523292
transform 1 0 44988 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1621523292
transform 1 0 45724 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_486
timestamp 1621523292
transform 1 0 45816 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_498
timestamp 1621523292
transform 1 0 46920 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_510
timestamp 1621523292
transform 1 0 48024 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_522
timestamp 1621523292
transform 1 0 49128 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1621523292
transform 1 0 50968 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_534
timestamp 1621523292
transform 1 0 50232 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_543
timestamp 1621523292
transform 1 0 51060 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_555
timestamp 1621523292
transform 1 0 52164 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_567
timestamp 1621523292
transform 1 0 53268 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_579
timestamp 1621523292
transform 1 0 54372 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1194_
timestamp 1621523292
transform 1 0 55568 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1301_
timestamp 1621523292
transform 1 0 57040 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1621523292
transform 1 0 56212 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_591
timestamp 1621523292
transform 1 0 55476 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_595
timestamp 1621523292
transform 1 0 55844 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_600
timestamp 1621523292
transform 1 0 56304 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1621523292
transform -1 0 58880 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_616
timestamp 1621523292
transform 1 0 57776 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_624
timestamp 1621523292
transform 1 0 58512 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1621523292
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1621523292
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1621523292
transform 1 0 1380 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1621523292
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1621523292
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_6
timestamp 1621523292
transform 1 0 1656 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 1621523292
transform 1 0 2760 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1621523292
transform 1 0 3772 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1621523292
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1621523292
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_26
timestamp 1621523292
transform 1 0 3496 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_30
timestamp 1621523292
transform 1 0 3864 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_42
timestamp 1621523292
transform 1 0 4968 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1621523292
transform 1 0 6348 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_51
timestamp 1621523292
transform 1 0 5796 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_58
timestamp 1621523292
transform 1 0 6440 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_54
timestamp 1621523292
transform 1 0 6072 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1621523292
transform 1 0 9016 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_70
timestamp 1621523292
transform 1 0 7544 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_82
timestamp 1621523292
transform 1 0 8648 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_66
timestamp 1621523292
transform 1 0 7176 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_78
timestamp 1621523292
transform 1 0 8280 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_87
timestamp 1621523292
transform 1 0 9108 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_94
timestamp 1621523292
transform 1 0 9752 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_106
timestamp 1621523292
transform 1 0 10856 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_99
timestamp 1621523292
transform 1 0 10212 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1621523292
transform 1 0 11592 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_115
timestamp 1621523292
transform 1 0 11684 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_127
timestamp 1621523292
transform 1 0 12788 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_111
timestamp 1621523292
transform 1 0 11316 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_123
timestamp 1621523292
transform 1 0 12420 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1621523292
transform 1 0 14260 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_139
timestamp 1621523292
transform 1 0 13892 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_151
timestamp 1621523292
transform 1 0 14996 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_135
timestamp 1621523292
transform 1 0 13524 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_144
timestamp 1621523292
transform 1 0 14352 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1621523292
transform 1 0 16836 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_163
timestamp 1621523292
transform 1 0 16100 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_172
timestamp 1621523292
transform 1 0 16928 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_156
timestamp 1621523292
transform 1 0 15456 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_168
timestamp 1621523292
transform 1 0 16560 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_184
timestamp 1621523292
transform 1 0 18032 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_196
timestamp 1621523292
transform 1 0 19136 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_180
timestamp 1621523292
transform 1 0 17664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_192
timestamp 1621523292
transform 1 0 18768 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1621523292
transform 1 0 19504 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_208
timestamp 1621523292
transform 1 0 20240 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_201
timestamp 1621523292
transform 1 0 19596 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_213
timestamp 1621523292
transform 1 0 20700 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1621523292
transform 1 0 22080 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_220
timestamp 1621523292
transform 1 0 21344 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_229
timestamp 1621523292
transform 1 0 22172 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_225
timestamp 1621523292
transform 1 0 21804 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_237
timestamp 1621523292
transform 1 0 22908 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1621523292
transform 1 0 24748 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_241
timestamp 1621523292
transform 1 0 23276 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_253
timestamp 1621523292
transform 1 0 24380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_249
timestamp 1621523292
transform 1 0 24012 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_258
timestamp 1621523292
transform 1 0 24840 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_265
timestamp 1621523292
transform 1 0 25484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_277
timestamp 1621523292
transform 1 0 26588 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_270
timestamp 1621523292
transform 1 0 25944 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_282
timestamp 1621523292
transform 1 0 27048 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1621523292
transform 1 0 27324 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_286
timestamp 1621523292
transform 1 0 27416 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_298
timestamp 1621523292
transform 1 0 28520 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_294
timestamp 1621523292
transform 1 0 28152 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1621523292
transform 1 0 29992 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_310
timestamp 1621523292
transform 1 0 29624 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_322
timestamp 1621523292
transform 1 0 30728 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_306
timestamp 1621523292
transform 1 0 29256 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_315
timestamp 1621523292
transform 1 0 30084 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_327
timestamp 1621523292
transform 1 0 31188 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1621523292
transform 1 0 32568 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_334
timestamp 1621523292
transform 1 0 31832 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_343
timestamp 1621523292
transform 1 0 32660 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_339
timestamp 1621523292
transform 1 0 32292 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1621523292
transform 1 0 35236 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_355
timestamp 1621523292
transform 1 0 33764 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1621523292
transform 1 0 34868 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_351
timestamp 1621523292
transform 1 0 33396 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_363
timestamp 1621523292
transform 1 0 34500 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_379
timestamp 1621523292
transform 1 0 35972 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_391
timestamp 1621523292
transform 1 0 37076 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_372
timestamp 1621523292
transform 1 0 35328 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_384
timestamp 1621523292
transform 1 0 36432 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1621523292
transform 1 0 37812 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_400
timestamp 1621523292
transform 1 0 37904 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_412
timestamp 1621523292
transform 1 0 39008 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_396
timestamp 1621523292
transform 1 0 37536 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_408
timestamp 1621523292
transform 1 0 38640 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1621523292
transform 1 0 40480 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_424
timestamp 1621523292
transform 1 0 40112 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_436
timestamp 1621523292
transform 1 0 41216 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_420
timestamp 1621523292
transform 1 0 39744 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_429
timestamp 1621523292
transform 1 0 40572 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1621523292
transform 1 0 43056 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_448
timestamp 1621523292
transform 1 0 42320 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_457
timestamp 1621523292
transform 1 0 43148 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_441
timestamp 1621523292
transform 1 0 41676 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_453
timestamp 1621523292
transform 1 0 42780 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_469
timestamp 1621523292
transform 1 0 44252 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_465
timestamp 1621523292
transform 1 0 43884 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_477
timestamp 1621523292
transform 1 0 44988 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1621523292
transform 1 0 45724 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_481
timestamp 1621523292
transform 1 0 45356 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_493
timestamp 1621523292
transform 1 0 46460 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_486
timestamp 1621523292
transform 1 0 45816 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_498
timestamp 1621523292
transform 1 0 46920 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1621523292
transform 1 0 48300 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_505
timestamp 1621523292
transform 1 0 47564 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_514
timestamp 1621523292
transform 1 0 48392 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_510
timestamp 1621523292
transform 1 0 48024 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_522
timestamp 1621523292
transform 1 0 49128 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1621523292
transform 1 0 50968 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_526
timestamp 1621523292
transform 1 0 49496 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_538
timestamp 1621523292
transform 1 0 50600 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_534
timestamp 1621523292
transform 1 0 50232 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_543
timestamp 1621523292
transform 1 0 51060 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_550
timestamp 1621523292
transform 1 0 51704 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_562
timestamp 1621523292
transform 1 0 52808 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_555
timestamp 1621523292
transform 1 0 52164 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_567
timestamp 1621523292
transform 1 0 53268 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1621523292
transform 1 0 53544 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_571
timestamp 1621523292
transform 1 0 53636 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_583
timestamp 1621523292
transform 1 0 54740 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_579
timestamp 1621523292
transform 1 0 54372 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_595
timestamp 1621523292
transform 1 0 55844 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_591
timestamp 1621523292
transform 1 0 55476 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_594
timestamp 1621523292
transform 1 0 55752 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1621523292
transform 1 0 55476 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1195_
timestamp 1621523292
transform 1 0 55568 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1157_
timestamp 1621523292
transform 1 0 56120 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_86_600
timestamp 1621523292
transform 1 0 56304 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_601
timestamp 1621523292
transform 1 0 56396 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output238
timestamp 1621523292
transform 1 0 56764 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1621523292
transform 1 0 56212 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_608
timestamp 1621523292
transform 1 0 57040 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_609
timestamp 1621523292
transform 1 0 57132 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1621523292
transform 1 0 57224 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1339_
timestamp 1621523292
transform 1 0 57500 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1621523292
transform -1 0 58880 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1621523292
transform -1 0 58880 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output200
timestamp 1621523292
transform 1 0 57868 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1621523292
transform 1 0 58236 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_613
timestamp 1621523292
transform 1 0 57500 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_621
timestamp 1621523292
transform 1 0 58236 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1621523292
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1621523292
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1621523292
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1621523292
transform 1 0 3588 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1621523292
transform 1 0 4692 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1621523292
transform 1 0 6348 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_51
timestamp 1621523292
transform 1 0 5796 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_58
timestamp 1621523292
transform 1 0 6440 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_70
timestamp 1621523292
transform 1 0 7544 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_82
timestamp 1621523292
transform 1 0 8648 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_94
timestamp 1621523292
transform 1 0 9752 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_106
timestamp 1621523292
transform 1 0 10856 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1621523292
transform 1 0 11592 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_115
timestamp 1621523292
transform 1 0 11684 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_127
timestamp 1621523292
transform 1 0 12788 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_139
timestamp 1621523292
transform 1 0 13892 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_151
timestamp 1621523292
transform 1 0 14996 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1621523292
transform 1 0 16836 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_163
timestamp 1621523292
transform 1 0 16100 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_172
timestamp 1621523292
transform 1 0 16928 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_184
timestamp 1621523292
transform 1 0 18032 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_196
timestamp 1621523292
transform 1 0 19136 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_208
timestamp 1621523292
transform 1 0 20240 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1621523292
transform 1 0 22080 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_220
timestamp 1621523292
transform 1 0 21344 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_229
timestamp 1621523292
transform 1 0 22172 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_241
timestamp 1621523292
transform 1 0 23276 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_253
timestamp 1621523292
transform 1 0 24380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_265
timestamp 1621523292
transform 1 0 25484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_277
timestamp 1621523292
transform 1 0 26588 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1621523292
transform 1 0 27324 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_286
timestamp 1621523292
transform 1 0 27416 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_298
timestamp 1621523292
transform 1 0 28520 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_310
timestamp 1621523292
transform 1 0 29624 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_322
timestamp 1621523292
transform 1 0 30728 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1621523292
transform 1 0 32568 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_334
timestamp 1621523292
transform 1 0 31832 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_343
timestamp 1621523292
transform 1 0 32660 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_355
timestamp 1621523292
transform 1 0 33764 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_367
timestamp 1621523292
transform 1 0 34868 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_379
timestamp 1621523292
transform 1 0 35972 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_391
timestamp 1621523292
transform 1 0 37076 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1621523292
transform 1 0 37812 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_400
timestamp 1621523292
transform 1 0 37904 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_412
timestamp 1621523292
transform 1 0 39008 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_424
timestamp 1621523292
transform 1 0 40112 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_436
timestamp 1621523292
transform 1 0 41216 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1621523292
transform 1 0 43056 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_448
timestamp 1621523292
transform 1 0 42320 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_457
timestamp 1621523292
transform 1 0 43148 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_469
timestamp 1621523292
transform 1 0 44252 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_481
timestamp 1621523292
transform 1 0 45356 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_493
timestamp 1621523292
transform 1 0 46460 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1621523292
transform 1 0 48300 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_505
timestamp 1621523292
transform 1 0 47564 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_514
timestamp 1621523292
transform 1 0 48392 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_526
timestamp 1621523292
transform 1 0 49496 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_538
timestamp 1621523292
transform 1 0 50600 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_550
timestamp 1621523292
transform 1 0 51704 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_562
timestamp 1621523292
transform 1 0 52808 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1621523292
transform 1 0 53544 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1621523292
transform 1 0 55200 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_571
timestamp 1621523292
transform 1 0 53636 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_583
timestamp 1621523292
transform 1 0 54740 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_587
timestamp 1621523292
transform 1 0 55108 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1621523292
transform 1 0 56488 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0931_
timestamp 1621523292
transform 1 0 55844 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1302_
timestamp 1621523292
transform 1 0 57132 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_87_591
timestamp 1621523292
transform 1 0 55476 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_598
timestamp 1621523292
transform 1 0 56120 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_605
timestamp 1621523292
transform 1 0 56764 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1621523292
transform -1 0 58880 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_617
timestamp 1621523292
transform 1 0 57868 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1621523292
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1621523292
transform 1 0 1380 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_6
timestamp 1621523292
transform 1 0 1656 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1621523292
transform 1 0 2760 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1621523292
transform 1 0 3772 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_26
timestamp 1621523292
transform 1 0 3496 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_30
timestamp 1621523292
transform 1 0 3864 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_42
timestamp 1621523292
transform 1 0 4968 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_54
timestamp 1621523292
transform 1 0 6072 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1621523292
transform 1 0 9016 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_66
timestamp 1621523292
transform 1 0 7176 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_78
timestamp 1621523292
transform 1 0 8280 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_87
timestamp 1621523292
transform 1 0 9108 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_99
timestamp 1621523292
transform 1 0 10212 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_111
timestamp 1621523292
transform 1 0 11316 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_123
timestamp 1621523292
transform 1 0 12420 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1621523292
transform 1 0 14260 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_135
timestamp 1621523292
transform 1 0 13524 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_144
timestamp 1621523292
transform 1 0 14352 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_156
timestamp 1621523292
transform 1 0 15456 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_168
timestamp 1621523292
transform 1 0 16560 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_180
timestamp 1621523292
transform 1 0 17664 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_192
timestamp 1621523292
transform 1 0 18768 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1621523292
transform 1 0 19504 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_201
timestamp 1621523292
transform 1 0 19596 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_213
timestamp 1621523292
transform 1 0 20700 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_225
timestamp 1621523292
transform 1 0 21804 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_237
timestamp 1621523292
transform 1 0 22908 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1621523292
transform 1 0 24748 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_249
timestamp 1621523292
transform 1 0 24012 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_258
timestamp 1621523292
transform 1 0 24840 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_270
timestamp 1621523292
transform 1 0 25944 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_282
timestamp 1621523292
transform 1 0 27048 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_294
timestamp 1621523292
transform 1 0 28152 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1621523292
transform 1 0 29992 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_306
timestamp 1621523292
transform 1 0 29256 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_315
timestamp 1621523292
transform 1 0 30084 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_327
timestamp 1621523292
transform 1 0 31188 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_339
timestamp 1621523292
transform 1 0 32292 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1621523292
transform 1 0 35236 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_351
timestamp 1621523292
transform 1 0 33396 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_363
timestamp 1621523292
transform 1 0 34500 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_372
timestamp 1621523292
transform 1 0 35328 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_384
timestamp 1621523292
transform 1 0 36432 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_396
timestamp 1621523292
transform 1 0 37536 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_408
timestamp 1621523292
transform 1 0 38640 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1621523292
transform 1 0 40480 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_420
timestamp 1621523292
transform 1 0 39744 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_429
timestamp 1621523292
transform 1 0 40572 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_441
timestamp 1621523292
transform 1 0 41676 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_453
timestamp 1621523292
transform 1 0 42780 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_465
timestamp 1621523292
transform 1 0 43884 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_477
timestamp 1621523292
transform 1 0 44988 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1621523292
transform 1 0 45724 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_486
timestamp 1621523292
transform 1 0 45816 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_498
timestamp 1621523292
transform 1 0 46920 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_510
timestamp 1621523292
transform 1 0 48024 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_522
timestamp 1621523292
transform 1 0 49128 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1621523292
transform 1 0 50968 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_534
timestamp 1621523292
transform 1 0 50232 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_543
timestamp 1621523292
transform 1 0 51060 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_555
timestamp 1621523292
transform 1 0 52164 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_567
timestamp 1621523292
transform 1 0 53268 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_579
timestamp 1621523292
transform 1 0 54372 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1158_
timestamp 1621523292
transform 1 0 55568 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1621523292
transform 1 0 56212 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output239
timestamp 1621523292
transform 1 0 56764 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_591
timestamp 1621523292
transform 1 0 55476 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_595
timestamp 1621523292
transform 1 0 55844 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_600
timestamp 1621523292
transform 1 0 56304 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_604
timestamp 1621523292
transform 1 0 56672 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_609
timestamp 1621523292
transform 1 0 57132 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1340_
timestamp 1621523292
transform 1 0 57500 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1621523292
transform -1 0 58880 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_621
timestamp 1621523292
transform 1 0 58236 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1621523292
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1621523292
transform 1 0 1380 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_6
timestamp 1621523292
transform 1 0 1656 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_18
timestamp 1621523292
transform 1 0 2760 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_30
timestamp 1621523292
transform 1 0 3864 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_42
timestamp 1621523292
transform 1 0 4968 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1621523292
transform 1 0 6348 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_89_54
timestamp 1621523292
transform 1 0 6072 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_58
timestamp 1621523292
transform 1 0 6440 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_70
timestamp 1621523292
transform 1 0 7544 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_82
timestamp 1621523292
transform 1 0 8648 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_94
timestamp 1621523292
transform 1 0 9752 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_106
timestamp 1621523292
transform 1 0 10856 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1621523292
transform 1 0 11592 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_115
timestamp 1621523292
transform 1 0 11684 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_127
timestamp 1621523292
transform 1 0 12788 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_139
timestamp 1621523292
transform 1 0 13892 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_151
timestamp 1621523292
transform 1 0 14996 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1621523292
transform 1 0 16836 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_163
timestamp 1621523292
transform 1 0 16100 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_172
timestamp 1621523292
transform 1 0 16928 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_184
timestamp 1621523292
transform 1 0 18032 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_196
timestamp 1621523292
transform 1 0 19136 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_208
timestamp 1621523292
transform 1 0 20240 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1621523292
transform 1 0 22080 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_220
timestamp 1621523292
transform 1 0 21344 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_229
timestamp 1621523292
transform 1 0 22172 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_241
timestamp 1621523292
transform 1 0 23276 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_253
timestamp 1621523292
transform 1 0 24380 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_265
timestamp 1621523292
transform 1 0 25484 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_277
timestamp 1621523292
transform 1 0 26588 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1621523292
transform 1 0 27324 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_286
timestamp 1621523292
transform 1 0 27416 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_298
timestamp 1621523292
transform 1 0 28520 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_310
timestamp 1621523292
transform 1 0 29624 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_322
timestamp 1621523292
transform 1 0 30728 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1621523292
transform 1 0 32568 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_334
timestamp 1621523292
transform 1 0 31832 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_343
timestamp 1621523292
transform 1 0 32660 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_355
timestamp 1621523292
transform 1 0 33764 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_367
timestamp 1621523292
transform 1 0 34868 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_379
timestamp 1621523292
transform 1 0 35972 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_391
timestamp 1621523292
transform 1 0 37076 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1621523292
transform 1 0 37812 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_400
timestamp 1621523292
transform 1 0 37904 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_412
timestamp 1621523292
transform 1 0 39008 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_424
timestamp 1621523292
transform 1 0 40112 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_436
timestamp 1621523292
transform 1 0 41216 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1621523292
transform 1 0 43056 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_448
timestamp 1621523292
transform 1 0 42320 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_457
timestamp 1621523292
transform 1 0 43148 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_469
timestamp 1621523292
transform 1 0 44252 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_481
timestamp 1621523292
transform 1 0 45356 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_493
timestamp 1621523292
transform 1 0 46460 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1621523292
transform 1 0 48300 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_505
timestamp 1621523292
transform 1 0 47564 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_514
timestamp 1621523292
transform 1 0 48392 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_526
timestamp 1621523292
transform 1 0 49496 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_538
timestamp 1621523292
transform 1 0 50600 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_550
timestamp 1621523292
transform 1 0 51704 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_562
timestamp 1621523292
transform 1 0 52808 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1621523292
transform 1 0 53544 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_571
timestamp 1621523292
transform 1 0 53636 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_583
timestamp 1621523292
transform 1 0 54740 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _0886_
timestamp 1621523292
transform 1 0 57224 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0930_
timestamp 1621523292
transform 1 0 56580 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1196_
timestamp 1621523292
transform 1 0 55936 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_89_595
timestamp 1621523292
transform 1 0 55844 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_599
timestamp 1621523292
transform 1 0 56212 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_606
timestamp 1621523292
transform 1 0 56856 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1621523292
transform -1 0 58880 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output201
timestamp 1621523292
transform 1 0 57868 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_613
timestamp 1621523292
transform 1 0 57500 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_621
timestamp 1621523292
transform 1 0 58236 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1621523292
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1621523292
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1621523292
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1621523292
transform 1 0 3772 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_27
timestamp 1621523292
transform 1 0 3588 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_90_30
timestamp 1621523292
transform 1 0 3864 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_42
timestamp 1621523292
transform 1 0 4968 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_54
timestamp 1621523292
transform 1 0 6072 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1621523292
transform 1 0 9016 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_66
timestamp 1621523292
transform 1 0 7176 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_78
timestamp 1621523292
transform 1 0 8280 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_87
timestamp 1621523292
transform 1 0 9108 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_99
timestamp 1621523292
transform 1 0 10212 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_111
timestamp 1621523292
transform 1 0 11316 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_123
timestamp 1621523292
transform 1 0 12420 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1621523292
transform 1 0 14260 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_135
timestamp 1621523292
transform 1 0 13524 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_144
timestamp 1621523292
transform 1 0 14352 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_156
timestamp 1621523292
transform 1 0 15456 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_168
timestamp 1621523292
transform 1 0 16560 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_180
timestamp 1621523292
transform 1 0 17664 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_192
timestamp 1621523292
transform 1 0 18768 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1621523292
transform 1 0 19504 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_201
timestamp 1621523292
transform 1 0 19596 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_213
timestamp 1621523292
transform 1 0 20700 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_225
timestamp 1621523292
transform 1 0 21804 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_237
timestamp 1621523292
transform 1 0 22908 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1621523292
transform 1 0 24748 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_249
timestamp 1621523292
transform 1 0 24012 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_258
timestamp 1621523292
transform 1 0 24840 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_270
timestamp 1621523292
transform 1 0 25944 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_282
timestamp 1621523292
transform 1 0 27048 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_294
timestamp 1621523292
transform 1 0 28152 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1621523292
transform 1 0 29992 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_306
timestamp 1621523292
transform 1 0 29256 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_315
timestamp 1621523292
transform 1 0 30084 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_327
timestamp 1621523292
transform 1 0 31188 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_339
timestamp 1621523292
transform 1 0 32292 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1621523292
transform 1 0 35236 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_351
timestamp 1621523292
transform 1 0 33396 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_363
timestamp 1621523292
transform 1 0 34500 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_372
timestamp 1621523292
transform 1 0 35328 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_384
timestamp 1621523292
transform 1 0 36432 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_396
timestamp 1621523292
transform 1 0 37536 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_408
timestamp 1621523292
transform 1 0 38640 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1621523292
transform 1 0 40480 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_420
timestamp 1621523292
transform 1 0 39744 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_429
timestamp 1621523292
transform 1 0 40572 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_441
timestamp 1621523292
transform 1 0 41676 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_453
timestamp 1621523292
transform 1 0 42780 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_465
timestamp 1621523292
transform 1 0 43884 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_477
timestamp 1621523292
transform 1 0 44988 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1621523292
transform 1 0 45724 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_486
timestamp 1621523292
transform 1 0 45816 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_498
timestamp 1621523292
transform 1 0 46920 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_510
timestamp 1621523292
transform 1 0 48024 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_522
timestamp 1621523292
transform 1 0 49128 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1621523292
transform 1 0 50968 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_534
timestamp 1621523292
transform 1 0 50232 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_543
timestamp 1621523292
transform 1 0 51060 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_555
timestamp 1621523292
transform 1 0 52164 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_567
timestamp 1621523292
transform 1 0 53268 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _1197_
timestamp 1621523292
transform 1 0 54924 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_90_579
timestamp 1621523292
transform 1 0 54372 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_588
timestamp 1621523292
transform 1 0 55200 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1159_
timestamp 1621523292
transform 1 0 55568 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1303_
timestamp 1621523292
transform 1 0 57040 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1621523292
transform 1 0 56212 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_595
timestamp 1621523292
transform 1 0 55844 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_600
timestamp 1621523292
transform 1 0 56304 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1621523292
transform -1 0 58880 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_90_616
timestamp 1621523292
transform 1 0 57776 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_624
timestamp 1621523292
transform 1 0 58512 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1621523292
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1621523292
transform 1 0 1380 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_6
timestamp 1621523292
transform 1 0 1656 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_18
timestamp 1621523292
transform 1 0 2760 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_30
timestamp 1621523292
transform 1 0 3864 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_42
timestamp 1621523292
transform 1 0 4968 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1621523292
transform 1 0 6348 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_54
timestamp 1621523292
transform 1 0 6072 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_58
timestamp 1621523292
transform 1 0 6440 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_70
timestamp 1621523292
transform 1 0 7544 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_82
timestamp 1621523292
transform 1 0 8648 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_94
timestamp 1621523292
transform 1 0 9752 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_106
timestamp 1621523292
transform 1 0 10856 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1621523292
transform 1 0 11592 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_115
timestamp 1621523292
transform 1 0 11684 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_127
timestamp 1621523292
transform 1 0 12788 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_139
timestamp 1621523292
transform 1 0 13892 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_151
timestamp 1621523292
transform 1 0 14996 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1621523292
transform 1 0 16836 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_163
timestamp 1621523292
transform 1 0 16100 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_172
timestamp 1621523292
transform 1 0 16928 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_184
timestamp 1621523292
transform 1 0 18032 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_196
timestamp 1621523292
transform 1 0 19136 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_208
timestamp 1621523292
transform 1 0 20240 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1621523292
transform 1 0 22080 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_220
timestamp 1621523292
transform 1 0 21344 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_229
timestamp 1621523292
transform 1 0 22172 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_241
timestamp 1621523292
transform 1 0 23276 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_253
timestamp 1621523292
transform 1 0 24380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_265
timestamp 1621523292
transform 1 0 25484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_277
timestamp 1621523292
transform 1 0 26588 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1621523292
transform 1 0 27324 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_286
timestamp 1621523292
transform 1 0 27416 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_298
timestamp 1621523292
transform 1 0 28520 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_310
timestamp 1621523292
transform 1 0 29624 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_322
timestamp 1621523292
transform 1 0 30728 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1621523292
transform 1 0 32568 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_334
timestamp 1621523292
transform 1 0 31832 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_343
timestamp 1621523292
transform 1 0 32660 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_355
timestamp 1621523292
transform 1 0 33764 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_367
timestamp 1621523292
transform 1 0 34868 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_379
timestamp 1621523292
transform 1 0 35972 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_391
timestamp 1621523292
transform 1 0 37076 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1621523292
transform 1 0 37812 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_400
timestamp 1621523292
transform 1 0 37904 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_412
timestamp 1621523292
transform 1 0 39008 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_424
timestamp 1621523292
transform 1 0 40112 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_436
timestamp 1621523292
transform 1 0 41216 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1621523292
transform 1 0 43056 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_448
timestamp 1621523292
transform 1 0 42320 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_457
timestamp 1621523292
transform 1 0 43148 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_469
timestamp 1621523292
transform 1 0 44252 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_481
timestamp 1621523292
transform 1 0 45356 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_493
timestamp 1621523292
transform 1 0 46460 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1621523292
transform 1 0 48300 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_505
timestamp 1621523292
transform 1 0 47564 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_514
timestamp 1621523292
transform 1 0 48392 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_526
timestamp 1621523292
transform 1 0 49496 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_538
timestamp 1621523292
transform 1 0 50600 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_550
timestamp 1621523292
transform 1 0 51704 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_562
timestamp 1621523292
transform 1 0 52808 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1621523292
transform 1 0 53544 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_571
timestamp 1621523292
transform 1 0 53636 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_583
timestamp 1621523292
transform 1 0 54740 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0885_
timestamp 1621523292
transform 1 0 56120 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1621523292
transform 1 0 55476 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output240
timestamp 1621523292
transform 1 0 56764 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_594
timestamp 1621523292
transform 1 0 55752 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_601
timestamp 1621523292
transform 1 0 56396 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_609
timestamp 1621523292
transform 1 0 57132 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1341_
timestamp 1621523292
transform 1 0 57500 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1621523292
transform -1 0 58880 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_621
timestamp 1621523292
transform 1 0 58236 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1621523292
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1621523292
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1621523292
transform 1 0 1380 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1621523292
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1621523292
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_6
timestamp 1621523292
transform 1 0 1656 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_18
timestamp 1621523292
transform 1 0 2760 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1621523292
transform 1 0 3772 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_27
timestamp 1621523292
transform 1 0 3588 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_30
timestamp 1621523292
transform 1 0 3864 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_42
timestamp 1621523292
transform 1 0 4968 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_30
timestamp 1621523292
transform 1 0 3864 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_42
timestamp 1621523292
transform 1 0 4968 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1621523292
transform 1 0 6348 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_54
timestamp 1621523292
transform 1 0 6072 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_54
timestamp 1621523292
transform 1 0 6072 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_58
timestamp 1621523292
transform 1 0 6440 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1621523292
transform 1 0 9016 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_66
timestamp 1621523292
transform 1 0 7176 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_78
timestamp 1621523292
transform 1 0 8280 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_87
timestamp 1621523292
transform 1 0 9108 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_70
timestamp 1621523292
transform 1 0 7544 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_82
timestamp 1621523292
transform 1 0 8648 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_99
timestamp 1621523292
transform 1 0 10212 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_94
timestamp 1621523292
transform 1 0 9752 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_106
timestamp 1621523292
transform 1 0 10856 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1621523292
transform 1 0 11592 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_111
timestamp 1621523292
transform 1 0 11316 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_123
timestamp 1621523292
transform 1 0 12420 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_115
timestamp 1621523292
transform 1 0 11684 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_127
timestamp 1621523292
transform 1 0 12788 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1621523292
transform 1 0 14260 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_135
timestamp 1621523292
transform 1 0 13524 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_144
timestamp 1621523292
transform 1 0 14352 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_139
timestamp 1621523292
transform 1 0 13892 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_151
timestamp 1621523292
transform 1 0 14996 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1621523292
transform 1 0 16836 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_156
timestamp 1621523292
transform 1 0 15456 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_168
timestamp 1621523292
transform 1 0 16560 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_163
timestamp 1621523292
transform 1 0 16100 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_172
timestamp 1621523292
transform 1 0 16928 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_180
timestamp 1621523292
transform 1 0 17664 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_192
timestamp 1621523292
transform 1 0 18768 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_184
timestamp 1621523292
transform 1 0 18032 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_196
timestamp 1621523292
transform 1 0 19136 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1621523292
transform 1 0 19504 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_201
timestamp 1621523292
transform 1 0 19596 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_213
timestamp 1621523292
transform 1 0 20700 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_208
timestamp 1621523292
transform 1 0 20240 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1621523292
transform 1 0 22080 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_225
timestamp 1621523292
transform 1 0 21804 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_237
timestamp 1621523292
transform 1 0 22908 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_220
timestamp 1621523292
transform 1 0 21344 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_229
timestamp 1621523292
transform 1 0 22172 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1621523292
transform 1 0 24748 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_249
timestamp 1621523292
transform 1 0 24012 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_258
timestamp 1621523292
transform 1 0 24840 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_241
timestamp 1621523292
transform 1 0 23276 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_253
timestamp 1621523292
transform 1 0 24380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_270
timestamp 1621523292
transform 1 0 25944 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_282
timestamp 1621523292
transform 1 0 27048 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_265
timestamp 1621523292
transform 1 0 25484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_277
timestamp 1621523292
transform 1 0 26588 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1621523292
transform 1 0 27324 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_294
timestamp 1621523292
transform 1 0 28152 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_286
timestamp 1621523292
transform 1 0 27416 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_298
timestamp 1621523292
transform 1 0 28520 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1621523292
transform 1 0 29992 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_306
timestamp 1621523292
transform 1 0 29256 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_315
timestamp 1621523292
transform 1 0 30084 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_327
timestamp 1621523292
transform 1 0 31188 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_310
timestamp 1621523292
transform 1 0 29624 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_322
timestamp 1621523292
transform 1 0 30728 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1621523292
transform 1 0 32568 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_339
timestamp 1621523292
transform 1 0 32292 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_334
timestamp 1621523292
transform 1 0 31832 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_343
timestamp 1621523292
transform 1 0 32660 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1621523292
transform 1 0 35236 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_351
timestamp 1621523292
transform 1 0 33396 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_363
timestamp 1621523292
transform 1 0 34500 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_355
timestamp 1621523292
transform 1 0 33764 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_367
timestamp 1621523292
transform 1 0 34868 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_372
timestamp 1621523292
transform 1 0 35328 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_384
timestamp 1621523292
transform 1 0 36432 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_379
timestamp 1621523292
transform 1 0 35972 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_391
timestamp 1621523292
transform 1 0 37076 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1621523292
transform 1 0 37812 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_396
timestamp 1621523292
transform 1 0 37536 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_408
timestamp 1621523292
transform 1 0 38640 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_400
timestamp 1621523292
transform 1 0 37904 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_412
timestamp 1621523292
transform 1 0 39008 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1621523292
transform 1 0 40480 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_420
timestamp 1621523292
transform 1 0 39744 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_429
timestamp 1621523292
transform 1 0 40572 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_424
timestamp 1621523292
transform 1 0 40112 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_436
timestamp 1621523292
transform 1 0 41216 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1621523292
transform 1 0 43056 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_441
timestamp 1621523292
transform 1 0 41676 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_453
timestamp 1621523292
transform 1 0 42780 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_448
timestamp 1621523292
transform 1 0 42320 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_457
timestamp 1621523292
transform 1 0 43148 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_465
timestamp 1621523292
transform 1 0 43884 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_477
timestamp 1621523292
transform 1 0 44988 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_469
timestamp 1621523292
transform 1 0 44252 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1621523292
transform 1 0 45724 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_486
timestamp 1621523292
transform 1 0 45816 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_498
timestamp 1621523292
transform 1 0 46920 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_481
timestamp 1621523292
transform 1 0 45356 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_493
timestamp 1621523292
transform 1 0 46460 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1621523292
transform 1 0 48300 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_510
timestamp 1621523292
transform 1 0 48024 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_522
timestamp 1621523292
transform 1 0 49128 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_505
timestamp 1621523292
transform 1 0 47564 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_514
timestamp 1621523292
transform 1 0 48392 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1621523292
transform 1 0 50968 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_534
timestamp 1621523292
transform 1 0 50232 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_543
timestamp 1621523292
transform 1 0 51060 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_526
timestamp 1621523292
transform 1 0 49496 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_538
timestamp 1621523292
transform 1 0 50600 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_555
timestamp 1621523292
transform 1 0 52164 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_567
timestamp 1621523292
transform 1 0 53268 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_550
timestamp 1621523292
transform 1 0 51704 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_562
timestamp 1621523292
transform 1 0 52808 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1621523292
transform 1 0 53544 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_579
timestamp 1621523292
transform 1 0 54372 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_571
timestamp 1621523292
transform 1 0 53636 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_583
timestamp 1621523292
transform 1 0 54740 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_595
timestamp 1621523292
transform 1 0 55844 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_591
timestamp 1621523292
transform 1 0 55476 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_591
timestamp 1621523292
transform 1 0 55476 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1198_
timestamp 1621523292
transform 1 0 55568 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_602
timestamp 1621523292
transform 1 0 56488 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_92_600
timestamp 1621523292
transform 1 0 56304 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1621523292
transform 1 0 56212 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _1160_
timestamp 1621523292
transform 1 0 56212 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0929_
timestamp 1621523292
transform 1 0 56856 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_609
timestamp 1621523292
transform 1 0 57132 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_92_608
timestamp 1621523292
transform 1 0 57040 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1621523292
transform 1 0 57224 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1342_
timestamp 1621523292
transform 1 0 57500 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1621523292
transform -1 0 58880 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1621523292
transform -1 0 58880 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output202
timestamp 1621523292
transform 1 0 57868 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1621523292
transform 1 0 57500 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1621523292
transform 1 0 58236 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_621
timestamp 1621523292
transform 1 0 58236 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1621523292
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1621523292
transform 1 0 1380 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_6
timestamp 1621523292
transform 1 0 1656 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_18
timestamp 1621523292
transform 1 0 2760 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1621523292
transform 1 0 3772 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_94_26
timestamp 1621523292
transform 1 0 3496 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_30
timestamp 1621523292
transform 1 0 3864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_42
timestamp 1621523292
transform 1 0 4968 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_54
timestamp 1621523292
transform 1 0 6072 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1621523292
transform 1 0 9016 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_66
timestamp 1621523292
transform 1 0 7176 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_78
timestamp 1621523292
transform 1 0 8280 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_87
timestamp 1621523292
transform 1 0 9108 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_99
timestamp 1621523292
transform 1 0 10212 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_111
timestamp 1621523292
transform 1 0 11316 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_123
timestamp 1621523292
transform 1 0 12420 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1621523292
transform 1 0 14260 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_135
timestamp 1621523292
transform 1 0 13524 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_144
timestamp 1621523292
transform 1 0 14352 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_156
timestamp 1621523292
transform 1 0 15456 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_168
timestamp 1621523292
transform 1 0 16560 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_180
timestamp 1621523292
transform 1 0 17664 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_192
timestamp 1621523292
transform 1 0 18768 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1621523292
transform 1 0 19504 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_201
timestamp 1621523292
transform 1 0 19596 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_213
timestamp 1621523292
transform 1 0 20700 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_225
timestamp 1621523292
transform 1 0 21804 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_237
timestamp 1621523292
transform 1 0 22908 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1621523292
transform 1 0 24748 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_249
timestamp 1621523292
transform 1 0 24012 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_258
timestamp 1621523292
transform 1 0 24840 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_270
timestamp 1621523292
transform 1 0 25944 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_282
timestamp 1621523292
transform 1 0 27048 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_294
timestamp 1621523292
transform 1 0 28152 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1621523292
transform 1 0 29992 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_306
timestamp 1621523292
transform 1 0 29256 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_315
timestamp 1621523292
transform 1 0 30084 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_327
timestamp 1621523292
transform 1 0 31188 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_339
timestamp 1621523292
transform 1 0 32292 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1621523292
transform 1 0 35236 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_351
timestamp 1621523292
transform 1 0 33396 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_363
timestamp 1621523292
transform 1 0 34500 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_372
timestamp 1621523292
transform 1 0 35328 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_384
timestamp 1621523292
transform 1 0 36432 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_396
timestamp 1621523292
transform 1 0 37536 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_408
timestamp 1621523292
transform 1 0 38640 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1621523292
transform 1 0 40480 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_420
timestamp 1621523292
transform 1 0 39744 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_429
timestamp 1621523292
transform 1 0 40572 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_441
timestamp 1621523292
transform 1 0 41676 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_453
timestamp 1621523292
transform 1 0 42780 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_465
timestamp 1621523292
transform 1 0 43884 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_477
timestamp 1621523292
transform 1 0 44988 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1621523292
transform 1 0 45724 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_486
timestamp 1621523292
transform 1 0 45816 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_498
timestamp 1621523292
transform 1 0 46920 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_510
timestamp 1621523292
transform 1 0 48024 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_522
timestamp 1621523292
transform 1 0 49128 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1621523292
transform 1 0 50968 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_534
timestamp 1621523292
transform 1 0 50232 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_543
timestamp 1621523292
transform 1 0 51060 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_555
timestamp 1621523292
transform 1 0 52164 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_567
timestamp 1621523292
transform 1 0 53268 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_579
timestamp 1621523292
transform 1 0 54372 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_1  _1304_
timestamp 1621523292
transform 1 0 57040 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1621523292
transform 1 0 56212 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1621523292
transform 1 0 55568 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_94_591
timestamp 1621523292
transform 1 0 55476 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_595
timestamp 1621523292
transform 1 0 55844 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_600
timestamp 1621523292
transform 1 0 56304 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1621523292
transform -1 0 58880 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_94_616
timestamp 1621523292
transform 1 0 57776 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_624
timestamp 1621523292
transform 1 0 58512 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1621523292
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1621523292
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1621523292
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1621523292
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1621523292
transform 1 0 4692 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1621523292
transform 1 0 6348 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_51
timestamp 1621523292
transform 1 0 5796 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_95_58
timestamp 1621523292
transform 1 0 6440 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_70
timestamp 1621523292
transform 1 0 7544 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_82
timestamp 1621523292
transform 1 0 8648 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_94
timestamp 1621523292
transform 1 0 9752 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_106
timestamp 1621523292
transform 1 0 10856 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1621523292
transform 1 0 11592 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_115
timestamp 1621523292
transform 1 0 11684 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_127
timestamp 1621523292
transform 1 0 12788 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_139
timestamp 1621523292
transform 1 0 13892 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_151
timestamp 1621523292
transform 1 0 14996 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1621523292
transform 1 0 16836 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_163
timestamp 1621523292
transform 1 0 16100 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_172
timestamp 1621523292
transform 1 0 16928 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_184
timestamp 1621523292
transform 1 0 18032 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_196
timestamp 1621523292
transform 1 0 19136 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_208
timestamp 1621523292
transform 1 0 20240 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1621523292
transform 1 0 22080 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_220
timestamp 1621523292
transform 1 0 21344 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_229
timestamp 1621523292
transform 1 0 22172 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_241
timestamp 1621523292
transform 1 0 23276 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_253
timestamp 1621523292
transform 1 0 24380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_265
timestamp 1621523292
transform 1 0 25484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_277
timestamp 1621523292
transform 1 0 26588 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1621523292
transform 1 0 27324 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_286
timestamp 1621523292
transform 1 0 27416 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_298
timestamp 1621523292
transform 1 0 28520 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_310
timestamp 1621523292
transform 1 0 29624 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_322
timestamp 1621523292
transform 1 0 30728 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1621523292
transform 1 0 32568 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_334
timestamp 1621523292
transform 1 0 31832 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_343
timestamp 1621523292
transform 1 0 32660 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_355
timestamp 1621523292
transform 1 0 33764 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_367
timestamp 1621523292
transform 1 0 34868 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_379
timestamp 1621523292
transform 1 0 35972 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_391
timestamp 1621523292
transform 1 0 37076 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1621523292
transform 1 0 37812 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_400
timestamp 1621523292
transform 1 0 37904 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_412
timestamp 1621523292
transform 1 0 39008 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_424
timestamp 1621523292
transform 1 0 40112 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_436
timestamp 1621523292
transform 1 0 41216 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1621523292
transform 1 0 43056 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_448
timestamp 1621523292
transform 1 0 42320 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_457
timestamp 1621523292
transform 1 0 43148 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_469
timestamp 1621523292
transform 1 0 44252 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_481
timestamp 1621523292
transform 1 0 45356 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_493
timestamp 1621523292
transform 1 0 46460 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1621523292
transform 1 0 48300 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_505
timestamp 1621523292
transform 1 0 47564 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_514
timestamp 1621523292
transform 1 0 48392 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_526
timestamp 1621523292
transform 1 0 49496 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_538
timestamp 1621523292
transform 1 0 50600 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_550
timestamp 1621523292
transform 1 0 51704 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_562
timestamp 1621523292
transform 1 0 52808 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1621523292
transform 1 0 53544 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_571
timestamp 1621523292
transform 1 0 53636 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_583
timestamp 1621523292
transform 1 0 54740 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0927_
timestamp 1621523292
transform 1 0 56120 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1621523292
transform 1 0 55476 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output241
timestamp 1621523292
transform 1 0 56764 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_594
timestamp 1621523292
transform 1 0 55752 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_601
timestamp 1621523292
transform 1 0 56396 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_609
timestamp 1621523292
transform 1 0 57132 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1305_
timestamp 1621523292
transform 1 0 57500 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1621523292
transform -1 0 58880 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1621523292
transform 1 0 58236 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1621523292
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1621523292
transform 1 0 1380 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_6
timestamp 1621523292
transform 1 0 1656 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_18
timestamp 1621523292
transform 1 0 2760 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1621523292
transform 1 0 3772 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_26
timestamp 1621523292
transform 1 0 3496 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_30
timestamp 1621523292
transform 1 0 3864 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_42
timestamp 1621523292
transform 1 0 4968 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_54
timestamp 1621523292
transform 1 0 6072 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1621523292
transform 1 0 9016 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_66
timestamp 1621523292
transform 1 0 7176 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_78
timestamp 1621523292
transform 1 0 8280 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_87
timestamp 1621523292
transform 1 0 9108 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_99
timestamp 1621523292
transform 1 0 10212 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_111
timestamp 1621523292
transform 1 0 11316 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_123
timestamp 1621523292
transform 1 0 12420 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1621523292
transform 1 0 14260 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_135
timestamp 1621523292
transform 1 0 13524 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_144
timestamp 1621523292
transform 1 0 14352 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_156
timestamp 1621523292
transform 1 0 15456 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_168
timestamp 1621523292
transform 1 0 16560 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_180
timestamp 1621523292
transform 1 0 17664 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_192
timestamp 1621523292
transform 1 0 18768 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1621523292
transform 1 0 19504 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_201
timestamp 1621523292
transform 1 0 19596 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_213
timestamp 1621523292
transform 1 0 20700 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_225
timestamp 1621523292
transform 1 0 21804 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_237
timestamp 1621523292
transform 1 0 22908 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1621523292
transform 1 0 24748 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_249
timestamp 1621523292
transform 1 0 24012 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_258
timestamp 1621523292
transform 1 0 24840 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_270
timestamp 1621523292
transform 1 0 25944 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_282
timestamp 1621523292
transform 1 0 27048 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_294
timestamp 1621523292
transform 1 0 28152 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1621523292
transform 1 0 29992 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_306
timestamp 1621523292
transform 1 0 29256 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_315
timestamp 1621523292
transform 1 0 30084 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_327
timestamp 1621523292
transform 1 0 31188 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_339
timestamp 1621523292
transform 1 0 32292 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1621523292
transform 1 0 35236 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_351
timestamp 1621523292
transform 1 0 33396 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_363
timestamp 1621523292
transform 1 0 34500 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_372
timestamp 1621523292
transform 1 0 35328 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_384
timestamp 1621523292
transform 1 0 36432 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_396
timestamp 1621523292
transform 1 0 37536 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_408
timestamp 1621523292
transform 1 0 38640 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1621523292
transform 1 0 40480 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_420
timestamp 1621523292
transform 1 0 39744 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_429
timestamp 1621523292
transform 1 0 40572 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_441
timestamp 1621523292
transform 1 0 41676 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_453
timestamp 1621523292
transform 1 0 42780 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_465
timestamp 1621523292
transform 1 0 43884 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_477
timestamp 1621523292
transform 1 0 44988 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1621523292
transform 1 0 45724 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_486
timestamp 1621523292
transform 1 0 45816 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_498
timestamp 1621523292
transform 1 0 46920 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_510
timestamp 1621523292
transform 1 0 48024 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_522
timestamp 1621523292
transform 1 0 49128 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1621523292
transform 1 0 50968 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_534
timestamp 1621523292
transform 1 0 50232 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_543
timestamp 1621523292
transform 1 0 51060 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_555
timestamp 1621523292
transform 1 0 52164 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_567
timestamp 1621523292
transform 1 0 53268 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0928_
timestamp 1621523292
transform 1 0 54924 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input161
timestamp 1621523292
transform 1 0 54280 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_96_575
timestamp 1621523292
transform 1 0 54004 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_581
timestamp 1621523292
transform 1 0 54556 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_588
timestamp 1621523292
transform 1 0 55200 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0877_
timestamp 1621523292
transform 1 0 55568 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _1343_
timestamp 1621523292
transform 1 0 56672 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1621523292
transform 1 0 56212 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_595
timestamp 1621523292
transform 1 0 55844 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_600
timestamp 1621523292
transform 1 0 56304 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1621523292
transform -1 0 58880 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output203
timestamp 1621523292
transform 1 0 57868 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_612
timestamp 1621523292
transform 1 0 57408 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_616
timestamp 1621523292
transform 1 0 57776 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_621
timestamp 1621523292
transform 1 0 58236 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1621523292
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1621523292
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1621523292
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1621523292
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1621523292
transform 1 0 4692 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1621523292
transform 1 0 6348 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_51
timestamp 1621523292
transform 1 0 5796 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_58
timestamp 1621523292
transform 1 0 6440 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_70
timestamp 1621523292
transform 1 0 7544 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_82
timestamp 1621523292
transform 1 0 8648 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_94
timestamp 1621523292
transform 1 0 9752 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_106
timestamp 1621523292
transform 1 0 10856 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1621523292
transform 1 0 11592 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_115
timestamp 1621523292
transform 1 0 11684 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_127
timestamp 1621523292
transform 1 0 12788 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_139
timestamp 1621523292
transform 1 0 13892 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_151
timestamp 1621523292
transform 1 0 14996 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1621523292
transform 1 0 16836 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_163
timestamp 1621523292
transform 1 0 16100 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_172
timestamp 1621523292
transform 1 0 16928 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_184
timestamp 1621523292
transform 1 0 18032 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_196
timestamp 1621523292
transform 1 0 19136 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_208
timestamp 1621523292
transform 1 0 20240 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1621523292
transform 1 0 22080 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_220
timestamp 1621523292
transform 1 0 21344 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_229
timestamp 1621523292
transform 1 0 22172 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_241
timestamp 1621523292
transform 1 0 23276 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_253
timestamp 1621523292
transform 1 0 24380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_265
timestamp 1621523292
transform 1 0 25484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_277
timestamp 1621523292
transform 1 0 26588 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1621523292
transform 1 0 27324 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_286
timestamp 1621523292
transform 1 0 27416 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_298
timestamp 1621523292
transform 1 0 28520 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_310
timestamp 1621523292
transform 1 0 29624 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_322
timestamp 1621523292
transform 1 0 30728 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1621523292
transform 1 0 32568 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_334
timestamp 1621523292
transform 1 0 31832 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_343
timestamp 1621523292
transform 1 0 32660 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_355
timestamp 1621523292
transform 1 0 33764 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_367
timestamp 1621523292
transform 1 0 34868 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_379
timestamp 1621523292
transform 1 0 35972 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_391
timestamp 1621523292
transform 1 0 37076 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1621523292
transform 1 0 37812 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_400
timestamp 1621523292
transform 1 0 37904 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_412
timestamp 1621523292
transform 1 0 39008 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_424
timestamp 1621523292
transform 1 0 40112 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_436
timestamp 1621523292
transform 1 0 41216 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1621523292
transform 1 0 43056 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_448
timestamp 1621523292
transform 1 0 42320 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_457
timestamp 1621523292
transform 1 0 43148 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_469
timestamp 1621523292
transform 1 0 44252 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_481
timestamp 1621523292
transform 1 0 45356 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_493
timestamp 1621523292
transform 1 0 46460 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1621523292
transform 1 0 48300 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_505
timestamp 1621523292
transform 1 0 47564 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_514
timestamp 1621523292
transform 1 0 48392 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_526
timestamp 1621523292
transform 1 0 49496 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_538
timestamp 1621523292
transform 1 0 50600 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_550
timestamp 1621523292
transform 1 0 51704 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_562
timestamp 1621523292
transform 1 0 52808 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1162_
timestamp 1621523292
transform 1 0 54832 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1621523292
transform 1 0 53544 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input156
timestamp 1621523292
transform 1 0 54188 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_571
timestamp 1621523292
transform 1 0 53636 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_97_580
timestamp 1621523292
transform 1 0 54464 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_587
timestamp 1621523292
transform 1 0 55108 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1621523292
transform 1 0 56120 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1161_
timestamp 1621523292
transform 1 0 55476 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output242
timestamp 1621523292
transform 1 0 56764 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_594
timestamp 1621523292
transform 1 0 55752 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_601
timestamp 1621523292
transform 1 0 56396 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_609
timestamp 1621523292
transform 1 0 57132 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1306_
timestamp 1621523292
transform 1 0 57500 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1621523292
transform -1 0 58880 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1621523292
transform 1 0 58236 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1621523292
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1621523292
transform 1 0 1380 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_6
timestamp 1621523292
transform 1 0 1656 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_18
timestamp 1621523292
transform 1 0 2760 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1621523292
transform 1 0 3772 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input175
timestamp 1621523292
transform 1 0 4232 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_98_26
timestamp 1621523292
transform 1 0 3496 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_30
timestamp 1621523292
transform 1 0 3864 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_37
timestamp 1621523292
transform 1 0 4508 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_49
timestamp 1621523292
transform 1 0 5612 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_61
timestamp 1621523292
transform 1 0 6716 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1621523292
transform 1 0 9016 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_73
timestamp 1621523292
transform 1 0 7820 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_85
timestamp 1621523292
transform 1 0 8924 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_87
timestamp 1621523292
transform 1 0 9108 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_99
timestamp 1621523292
transform 1 0 10212 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_111
timestamp 1621523292
transform 1 0 11316 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_123
timestamp 1621523292
transform 1 0 12420 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1621523292
transform 1 0 14260 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_135
timestamp 1621523292
transform 1 0 13524 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_144
timestamp 1621523292
transform 1 0 14352 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_156
timestamp 1621523292
transform 1 0 15456 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_168
timestamp 1621523292
transform 1 0 16560 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_180
timestamp 1621523292
transform 1 0 17664 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_192
timestamp 1621523292
transform 1 0 18768 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1621523292
transform 1 0 19504 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_201
timestamp 1621523292
transform 1 0 19596 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_213
timestamp 1621523292
transform 1 0 20700 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_225
timestamp 1621523292
transform 1 0 21804 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_237
timestamp 1621523292
transform 1 0 22908 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1621523292
transform 1 0 24748 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_249
timestamp 1621523292
transform 1 0 24012 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_258
timestamp 1621523292
transform 1 0 24840 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_270
timestamp 1621523292
transform 1 0 25944 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_282
timestamp 1621523292
transform 1 0 27048 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_294
timestamp 1621523292
transform 1 0 28152 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1621523292
transform 1 0 29992 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_306
timestamp 1621523292
transform 1 0 29256 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_315
timestamp 1621523292
transform 1 0 30084 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_327
timestamp 1621523292
transform 1 0 31188 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_339
timestamp 1621523292
transform 1 0 32292 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1621523292
transform 1 0 35236 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_351
timestamp 1621523292
transform 1 0 33396 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_363
timestamp 1621523292
transform 1 0 34500 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_372
timestamp 1621523292
transform 1 0 35328 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_384
timestamp 1621523292
transform 1 0 36432 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_396
timestamp 1621523292
transform 1 0 37536 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_408
timestamp 1621523292
transform 1 0 38640 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1621523292
transform 1 0 40480 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_420
timestamp 1621523292
transform 1 0 39744 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_429
timestamp 1621523292
transform 1 0 40572 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_441
timestamp 1621523292
transform 1 0 41676 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_453
timestamp 1621523292
transform 1 0 42780 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_465
timestamp 1621523292
transform 1 0 43884 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_477
timestamp 1621523292
transform 1 0 44988 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1621523292
transform 1 0 45724 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_486
timestamp 1621523292
transform 1 0 45816 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_498
timestamp 1621523292
transform 1 0 46920 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_510
timestamp 1621523292
transform 1 0 48024 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_522
timestamp 1621523292
transform 1 0 49128 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1621523292
transform 1 0 50968 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_534
timestamp 1621523292
transform 1 0 50232 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_543
timestamp 1621523292
transform 1 0 51060 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1621523292
transform 1 0 52992 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1621523292
transform 1 0 52348 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_555
timestamp 1621523292
transform 1 0 52164 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_560
timestamp 1621523292
transform 1 0 52624 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_567
timestamp 1621523292
transform 1 0 53268 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1199_
timestamp 1621523292
transform 1 0 54924 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1621523292
transform 1 0 54280 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input155
timestamp 1621523292
transform 1 0 53636 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_574
timestamp 1621523292
transform 1 0 53912 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_581
timestamp 1621523292
transform 1 0 54556 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_588
timestamp 1621523292
transform 1 0 55200 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0880_
timestamp 1621523292
transform 1 0 55568 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1621523292
transform 1 0 56212 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output244
timestamp 1621523292
transform 1 0 57132 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_595
timestamp 1621523292
transform 1 0 55844 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_600
timestamp 1621523292
transform 1 0 56304 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_608
timestamp 1621523292
transform 1 0 57040 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1621523292
transform -1 0 58880 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output204
timestamp 1621523292
transform 1 0 57868 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_613
timestamp 1621523292
transform 1 0 57500 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_621
timestamp 1621523292
transform 1 0 58236 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_6
timestamp 1621523292
transform 1 0 1656 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_6
timestamp 1621523292
transform 1 0 1656 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1621523292
transform 1 0 1380 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1621523292
transform 1 0 1380 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1621523292
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1621523292
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_14
timestamp 1621523292
transform 1 0 2392 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_13
timestamp 1621523292
transform 1 0 2300 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input174
timestamp 1621523292
transform 1 0 2024 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1621523292
transform 1 0 2484 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_18
timestamp 1621523292
transform 1 0 2760 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1621523292
transform 1 0 2852 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_30
timestamp 1621523292
transform 1 0 3864 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_25
timestamp 1621523292
transform 1 0 3404 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_22
timestamp 1621523292
transform 1 0 3128 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1621523292
transform 1 0 3772 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1205_
timestamp 1621523292
transform 1 0 3496 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _1092_
timestamp 1621523292
transform 1 0 3128 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_36
timestamp 1621523292
transform 1 0 4416 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_41
timestamp 1621523292
transform 1 0 4876 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_34
timestamp 1621523292
transform 1 0 4232 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1048_
timestamp 1621523292
transform 1 0 4600 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4508 0 -1 57120
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _1202_
timestamp 1621523292
transform 1 0 5244 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1621523292
transform 1 0 6348 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_48
timestamp 1621523292
transform 1 0 5520 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_56
timestamp 1621523292
transform 1 0 6256 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_58
timestamp 1621523292
transform 1 0 6440 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_58
timestamp 1621523292
transform 1 0 6440 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1621523292
transform 1 0 9016 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_70
timestamp 1621523292
transform 1 0 7544 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_82
timestamp 1621523292
transform 1 0 8648 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_70
timestamp 1621523292
transform 1 0 7544 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_82
timestamp 1621523292
transform 1 0 8648 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_87
timestamp 1621523292
transform 1 0 9108 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_94
timestamp 1621523292
transform 1 0 9752 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_106
timestamp 1621523292
transform 1 0 10856 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_99
timestamp 1621523292
transform 1 0 10212 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1621523292
transform 1 0 11592 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_115
timestamp 1621523292
transform 1 0 11684 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_127
timestamp 1621523292
transform 1 0 12788 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_111
timestamp 1621523292
transform 1 0 11316 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_123
timestamp 1621523292
transform 1 0 12420 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1621523292
transform 1 0 14260 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_139
timestamp 1621523292
transform 1 0 13892 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_151
timestamp 1621523292
transform 1 0 14996 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_135
timestamp 1621523292
transform 1 0 13524 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_144
timestamp 1621523292
transform 1 0 14352 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1621523292
transform 1 0 16836 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input136
timestamp 1621523292
transform 1 0 16100 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_163
timestamp 1621523292
transform 1 0 16100 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_172
timestamp 1621523292
transform 1 0 16928 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_156
timestamp 1621523292
transform 1 0 15456 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_162
timestamp 1621523292
transform 1 0 16008 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_166
timestamp 1621523292
transform 1 0 16376 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_184
timestamp 1621523292
transform 1 0 18032 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_196
timestamp 1621523292
transform 1 0 19136 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_178
timestamp 1621523292
transform 1 0 17480 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_190
timestamp 1621523292
transform 1 0 18584 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1621523292
transform 1 0 19504 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_208
timestamp 1621523292
transform 1 0 20240 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_198
timestamp 1621523292
transform 1 0 19320 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_201
timestamp 1621523292
transform 1 0 19596 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_213
timestamp 1621523292
transform 1 0 20700 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1621523292
transform 1 0 22080 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_220
timestamp 1621523292
transform 1 0 21344 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_229
timestamp 1621523292
transform 1 0 22172 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_225
timestamp 1621523292
transform 1 0 21804 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_237
timestamp 1621523292
transform 1 0 22908 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1621523292
transform 1 0 24748 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_241
timestamp 1621523292
transform 1 0 23276 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_253
timestamp 1621523292
transform 1 0 24380 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_249
timestamp 1621523292
transform 1 0 24012 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_258
timestamp 1621523292
transform 1 0 24840 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input119
timestamp 1621523292
transform 1 0 26404 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_265
timestamp 1621523292
transform 1 0 25484 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_277
timestamp 1621523292
transform 1 0 26588 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_270
timestamp 1621523292
transform 1 0 25944 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_274
timestamp 1621523292
transform 1 0 26312 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_278
timestamp 1621523292
transform 1 0 26680 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1621523292
transform 1 0 27324 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_286
timestamp 1621523292
transform 1 0 27416 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_298
timestamp 1621523292
transform 1 0 28520 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_290
timestamp 1621523292
transform 1 0 27784 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_302
timestamp 1621523292
transform 1 0 28888 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1621523292
transform 1 0 29992 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_310
timestamp 1621523292
transform 1 0 29624 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_322
timestamp 1621523292
transform 1 0 30728 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_315
timestamp 1621523292
transform 1 0 30084 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_327
timestamp 1621523292
transform 1 0 31188 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1621523292
transform 1 0 32568 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_334
timestamp 1621523292
transform 1 0 31832 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_343
timestamp 1621523292
transform 1 0 32660 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_339
timestamp 1621523292
transform 1 0 32292 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1621523292
transform 1 0 35236 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1621523292
transform 1 0 34224 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_355
timestamp 1621523292
transform 1 0 33764 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1621523292
transform 1 0 34868 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_351
timestamp 1621523292
transform 1 0 33396 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_359
timestamp 1621523292
transform 1 0 34132 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_363
timestamp 1621523292
transform 1 0 34500 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1621523292
transform 1 0 35972 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_391
timestamp 1621523292
transform 1 0 37076 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_372
timestamp 1621523292
transform 1 0 35328 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_384
timestamp 1621523292
transform 1 0 36432 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1621523292
transform 1 0 37812 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_400
timestamp 1621523292
transform 1 0 37904 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_412
timestamp 1621523292
transform 1 0 39008 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_396
timestamp 1621523292
transform 1 0 37536 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_408
timestamp 1621523292
transform 1 0 38640 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1621523292
transform 1 0 40480 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1621523292
transform 1 0 39744 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1621523292
transform 1 0 40940 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_424
timestamp 1621523292
transform 1 0 40112 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_436
timestamp 1621523292
transform 1 0 41216 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_423
timestamp 1621523292
transform 1 0 40020 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_427
timestamp 1621523292
transform 1 0 40388 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_429
timestamp 1621523292
transform 1 0 40572 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_436
timestamp 1621523292
transform 1 0 41216 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1621523292
transform 1 0 43056 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1621523292
transform 1 0 41584 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_448
timestamp 1621523292
transform 1 0 42320 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_457
timestamp 1621523292
transform 1 0 43148 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_443
timestamp 1621523292
transform 1 0 41860 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_455
timestamp 1621523292
transform 1 0 42964 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_469
timestamp 1621523292
transform 1 0 44252 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_467
timestamp 1621523292
transform 1 0 44068 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_479
timestamp 1621523292
transform 1 0 45172 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1621523292
transform 1 0 45724 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_481
timestamp 1621523292
transform 1 0 45356 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_493
timestamp 1621523292
transform 1 0 46460 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_486
timestamp 1621523292
transform 1 0 45816 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_498
timestamp 1621523292
transform 1 0 46920 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1621523292
transform 1 0 48300 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_505
timestamp 1621523292
transform 1 0 47564 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_514
timestamp 1621523292
transform 1 0 48392 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_510
timestamp 1621523292
transform 1 0 48024 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_522
timestamp 1621523292
transform 1 0 49128 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1621523292
transform 1 0 50968 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_526
timestamp 1621523292
transform 1 0 49496 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_538
timestamp 1621523292
transform 1 0 50600 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_534
timestamp 1621523292
transform 1 0 50232 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_543
timestamp 1621523292
transform 1 0 51060 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_550
timestamp 1621523292
transform 1 0 51704 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_552
timestamp 1621523292
transform 1 0 51888 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_546
timestamp 1621523292
transform 1 0 51336 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1621523292
transform 1 0 51612 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1621523292
transform 1 0 51428 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_557
timestamp 1621523292
transform 1 0 52348 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_559
timestamp 1621523292
transform 1 0 52532 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1621523292
transform 1 0 52256 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1621523292
transform 1 0 52072 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_564
timestamp 1621523292
transform 1 0 52992 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_566
timestamp 1621523292
transform 1 0 53176 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input154
timestamp 1621523292
transform 1 0 52900 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input153
timestamp 1621523292
transform 1 0 52716 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_574
timestamp 1621523292
transform 1 0 53912 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_570
timestamp 1621523292
transform 1 0 53544 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_571
timestamp 1621523292
transform 1 0 53636 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1621523292
transform 1 0 53636 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1621523292
transform 1 0 53544 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_581
timestamp 1621523292
transform 1 0 54556 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_580
timestamp 1621523292
transform 1 0 54464 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1204_
timestamp 1621523292
transform 1 0 54188 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1203_
timestamp 1621523292
transform 1 0 54280 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_588
timestamp 1621523292
transform 1 0 55200 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_587
timestamp 1621523292
transform 1 0 55108 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1201_
timestamp 1621523292
transform 1 0 54924 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1200_
timestamp 1621523292
transform 1 0 54832 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_595
timestamp 1621523292
transform 1 0 55844 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_594
timestamp 1621523292
transform 1 0 55752 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1347_
timestamp 1621523292
transform 1 0 56120 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _0879_
timestamp 1621523292
transform 1 0 55568 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1621523292
transform 1 0 55476 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_604
timestamp 1621523292
transform 1 0 56672 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_600
timestamp 1621523292
transform 1 0 56304 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_606
timestamp 1621523292
transform 1 0 56856 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output243
timestamp 1621523292
transform 1 0 56764 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1621523292
transform 1 0 56212 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_609
timestamp 1621523292
transform 1 0 57132 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _1344_
timestamp 1621523292
transform 1 0 57500 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _1345_
timestamp 1621523292
transform 1 0 57500 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1621523292
transform -1 0 58880 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1621523292
transform -1 0 58880 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_99_612
timestamp 1621523292
transform 1 0 57408 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_621
timestamp 1621523292
transform 1 0 58236 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1621523292
transform 1 0 58236 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1621523292
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1621523292
transform 1 0 1380 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1621523292
transform 1 0 2024 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1621523292
transform 1 0 2668 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_6
timestamp 1621523292
transform 1 0 1656 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_13
timestamp 1621523292
transform 1 0 2300 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_20
timestamp 1621523292
transform 1 0 2944 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1621523292
transform 1 0 3772 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1621523292
transform 1 0 5060 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output287
timestamp 1621523292
transform 1 0 4232 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_28
timestamp 1621523292
transform 1 0 3680 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_30
timestamp 1621523292
transform 1 0 3864 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_38
timestamp 1621523292
transform 1 0 4600 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_42
timestamp 1621523292
transform 1 0 4968 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1621523292
transform 1 0 6440 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1621523292
transform 1 0 5796 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1621523292
transform 1 0 6900 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_47
timestamp 1621523292
transform 1 0 5428 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_54
timestamp 1621523292
transform 1 0 6072 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_59
timestamp 1621523292
transform 1 0 6532 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1621523292
transform 1 0 9108 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1621523292
transform 1 0 7544 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input173
timestamp 1621523292
transform 1 0 8188 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_66
timestamp 1621523292
transform 1 0 7176 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_73
timestamp 1621523292
transform 1 0 7820 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_80
timestamp 1621523292
transform 1 0 8464 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_86
timestamp 1621523292
transform 1 0 9016 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1621523292
transform 1 0 9568 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1621523292
transform 1 0 10212 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input127
timestamp 1621523292
transform 1 0 10856 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_88
timestamp 1621523292
transform 1 0 9200 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_95
timestamp 1621523292
transform 1 0 9844 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_102
timestamp 1621523292
transform 1 0 10488 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_109
timestamp 1621523292
transform 1 0 11132 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1621523292
transform 1 0 11776 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input130
timestamp 1621523292
transform 1 0 12236 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input131
timestamp 1621523292
transform 1 0 12880 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_115
timestamp 1621523292
transform 1 0 11684 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_117
timestamp 1621523292
transform 1 0 11868 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_124
timestamp 1621523292
transform 1 0 12512 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_131
timestamp 1621523292
transform 1 0 13156 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1621523292
transform 1 0 14444 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input132
timestamp 1621523292
transform 1 0 13524 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input133
timestamp 1621523292
transform 1 0 14904 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_138
timestamp 1621523292
transform 1 0 13800 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_144
timestamp 1621523292
transform 1 0 14352 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_146
timestamp 1621523292
transform 1 0 14536 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1621523292
transform 1 0 17112 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input134
timestamp 1621523292
transform 1 0 15548 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input135
timestamp 1621523292
transform 1 0 16192 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_153
timestamp 1621523292
transform 1 0 15180 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_160
timestamp 1621523292
transform 1 0 15824 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_167
timestamp 1621523292
transform 1 0 16468 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_173
timestamp 1621523292
transform 1 0 17020 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1621523292
transform 1 0 17572 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1621523292
transform 1 0 18216 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1621523292
transform 1 0 18860 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_175
timestamp 1621523292
transform 1 0 17204 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_182
timestamp 1621523292
transform 1 0 17848 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_189
timestamp 1621523292
transform 1 0 18492 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_196
timestamp 1621523292
transform 1 0 19136 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1621523292
transform 1 0 19780 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 1621523292
transform 1 0 20240 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1621523292
transform 1 0 20884 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_202
timestamp 1621523292
transform 1 0 19688 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_204
timestamp 1621523292
transform 1 0 19872 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_211
timestamp 1621523292
transform 1 0 20516 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_218
timestamp 1621523292
transform 1 0 21160 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1621523292
transform 1 0 22448 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1621523292
transform 1 0 21528 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 1621523292
transform 1 0 22908 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_225
timestamp 1621523292
transform 1 0 21804 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_231
timestamp 1621523292
transform 1 0 22356 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_233
timestamp 1621523292
transform 1 0 22540 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_240
timestamp 1621523292
transform 1 0 23184 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1621523292
transform 1 0 25116 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1621523292
transform 1 0 23552 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 1621523292
transform 1 0 24196 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_247
timestamp 1621523292
transform 1 0 23828 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_254
timestamp 1621523292
transform 1 0 24472 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_260
timestamp 1621523292
transform 1 0 25024 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_262
timestamp 1621523292
transform 1 0 25208 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1621523292
transform 1 0 25576 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1621523292
transform 1 0 26220 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1621523292
transform 1 0 26864 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_269
timestamp 1621523292
transform 1 0 25852 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_276
timestamp 1621523292
transform 1 0 26496 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_283
timestamp 1621523292
transform 1 0 27140 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1621523292
transform 1 0 27784 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1621523292
transform 1 0 28244 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input121
timestamp 1621523292
transform 1 0 28888 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_289
timestamp 1621523292
transform 1 0 27692 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_291
timestamp 1621523292
transform 1 0 27876 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_298
timestamp 1621523292
transform 1 0 28520 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_305
timestamp 1621523292
transform 1 0 29164 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1621523292
transform 1 0 30452 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input122
timestamp 1621523292
transform 1 0 29532 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input123
timestamp 1621523292
transform 1 0 30912 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_312
timestamp 1621523292
transform 1 0 29808 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_318
timestamp 1621523292
transform 1 0 30360 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_320
timestamp 1621523292
transform 1 0 30544 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_327
timestamp 1621523292
transform 1 0 31188 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1621523292
transform 1 0 33120 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input124
timestamp 1621523292
transform 1 0 31556 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input125
timestamp 1621523292
transform 1 0 32200 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_334
timestamp 1621523292
transform 1 0 31832 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_341
timestamp 1621523292
transform 1 0 32476 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_347
timestamp 1621523292
transform 1 0 33028 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_349
timestamp 1621523292
transform 1 0 33212 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input126
timestamp 1621523292
transform 1 0 33580 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input128
timestamp 1621523292
transform 1 0 34224 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input129
timestamp 1621523292
transform 1 0 34868 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_356
timestamp 1621523292
transform 1 0 33856 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_363
timestamp 1621523292
transform 1 0 34500 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_370
timestamp 1621523292
transform 1 0 35144 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1621523292
transform 1 0 35788 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1621523292
transform 1 0 36248 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1621523292
transform 1 0 36892 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_376
timestamp 1621523292
transform 1 0 35696 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_378
timestamp 1621523292
transform 1 0 35880 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_385
timestamp 1621523292
transform 1 0 36524 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_392
timestamp 1621523292
transform 1 0 37168 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1621523292
transform 1 0 38456 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1621523292
transform 1 0 37536 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input164
timestamp 1621523292
transform 1 0 38916 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_399
timestamp 1621523292
transform 1 0 37812 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_405
timestamp 1621523292
transform 1 0 38364 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_407
timestamp 1621523292
transform 1 0 38548 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_414
timestamp 1621523292
transform 1 0 39192 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1621523292
transform 1 0 41124 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1621523292
transform 1 0 39560 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1621523292
transform 1 0 40204 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_421
timestamp 1621523292
transform 1 0 39836 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_428
timestamp 1621523292
transform 1 0 40480 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_434
timestamp 1621523292
transform 1 0 41032 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_436
timestamp 1621523292
transform 1 0 41216 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1621523292
transform 1 0 42136 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1621523292
transform 1 0 42964 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_444
timestamp 1621523292
transform 1 0 41952 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_449
timestamp 1621523292
transform 1 0 42412 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_458
timestamp 1621523292
transform 1 0 43240 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1621523292
transform 1 0 43792 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1621523292
transform 1 0 44252 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1621523292
transform 1 0 44896 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_465
timestamp 1621523292
transform 1 0 43884 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_472
timestamp 1621523292
transform 1 0 44528 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_479
timestamp 1621523292
transform 1 0 45172 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1621523292
transform 1 0 46460 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1621523292
transform 1 0 45540 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1621523292
transform 1 0 46920 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_486
timestamp 1621523292
transform 1 0 45816 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_492
timestamp 1621523292
transform 1 0 46368 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_494
timestamp 1621523292
transform 1 0 46552 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_501
timestamp 1621523292
transform 1 0 47196 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1621523292
transform 1 0 49128 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1621523292
transform 1 0 47564 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input146
timestamp 1621523292
transform 1 0 48208 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_508
timestamp 1621523292
transform 1 0 47840 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_515
timestamp 1621523292
transform 1 0 48484 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_521
timestamp 1621523292
transform 1 0 49036 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_523
timestamp 1621523292
transform 1 0 49220 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1621523292
transform 1 0 49588 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1621523292
transform 1 0 50232 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1621523292
transform 1 0 50876 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_530
timestamp 1621523292
transform 1 0 49864 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_537
timestamp 1621523292
transform 1 0 50508 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_544
timestamp 1621523292
transform 1 0 51152 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1621523292
transform 1 0 51796 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output253
timestamp 1621523292
transform 1 0 52992 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output254
timestamp 1621523292
transform 1 0 52256 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_550
timestamp 1621523292
transform 1 0 51704 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_552
timestamp 1621523292
transform 1 0 51888 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_560
timestamp 1621523292
transform 1 0 52624 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1621523292
transform 1 0 54464 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output206
timestamp 1621523292
transform 1 0 55200 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output252
timestamp 1621523292
transform 1 0 53728 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_568
timestamp 1621523292
transform 1 0 53360 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_576
timestamp 1621523292
transform 1 0 54096 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_581
timestamp 1621523292
transform 1 0 54556 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_587
timestamp 1621523292
transform 1 0 55108 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _1348_
timestamp 1621523292
transform 1 0 55936 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1621523292
transform 1 0 57132 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_592
timestamp 1621523292
transform 1 0 55568 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_604
timestamp 1621523292
transform 1 0 56672 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_608
timestamp 1621523292
transform 1 0 57040 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_610
timestamp 1621523292
transform 1 0 57224 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1621523292
transform -1 0 58880 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output205
timestamp 1621523292
transform 1 0 57868 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_616
timestamp 1621523292
transform 1 0 57776 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1621523292
transform 1 0 58236 0 1 57120
box -38 -48 406 592
<< labels >>
rlabel metal2 s 5078 59200 5134 60000 6 active
port 0 nsew signal input
rlabel metal3 s 59200 144 60000 264 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 59200 15648 60000 15768 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 59200 17144 60000 17264 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 59200 18640 60000 18760 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 59200 20272 60000 20392 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 59200 21768 60000 21888 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 59200 23400 60000 23520 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 59200 24896 60000 25016 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 59200 26392 60000 26512 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 59200 28024 60000 28144 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 59200 29520 60000 29640 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 59200 31152 60000 31272 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 59200 32648 60000 32768 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 59200 34144 60000 34264 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 59200 35776 60000 35896 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 59200 37272 60000 37392 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 59200 38904 60000 39024 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 59200 40400 60000 40520 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 59200 41896 60000 42016 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 59200 43528 60000 43648 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 59200 45024 60000 45144 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 59200 3136 60000 3256 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 59200 46656 60000 46776 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 59200 48152 60000 48272 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 59200 49648 60000 49768 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 59200 51280 60000 51400 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 59200 52776 60000 52896 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 59200 54408 60000 54528 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 59200 55904 60000 56024 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59200 57400 60000 57520 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 59200 4768 60000 4888 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59200 6264 60000 6384 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 59200 7896 60000 8016 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 59200 9392 60000 9512 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 59200 10888 60000 11008 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 59200 12520 60000 12640 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 59200 14016 60000 14136 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 59200 1096 60000 1216 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 59200 16600 60000 16720 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 59200 18232 60000 18352 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 59200 19728 60000 19848 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 59200 21224 60000 21344 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 59200 22856 60000 22976 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal3 s 59200 24352 60000 24472 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 59200 25984 60000 26104 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal3 s 59200 27480 60000 27600 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal3 s 59200 28976 60000 29096 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal3 s 59200 30608 60000 30728 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal3 s 59200 2728 60000 2848 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 59200 32104 60000 32224 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 59200 33736 60000 33856 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal3 s 59200 35232 60000 35352 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal3 s 59200 36728 60000 36848 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal3 s 59200 38360 60000 38480 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 59200 39856 60000 39976 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 59200 41488 60000 41608 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal3 s 59200 42984 60000 43104 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal3 s 59200 44480 60000 44600 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 59200 46112 60000 46232 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal3 s 59200 4224 60000 4344 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 59200 47608 60000 47728 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 59200 49240 60000 49360 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 59200 50736 60000 50856 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 59200 52232 60000 52352 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 59200 53864 60000 53984 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 59200 55360 60000 55480 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 59200 56992 60000 57112 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 59200 58488 60000 58608 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal3 s 59200 5720 60000 5840 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 59200 7352 60000 7472 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 59200 8848 60000 8968 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 59200 10480 60000 10600 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal3 s 59200 11976 60000 12096 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal3 s 59200 13472 60000 13592 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal3 s 59200 15104 60000 15224 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 59200 552 60000 672 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 59200 16056 60000 16176 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 59200 17688 60000 17808 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 59200 19184 60000 19304 6 io_out[12]
port 80 nsew signal tristate
rlabel metal3 s 59200 20816 60000 20936 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 59200 22312 60000 22432 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 59200 23808 60000 23928 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 59200 25440 60000 25560 6 io_out[16]
port 84 nsew signal tristate
rlabel metal3 s 59200 26936 60000 27056 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 59200 28568 60000 28688 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 59200 30064 60000 30184 6 io_out[19]
port 87 nsew signal tristate
rlabel metal3 s 59200 2184 60000 2304 6 io_out[1]
port 88 nsew signal tristate
rlabel metal3 s 59200 31560 60000 31680 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 59200 33192 60000 33312 6 io_out[21]
port 90 nsew signal tristate
rlabel metal3 s 59200 34688 60000 34808 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 59200 36320 60000 36440 6 io_out[23]
port 92 nsew signal tristate
rlabel metal3 s 59200 37816 60000 37936 6 io_out[24]
port 93 nsew signal tristate
rlabel metal3 s 59200 39312 60000 39432 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 59200 40944 60000 41064 6 io_out[26]
port 95 nsew signal tristate
rlabel metal3 s 59200 42440 60000 42560 6 io_out[27]
port 96 nsew signal tristate
rlabel metal3 s 59200 44072 60000 44192 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 59200 45568 60000 45688 6 io_out[29]
port 98 nsew signal tristate
rlabel metal3 s 59200 3680 60000 3800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 59200 47064 60000 47184 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 59200 48696 60000 48816 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 59200 50192 60000 50312 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 59200 51824 60000 51944 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 59200 53320 60000 53440 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 59200 54816 60000 54936 6 io_out[35]
port 105 nsew signal tristate
rlabel metal3 s 59200 56448 60000 56568 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 59200 57944 60000 58064 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 59200 5312 60000 5432 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 59200 6808 60000 6928 6 io_out[4]
port 109 nsew signal tristate
rlabel metal3 s 59200 8304 60000 8424 6 io_out[5]
port 110 nsew signal tristate
rlabel metal3 s 59200 9936 60000 10056 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 59200 11432 60000 11552 6 io_out[7]
port 112 nsew signal tristate
rlabel metal3 s 59200 13064 60000 13184 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 59200 14560 60000 14680 6 io_out[9]
port 114 nsew signal tristate
rlabel metal2 s 59542 59200 59598 60000 6 irq[0]
port 115 nsew signal tristate
rlabel metal3 s 59200 59032 60000 59152 6 irq[1]
port 116 nsew signal tristate
rlabel metal3 s 59200 59576 60000 59696 6 irq[2]
port 117 nsew signal tristate
rlabel metal2 s 478 0 534 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[3]
port 143 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_in[4]
port 144 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 la_data_in[5]
port 145 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 la_data_in[6]
port 146 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 la_data_in[7]
port 147 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 la_data_in[8]
port 148 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 la_data_in[9]
port 149 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_out[0]
port 150 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 la_data_out[10]
port 151 nsew signal tristate
rlabel metal2 s 40774 0 40830 800 6 la_data_out[11]
port 152 nsew signal tristate
rlabel metal2 s 41694 0 41750 800 6 la_data_out[12]
port 153 nsew signal tristate
rlabel metal2 s 42614 0 42670 800 6 la_data_out[13]
port 154 nsew signal tristate
rlabel metal2 s 43534 0 43590 800 6 la_data_out[14]
port 155 nsew signal tristate
rlabel metal2 s 44454 0 44510 800 6 la_data_out[15]
port 156 nsew signal tristate
rlabel metal2 s 45466 0 45522 800 6 la_data_out[16]
port 157 nsew signal tristate
rlabel metal2 s 46386 0 46442 800 6 la_data_out[17]
port 158 nsew signal tristate
rlabel metal2 s 47306 0 47362 800 6 la_data_out[18]
port 159 nsew signal tristate
rlabel metal2 s 48226 0 48282 800 6 la_data_out[19]
port 160 nsew signal tristate
rlabel metal2 s 31390 0 31446 800 6 la_data_out[1]
port 161 nsew signal tristate
rlabel metal2 s 49146 0 49202 800 6 la_data_out[20]
port 162 nsew signal tristate
rlabel metal2 s 50066 0 50122 800 6 la_data_out[21]
port 163 nsew signal tristate
rlabel metal2 s 51078 0 51134 800 6 la_data_out[22]
port 164 nsew signal tristate
rlabel metal2 s 51998 0 52054 800 6 la_data_out[23]
port 165 nsew signal tristate
rlabel metal2 s 52918 0 52974 800 6 la_data_out[24]
port 166 nsew signal tristate
rlabel metal2 s 53838 0 53894 800 6 la_data_out[25]
port 167 nsew signal tristate
rlabel metal2 s 54758 0 54814 800 6 la_data_out[26]
port 168 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 la_data_out[27]
port 169 nsew signal tristate
rlabel metal2 s 56690 0 56746 800 6 la_data_out[28]
port 170 nsew signal tristate
rlabel metal2 s 57610 0 57666 800 6 la_data_out[29]
port 171 nsew signal tristate
rlabel metal2 s 32310 0 32366 800 6 la_data_out[2]
port 172 nsew signal tristate
rlabel metal2 s 58530 0 58586 800 6 la_data_out[30]
port 173 nsew signal tristate
rlabel metal2 s 59450 0 59506 800 6 la_data_out[31]
port 174 nsew signal tristate
rlabel metal2 s 33230 0 33286 800 6 la_data_out[3]
port 175 nsew signal tristate
rlabel metal2 s 34150 0 34206 800 6 la_data_out[4]
port 176 nsew signal tristate
rlabel metal2 s 35070 0 35126 800 6 la_data_out[5]
port 177 nsew signal tristate
rlabel metal2 s 36082 0 36138 800 6 la_data_out[6]
port 178 nsew signal tristate
rlabel metal2 s 37002 0 37058 800 6 la_data_out[7]
port 179 nsew signal tristate
rlabel metal2 s 37922 0 37978 800 6 la_data_out[8]
port 180 nsew signal tristate
rlabel metal2 s 38842 0 38898 800 6 la_data_out[9]
port 181 nsew signal tristate
rlabel metal3 s 0 30336 800 30456 6 la_oenb[0]
port 182 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la_oenb[10]
port 183 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 la_oenb[11]
port 184 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 la_oenb[12]
port 185 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 la_oenb[13]
port 186 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 la_oenb[14]
port 187 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 la_oenb[15]
port 188 nsew signal input
rlabel metal3 s 0 45296 800 45416 6 la_oenb[16]
port 189 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 la_oenb[17]
port 190 nsew signal input
rlabel metal3 s 0 47200 800 47320 6 la_oenb[18]
port 191 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 la_oenb[19]
port 192 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la_oenb[1]
port 193 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 la_oenb[20]
port 194 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 la_oenb[21]
port 195 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 la_oenb[22]
port 196 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 la_oenb[23]
port 197 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 la_oenb[24]
port 198 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_oenb[25]
port 199 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 la_oenb[26]
port 200 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 la_oenb[27]
port 201 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la_oenb[28]
port 202 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 la_oenb[29]
port 203 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 la_oenb[2]
port 204 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 la_oenb[30]
port 205 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 la_oenb[31]
port 206 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 la_oenb[3]
port 207 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 la_oenb[4]
port 208 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 la_oenb[5]
port 209 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 la_oenb[6]
port 210 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 la_oenb[7]
port 211 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 la_oenb[8]
port 212 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_oenb[9]
port 213 nsew signal input
rlabel metal2 s 386 59200 442 60000 6 wb_clk_i
port 214 nsew signal input
rlabel metal2 s 1122 59200 1178 60000 6 wb_rst_i
port 215 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 wbs_ack_o
port 216 nsew signal tristate
rlabel metal2 s 9034 59200 9090 60000 6 wbs_adr_i[0]
port 217 nsew signal input
rlabel metal2 s 16946 59200 17002 60000 6 wbs_adr_i[10]
port 218 nsew signal input
rlabel metal2 s 17682 59200 17738 60000 6 wbs_adr_i[11]
port 219 nsew signal input
rlabel metal2 s 18510 59200 18566 60000 6 wbs_adr_i[12]
port 220 nsew signal input
rlabel metal2 s 19246 59200 19302 60000 6 wbs_adr_i[13]
port 221 nsew signal input
rlabel metal2 s 20074 59200 20130 60000 6 wbs_adr_i[14]
port 222 nsew signal input
rlabel metal2 s 20902 59200 20958 60000 6 wbs_adr_i[15]
port 223 nsew signal input
rlabel metal2 s 21638 59200 21694 60000 6 wbs_adr_i[16]
port 224 nsew signal input
rlabel metal2 s 22466 59200 22522 60000 6 wbs_adr_i[17]
port 225 nsew signal input
rlabel metal2 s 23202 59200 23258 60000 6 wbs_adr_i[18]
port 226 nsew signal input
rlabel metal2 s 24030 59200 24086 60000 6 wbs_adr_i[19]
port 227 nsew signal input
rlabel metal2 s 9770 59200 9826 60000 6 wbs_adr_i[1]
port 228 nsew signal input
rlabel metal2 s 24766 59200 24822 60000 6 wbs_adr_i[20]
port 229 nsew signal input
rlabel metal2 s 25594 59200 25650 60000 6 wbs_adr_i[21]
port 230 nsew signal input
rlabel metal2 s 26422 59200 26478 60000 6 wbs_adr_i[22]
port 231 nsew signal input
rlabel metal2 s 27158 59200 27214 60000 6 wbs_adr_i[23]
port 232 nsew signal input
rlabel metal2 s 27986 59200 28042 60000 6 wbs_adr_i[24]
port 233 nsew signal input
rlabel metal2 s 28722 59200 28778 60000 6 wbs_adr_i[25]
port 234 nsew signal input
rlabel metal2 s 29550 59200 29606 60000 6 wbs_adr_i[26]
port 235 nsew signal input
rlabel metal2 s 30378 59200 30434 60000 6 wbs_adr_i[27]
port 236 nsew signal input
rlabel metal2 s 31114 59200 31170 60000 6 wbs_adr_i[28]
port 237 nsew signal input
rlabel metal2 s 31942 59200 31998 60000 6 wbs_adr_i[29]
port 238 nsew signal input
rlabel metal2 s 10598 59200 10654 60000 6 wbs_adr_i[2]
port 239 nsew signal input
rlabel metal2 s 32678 59200 32734 60000 6 wbs_adr_i[30]
port 240 nsew signal input
rlabel metal2 s 33506 59200 33562 60000 6 wbs_adr_i[31]
port 241 nsew signal input
rlabel metal2 s 11426 59200 11482 60000 6 wbs_adr_i[3]
port 242 nsew signal input
rlabel metal2 s 12162 59200 12218 60000 6 wbs_adr_i[4]
port 243 nsew signal input
rlabel metal2 s 12990 59200 13046 60000 6 wbs_adr_i[5]
port 244 nsew signal input
rlabel metal2 s 13726 59200 13782 60000 6 wbs_adr_i[6]
port 245 nsew signal input
rlabel metal2 s 14554 59200 14610 60000 6 wbs_adr_i[7]
port 246 nsew signal input
rlabel metal2 s 15382 59200 15438 60000 6 wbs_adr_i[8]
port 247 nsew signal input
rlabel metal2 s 16118 59200 16174 60000 6 wbs_adr_i[9]
port 248 nsew signal input
rlabel metal2 s 2686 59200 2742 60000 6 wbs_cyc_i
port 249 nsew signal input
rlabel metal2 s 34242 59200 34298 60000 6 wbs_dat_i[0]
port 250 nsew signal input
rlabel metal2 s 42154 59200 42210 60000 6 wbs_dat_i[10]
port 251 nsew signal input
rlabel metal2 s 42982 59200 43038 60000 6 wbs_dat_i[11]
port 252 nsew signal input
rlabel metal2 s 43718 59200 43774 60000 6 wbs_dat_i[12]
port 253 nsew signal input
rlabel metal2 s 44546 59200 44602 60000 6 wbs_dat_i[13]
port 254 nsew signal input
rlabel metal2 s 45374 59200 45430 60000 6 wbs_dat_i[14]
port 255 nsew signal input
rlabel metal2 s 46110 59200 46166 60000 6 wbs_dat_i[15]
port 256 nsew signal input
rlabel metal2 s 46938 59200 46994 60000 6 wbs_dat_i[16]
port 257 nsew signal input
rlabel metal2 s 47674 59200 47730 60000 6 wbs_dat_i[17]
port 258 nsew signal input
rlabel metal2 s 48502 59200 48558 60000 6 wbs_dat_i[18]
port 259 nsew signal input
rlabel metal2 s 49238 59200 49294 60000 6 wbs_dat_i[19]
port 260 nsew signal input
rlabel metal2 s 35070 59200 35126 60000 6 wbs_dat_i[1]
port 261 nsew signal input
rlabel metal2 s 50066 59200 50122 60000 6 wbs_dat_i[20]
port 262 nsew signal input
rlabel metal2 s 50894 59200 50950 60000 6 wbs_dat_i[21]
port 263 nsew signal input
rlabel metal2 s 51630 59200 51686 60000 6 wbs_dat_i[22]
port 264 nsew signal input
rlabel metal2 s 52458 59200 52514 60000 6 wbs_dat_i[23]
port 265 nsew signal input
rlabel metal2 s 53194 59200 53250 60000 6 wbs_dat_i[24]
port 266 nsew signal input
rlabel metal2 s 54022 59200 54078 60000 6 wbs_dat_i[25]
port 267 nsew signal input
rlabel metal2 s 54758 59200 54814 60000 6 wbs_dat_i[26]
port 268 nsew signal input
rlabel metal2 s 55586 59200 55642 60000 6 wbs_dat_i[27]
port 269 nsew signal input
rlabel metal2 s 56414 59200 56470 60000 6 wbs_dat_i[28]
port 270 nsew signal input
rlabel metal2 s 57150 59200 57206 60000 6 wbs_dat_i[29]
port 271 nsew signal input
rlabel metal2 s 35898 59200 35954 60000 6 wbs_dat_i[2]
port 272 nsew signal input
rlabel metal2 s 57978 59200 58034 60000 6 wbs_dat_i[30]
port 273 nsew signal input
rlabel metal2 s 58714 59200 58770 60000 6 wbs_dat_i[31]
port 274 nsew signal input
rlabel metal2 s 36634 59200 36690 60000 6 wbs_dat_i[3]
port 275 nsew signal input
rlabel metal2 s 37462 59200 37518 60000 6 wbs_dat_i[4]
port 276 nsew signal input
rlabel metal2 s 38198 59200 38254 60000 6 wbs_dat_i[5]
port 277 nsew signal input
rlabel metal2 s 39026 59200 39082 60000 6 wbs_dat_i[6]
port 278 nsew signal input
rlabel metal2 s 39762 59200 39818 60000 6 wbs_dat_i[7]
port 279 nsew signal input
rlabel metal2 s 40590 59200 40646 60000 6 wbs_dat_i[8]
port 280 nsew signal input
rlabel metal2 s 41418 59200 41474 60000 6 wbs_dat_i[9]
port 281 nsew signal input
rlabel metal3 s 0 416 800 536 6 wbs_dat_o[0]
port 282 nsew signal tristate
rlabel metal3 s 0 9664 800 9784 6 wbs_dat_o[10]
port 283 nsew signal tristate
rlabel metal3 s 0 10616 800 10736 6 wbs_dat_o[11]
port 284 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 wbs_dat_o[12]
port 285 nsew signal tristate
rlabel metal3 s 0 12520 800 12640 6 wbs_dat_o[13]
port 286 nsew signal tristate
rlabel metal3 s 0 13472 800 13592 6 wbs_dat_o[14]
port 287 nsew signal tristate
rlabel metal3 s 0 14424 800 14544 6 wbs_dat_o[15]
port 288 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 wbs_dat_o[16]
port 289 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 wbs_dat_o[17]
port 290 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 wbs_dat_o[18]
port 291 nsew signal tristate
rlabel metal3 s 0 18096 800 18216 6 wbs_dat_o[19]
port 292 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 wbs_dat_o[1]
port 293 nsew signal tristate
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_o[20]
port 294 nsew signal tristate
rlabel metal3 s 0 20000 800 20120 6 wbs_dat_o[21]
port 295 nsew signal tristate
rlabel metal3 s 0 20952 800 21072 6 wbs_dat_o[22]
port 296 nsew signal tristate
rlabel metal3 s 0 21904 800 22024 6 wbs_dat_o[23]
port 297 nsew signal tristate
rlabel metal3 s 0 22856 800 22976 6 wbs_dat_o[24]
port 298 nsew signal tristate
rlabel metal3 s 0 23808 800 23928 6 wbs_dat_o[25]
port 299 nsew signal tristate
rlabel metal3 s 0 24760 800 24880 6 wbs_dat_o[26]
port 300 nsew signal tristate
rlabel metal3 s 0 25712 800 25832 6 wbs_dat_o[27]
port 301 nsew signal tristate
rlabel metal3 s 0 26528 800 26648 6 wbs_dat_o[28]
port 302 nsew signal tristate
rlabel metal3 s 0 27480 800 27600 6 wbs_dat_o[29]
port 303 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 wbs_dat_o[2]
port 304 nsew signal tristate
rlabel metal3 s 0 28432 800 28552 6 wbs_dat_o[30]
port 305 nsew signal tristate
rlabel metal3 s 0 29384 800 29504 6 wbs_dat_o[31]
port 306 nsew signal tristate
rlabel metal3 s 0 3136 800 3256 6 wbs_dat_o[3]
port 307 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[4]
port 308 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 wbs_dat_o[5]
port 309 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 wbs_dat_o[6]
port 310 nsew signal tristate
rlabel metal3 s 0 6944 800 7064 6 wbs_dat_o[7]
port 311 nsew signal tristate
rlabel metal3 s 0 7896 800 8016 6 wbs_dat_o[8]
port 312 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 wbs_dat_o[9]
port 313 nsew signal tristate
rlabel metal2 s 5906 59200 5962 60000 6 wbs_sel_i[0]
port 314 nsew signal input
rlabel metal2 s 6642 59200 6698 60000 6 wbs_sel_i[1]
port 315 nsew signal input
rlabel metal2 s 7470 59200 7526 60000 6 wbs_sel_i[2]
port 316 nsew signal input
rlabel metal2 s 8206 59200 8262 60000 6 wbs_sel_i[3]
port 317 nsew signal input
rlabel metal2 s 1950 59200 2006 60000 6 wbs_stb_i
port 318 nsew signal input
rlabel metal2 s 3514 59200 3570 60000 6 wbs_we_i
port 319 nsew signal input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 320 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 321 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 322 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 323 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 57664 6 vccd2
port 324 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 57664 6 vccd2
port 325 nsew power bidirectional
rlabel metal4 s 50948 2176 51268 57664 6 vssd2
port 326 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 57664 6 vssd2
port 327 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 57664 6 vdda1
port 328 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 57664 6 vdda1
port 329 nsew power bidirectional
rlabel metal4 s 51608 2176 51928 57664 6 vssa1
port 330 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 57664 6 vssa1
port 331 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 57664 6 vdda2
port 332 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 57664 6 vdda2
port 333 nsew power bidirectional
rlabel metal4 s 52268 2176 52588 57664 6 vssa2
port 334 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 57664 6 vssa2
port 335 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
