magic
tech sky130A
magscale 1 2
timestamp 1621574425
<< locali >>
rect 32045 31875 32079 31977
rect 15209 30583 15243 30753
rect 28457 30039 28491 30345
rect 27353 28407 27387 28645
rect 29009 24599 29043 24701
rect 21741 24191 21775 24361
rect 13185 23103 13219 23273
rect 4721 21471 4755 21573
rect 16773 19159 16807 19329
rect 56333 14943 56367 15113
<< viali >>
rect 3249 57545 3283 57579
rect 29745 57545 29779 57579
rect 32137 57545 32171 57579
rect 36277 57545 36311 57579
rect 2053 57477 2087 57511
rect 10425 57477 10459 57511
rect 26755 57477 26789 57511
rect 26893 57477 26927 57511
rect 37565 57477 37599 57511
rect 53297 57477 53331 57511
rect 55597 57477 55631 57511
rect 12725 57409 12759 57443
rect 24501 57409 24535 57443
rect 26985 57409 27019 57443
rect 29193 57409 29227 57443
rect 54033 57409 54067 57443
rect 58173 57409 58207 57443
rect 4261 57341 4295 57375
rect 4445 57341 4479 57375
rect 5365 57341 5399 57375
rect 6929 57341 6963 57375
rect 7573 57341 7607 57375
rect 8217 57341 8251 57375
rect 9597 57341 9631 57375
rect 10241 57341 10275 57375
rect 11069 57341 11103 57375
rect 12265 57341 12299 57375
rect 12817 57341 12851 57375
rect 13461 57341 13495 57375
rect 15117 57341 15151 57375
rect 15761 57341 15795 57375
rect 16405 57341 16439 57375
rect 17785 57341 17819 57375
rect 18429 57341 18463 57375
rect 19073 57341 19107 57375
rect 20453 57341 20487 57375
rect 21097 57341 21131 57375
rect 21741 57341 21775 57375
rect 23121 57341 23155 57375
rect 24317 57341 24351 57375
rect 24593 57341 24627 57375
rect 25973 57341 26007 57375
rect 26157 57341 26191 57375
rect 28449 57341 28483 57375
rect 29101 57341 29135 57375
rect 29929 57341 29963 57375
rect 31493 57341 31527 57375
rect 32321 57341 32355 57375
rect 33793 57341 33827 57375
rect 34437 57341 34471 57375
rect 35081 57341 35115 57375
rect 36461 57341 36495 57375
rect 37105 57341 37139 57375
rect 37749 57341 37783 57375
rect 39129 57341 39163 57375
rect 39773 57341 39807 57375
rect 40233 57341 40267 57375
rect 41613 57341 41647 57375
rect 42257 57341 42291 57375
rect 42993 57341 43027 57375
rect 44281 57341 44315 57375
rect 44925 57341 44959 57375
rect 45569 57341 45603 57375
rect 46949 57341 46983 57375
rect 47593 57341 47627 57375
rect 48237 57341 48271 57375
rect 49617 57341 49651 57375
rect 50261 57341 50295 57375
rect 50905 57341 50939 57375
rect 52377 57341 52411 57375
rect 56057 57341 56091 57375
rect 56241 57341 56275 57375
rect 1869 57273 1903 57307
rect 3157 57273 3191 57307
rect 4905 57273 4939 57307
rect 26617 57273 26651 57307
rect 53113 57273 53147 57307
rect 53849 57273 53883 57307
rect 55413 57273 55447 57307
rect 56701 57273 56735 57307
rect 57989 57273 58023 57307
rect 5549 57205 5583 57239
rect 9781 57205 9815 57239
rect 11253 57205 11287 57239
rect 12449 57205 12483 57239
rect 13645 57205 13679 57239
rect 14933 57205 14967 57239
rect 15577 57205 15611 57239
rect 16221 57205 16255 57239
rect 17601 57205 17635 57239
rect 18245 57205 18279 57239
rect 18889 57205 18923 57239
rect 20269 57205 20303 57239
rect 20913 57205 20947 57239
rect 21557 57205 21591 57239
rect 22937 57205 22971 57239
rect 24133 57205 24167 57239
rect 26065 57205 26099 57239
rect 27261 57205 27295 57239
rect 28273 57205 28307 57239
rect 31585 57205 31619 57239
rect 33609 57205 33643 57239
rect 34253 57205 34287 57239
rect 35265 57205 35299 57239
rect 36921 57205 36955 57239
rect 38945 57205 38979 57239
rect 39589 57205 39623 57239
rect 40417 57205 40451 57239
rect 4905 57001 4939 57035
rect 10609 57001 10643 57035
rect 16129 57001 16163 57035
rect 23673 57001 23707 57035
rect 27353 57001 27387 57035
rect 35725 57001 35759 57035
rect 55229 57001 55263 57035
rect 58173 57001 58207 57035
rect 4537 56933 4571 56967
rect 4629 56933 4663 56967
rect 13093 56933 13127 56967
rect 14749 56933 14783 56967
rect 17601 56933 17635 56967
rect 19993 56933 20027 56967
rect 23029 56933 23063 56967
rect 57069 56933 57103 56967
rect 1409 56865 1443 56899
rect 2145 56865 2179 56899
rect 3157 56865 3191 56899
rect 4746 56865 4780 56899
rect 8217 56865 8251 56899
rect 10793 56865 10827 56899
rect 11713 56865 11747 56899
rect 11989 56865 12023 56899
rect 14896 56865 14930 56899
rect 16313 56865 16347 56899
rect 17748 56865 17782 56899
rect 20729 56865 20763 56899
rect 21189 56865 21223 56899
rect 21336 56865 21370 56899
rect 22569 56865 22603 56899
rect 25789 56865 25823 56899
rect 26709 56865 26743 56899
rect 26856 56865 26890 56899
rect 27997 56865 28031 56899
rect 28641 56865 28675 56899
rect 31300 56865 31334 56899
rect 33600 56865 33634 56899
rect 35909 56865 35943 56899
rect 36553 56865 36587 56899
rect 37197 56865 37231 56899
rect 37841 56865 37875 56899
rect 39773 56865 39807 56899
rect 42165 56865 42199 56899
rect 51457 56865 51491 56899
rect 52101 56865 52135 56899
rect 54125 56865 54159 56899
rect 56885 56865 56919 56899
rect 4261 56797 4295 56831
rect 11805 56797 11839 56831
rect 12173 56797 12207 56831
rect 15117 56797 15151 56831
rect 17969 56797 18003 56831
rect 18337 56797 18371 56831
rect 20140 56797 20174 56831
rect 20361 56797 20395 56831
rect 21557 56797 21591 56831
rect 21925 56797 21959 56831
rect 23397 56797 23431 56831
rect 26065 56797 26099 56831
rect 27077 56797 27111 56831
rect 29193 56797 29227 56831
rect 29285 56797 29319 56831
rect 31033 56797 31067 56831
rect 33333 56797 33367 56831
rect 54585 56797 54619 56831
rect 54769 56797 54803 56831
rect 57529 56797 57563 56831
rect 57713 56797 57747 56831
rect 13277 56729 13311 56763
rect 15025 56729 15059 56763
rect 15393 56729 15427 56763
rect 17877 56729 17911 56763
rect 20269 56729 20303 56763
rect 22385 56729 22419 56763
rect 23305 56729 23339 56763
rect 29101 56729 29135 56763
rect 32413 56729 32447 56763
rect 37013 56729 37047 56763
rect 53481 56729 53515 56763
rect 3249 56661 3283 56695
rect 21465 56661 21499 56695
rect 23167 56661 23201 56695
rect 25605 56661 25639 56695
rect 25973 56661 26007 56695
rect 26985 56661 27019 56695
rect 28089 56661 28123 56695
rect 29009 56661 29043 56695
rect 34713 56661 34747 56695
rect 36369 56661 36403 56695
rect 37657 56661 37691 56695
rect 3801 56457 3835 56491
rect 4813 56457 4847 56491
rect 22845 56457 22879 56491
rect 24869 56457 24903 56491
rect 26709 56457 26743 56491
rect 31493 56457 31527 56491
rect 33222 56457 33256 56491
rect 33333 56457 33367 56491
rect 34989 56457 35023 56491
rect 54217 56457 54251 56491
rect 55137 56457 55171 56491
rect 2697 56389 2731 56423
rect 3341 56389 3375 56423
rect 3709 56389 3743 56423
rect 12173 56389 12207 56423
rect 33517 56389 33551 56423
rect 3893 56321 3927 56355
rect 33425 56321 33459 56355
rect 34538 56321 34572 56355
rect 55781 56321 55815 56355
rect 56241 56321 56275 56355
rect 1409 56253 1443 56287
rect 2053 56253 2087 56287
rect 2881 56253 2915 56287
rect 4997 56253 5031 56287
rect 12081 56253 12115 56287
rect 12357 56253 12391 56287
rect 23029 56253 23063 56287
rect 23489 56253 23523 56287
rect 23756 56253 23790 56287
rect 25329 56253 25363 56287
rect 25596 56253 25630 56287
rect 27813 56253 27847 56287
rect 29653 56253 29687 56287
rect 31677 56253 31711 56287
rect 32137 56253 32171 56287
rect 34253 56253 34287 56287
rect 34437 56253 34471 56287
rect 34621 56253 34655 56287
rect 34805 56253 34839 56287
rect 35633 56253 35667 56287
rect 36277 56253 36311 56287
rect 51825 56253 51859 56287
rect 52469 56253 52503 56287
rect 54401 56253 54435 56287
rect 55321 56253 55355 56287
rect 12817 56185 12851 56219
rect 28058 56185 28092 56219
rect 29920 56185 29954 56219
rect 31769 56185 31803 56219
rect 31861 56185 31895 56219
rect 31999 56185 32033 56219
rect 33057 56185 33091 56219
rect 55965 56185 55999 56219
rect 4169 56117 4203 56151
rect 29193 56117 29227 56151
rect 31033 56117 31067 56151
rect 35449 56117 35483 56151
rect 36093 56117 36127 56151
rect 2237 55913 2271 55947
rect 24317 55913 24351 55947
rect 25973 55913 26007 55947
rect 27905 55913 27939 55947
rect 30481 55913 30515 55947
rect 31585 55913 31619 55947
rect 32597 55913 32631 55947
rect 35725 55913 35759 55947
rect 56793 55913 56827 55947
rect 25329 55845 25363 55879
rect 28917 55845 28951 55879
rect 32689 55845 32723 55879
rect 1409 55777 1443 55811
rect 2053 55777 2087 55811
rect 4445 55777 4479 55811
rect 24133 55777 24167 55811
rect 24317 55777 24351 55811
rect 25237 55777 25271 55811
rect 25881 55777 25915 55811
rect 26709 55777 26743 55811
rect 28089 55777 28123 55811
rect 28825 55777 28859 55811
rect 29009 55777 29043 55811
rect 30665 55777 30699 55811
rect 31401 55777 31435 55811
rect 31585 55777 31619 55811
rect 33692 55777 33726 55811
rect 35909 55777 35943 55811
rect 52561 55777 52595 55811
rect 53205 55777 53239 55811
rect 53849 55777 53883 55811
rect 54677 55777 54711 55811
rect 55781 55777 55815 55811
rect 56977 55777 57011 55811
rect 26985 55709 27019 55743
rect 28365 55709 28399 55743
rect 30849 55709 30883 55743
rect 30941 55709 30975 55743
rect 32873 55709 32907 55743
rect 33425 55709 33459 55743
rect 57529 55709 57563 55743
rect 57713 55709 57747 55743
rect 4261 55641 4295 55675
rect 26525 55573 26559 55607
rect 26893 55573 26927 55607
rect 28273 55573 28307 55607
rect 32229 55573 32263 55607
rect 34805 55573 34839 55607
rect 57989 55573 58023 55607
rect 56057 55369 56091 55403
rect 57345 55369 57379 55403
rect 56517 55301 56551 55335
rect 58173 55301 58207 55335
rect 23765 55233 23799 55267
rect 32045 55233 32079 55267
rect 33425 55233 33459 55267
rect 33885 55233 33919 55267
rect 34805 55233 34839 55267
rect 22753 55165 22787 55199
rect 22937 55165 22971 55199
rect 23029 55165 23063 55199
rect 25789 55165 25823 55199
rect 26433 55165 26467 55199
rect 26525 55165 26559 55199
rect 27813 55165 27847 55199
rect 27997 55165 28031 55199
rect 29009 55165 29043 55199
rect 31769 55165 31803 55199
rect 33169 55165 33203 55199
rect 33333 55165 33367 55199
rect 33517 55165 33551 55199
rect 33701 55165 33735 55199
rect 54585 55165 54619 55199
rect 55229 55165 55263 55199
rect 56701 55165 56735 55199
rect 57989 55165 58023 55199
rect 24010 55097 24044 55131
rect 27905 55097 27939 55131
rect 29254 55097 29288 55131
rect 31861 55097 31895 55131
rect 35072 55097 35106 55131
rect 57253 55097 57287 55131
rect 22569 55029 22603 55063
rect 25145 55029 25179 55063
rect 25605 55029 25639 55063
rect 30389 55029 30423 55063
rect 31401 55029 31435 55063
rect 36185 55029 36219 55063
rect 23397 54825 23431 54859
rect 23857 54825 23891 54859
rect 27445 54825 27479 54859
rect 27997 54825 28031 54859
rect 32137 54825 32171 54859
rect 33793 54825 33827 54859
rect 58173 54825 58207 54859
rect 22284 54757 22318 54791
rect 26332 54757 26366 54791
rect 31024 54757 31058 54791
rect 1409 54689 1443 54723
rect 22017 54689 22051 54723
rect 24041 54689 24075 54723
rect 24317 54689 24351 54723
rect 26065 54689 26099 54723
rect 27905 54689 27939 54723
rect 28733 54689 28767 54723
rect 32597 54689 32631 54723
rect 32781 54689 32815 54723
rect 32873 54689 32907 54723
rect 33011 54689 33045 54723
rect 33149 54689 33183 54723
rect 34161 54689 34195 54723
rect 34253 54689 34287 54723
rect 36829 54689 36863 54723
rect 54309 54689 54343 54723
rect 54953 54689 54987 54723
rect 55597 54689 55631 54723
rect 29009 54621 29043 54655
rect 30757 54621 30791 54655
rect 34437 54621 34471 54655
rect 35725 54621 35759 54655
rect 57069 54621 57103 54655
rect 57529 54621 57563 54655
rect 57713 54621 57747 54655
rect 33333 54553 33367 54587
rect 36921 54553 36955 54587
rect 24225 54485 24259 54519
rect 28549 54485 28583 54519
rect 28917 54485 28951 54519
rect 36369 54485 36403 54519
rect 22661 54281 22695 54315
rect 23305 54281 23339 54315
rect 23949 54281 23983 54315
rect 24593 54281 24627 54315
rect 29009 54281 29043 54315
rect 31033 54281 31067 54315
rect 35265 54281 35299 54315
rect 57253 54281 57287 54315
rect 58173 54213 58207 54247
rect 25881 54145 25915 54179
rect 26801 54145 26835 54179
rect 26893 54145 26927 54179
rect 30481 54145 30515 54179
rect 32137 54145 32171 54179
rect 35909 54145 35943 54179
rect 36461 54145 36495 54179
rect 1409 54077 1443 54111
rect 22569 54077 22603 54111
rect 23213 54077 23247 54111
rect 23397 54077 23431 54111
rect 23857 54077 23891 54111
rect 24501 54077 24535 54111
rect 24685 54077 24719 54111
rect 25145 54077 25179 54111
rect 25789 54077 25823 54111
rect 26617 54077 26651 54111
rect 27813 54077 27847 54111
rect 27997 54077 28031 54111
rect 29193 54077 29227 54111
rect 29377 54077 29411 54111
rect 29515 54077 29549 54111
rect 29653 54077 29687 54111
rect 31493 54077 31527 54111
rect 33057 54077 33091 54111
rect 33241 54077 33275 54111
rect 33333 54077 33367 54111
rect 33425 54077 33459 54111
rect 33609 54077 33643 54111
rect 35449 54077 35483 54111
rect 35633 54077 35667 54111
rect 36369 54077 36403 54111
rect 36553 54077 36587 54111
rect 55597 54077 55631 54111
rect 56793 54077 56827 54111
rect 57437 54077 57471 54111
rect 27905 54009 27939 54043
rect 29285 54009 29319 54043
rect 35541 54009 35575 54043
rect 35771 54009 35805 54043
rect 57989 54009 58023 54043
rect 25237 53941 25271 53975
rect 26433 53941 26467 53975
rect 33793 53941 33827 53975
rect 27721 53737 27755 53771
rect 29561 53737 29595 53771
rect 34529 53737 34563 53771
rect 56977 53737 57011 53771
rect 58173 53737 58207 53771
rect 26586 53669 26620 53703
rect 28448 53669 28482 53703
rect 33416 53669 33450 53703
rect 56885 53669 56919 53703
rect 21189 53601 21223 53635
rect 21456 53601 21490 53635
rect 23673 53601 23707 53635
rect 25421 53601 25455 53635
rect 25605 53601 25639 53635
rect 26341 53601 26375 53635
rect 28181 53601 28215 53635
rect 30932 53601 30966 53635
rect 32505 53601 32539 53635
rect 33149 53601 33183 53635
rect 35909 53601 35943 53635
rect 36185 53601 36219 53635
rect 55597 53601 55631 53635
rect 57529 53601 57563 53635
rect 23949 53533 23983 53567
rect 25697 53533 25731 53567
rect 30665 53533 30699 53567
rect 57713 53533 57747 53567
rect 32597 53465 32631 53499
rect 22569 53397 22603 53431
rect 23489 53397 23523 53431
rect 23857 53397 23891 53431
rect 25237 53397 25271 53431
rect 32045 53397 32079 53431
rect 35725 53397 35759 53431
rect 36093 53397 36127 53431
rect 29285 53193 29319 53227
rect 29929 53193 29963 53227
rect 31125 53193 31159 53227
rect 32045 53193 32079 53227
rect 36093 53193 36127 53227
rect 57253 53193 57287 53227
rect 21557 53125 21591 53159
rect 26065 53125 26099 53159
rect 22845 53057 22879 53091
rect 1409 52989 1443 53023
rect 21465 52989 21499 53023
rect 21649 52989 21683 53023
rect 23112 52989 23146 53023
rect 24685 52989 24719 53023
rect 24952 52989 24986 53023
rect 26525 52989 26559 53023
rect 26709 52989 26743 53023
rect 27905 52989 27939 53023
rect 29193 52989 29227 53023
rect 29837 52989 29871 53023
rect 30021 52989 30055 53023
rect 30481 52989 30515 53023
rect 30629 52989 30663 53023
rect 30987 52989 31021 53023
rect 31769 52989 31803 53023
rect 31861 52989 31895 53023
rect 33057 52989 33091 53023
rect 33245 52989 33279 53023
rect 33333 52989 33367 53023
rect 33425 52989 33459 53023
rect 33609 52989 33643 53023
rect 34713 52989 34747 53023
rect 34980 52989 35014 53023
rect 56609 52989 56643 53023
rect 57437 52989 57471 53023
rect 26617 52921 26651 52955
rect 27997 52921 28031 52955
rect 30757 52921 30791 52955
rect 30849 52921 30883 52955
rect 57989 52921 58023 52955
rect 58173 52921 58207 52955
rect 24225 52853 24259 52887
rect 33793 52853 33827 52887
rect 21741 52649 21775 52683
rect 23121 52649 23155 52683
rect 23673 52649 23707 52683
rect 31217 52649 31251 52683
rect 31677 52649 31711 52683
rect 36737 52649 36771 52683
rect 58173 52649 58207 52683
rect 28448 52581 28482 52615
rect 33140 52581 33174 52615
rect 21097 52513 21131 52547
rect 21925 52513 21959 52547
rect 22201 52513 22235 52547
rect 22937 52513 22971 52547
rect 23121 52513 23155 52547
rect 23581 52513 23615 52547
rect 25697 52513 25731 52547
rect 25881 52513 25915 52547
rect 28181 52513 28215 52547
rect 30665 52513 30699 52547
rect 32045 52513 32079 52547
rect 32137 52513 32171 52547
rect 32873 52513 32907 52547
rect 35909 52513 35943 52547
rect 36645 52513 36679 52547
rect 21189 52445 21223 52479
rect 22109 52445 22143 52479
rect 32321 52445 32355 52479
rect 36185 52445 36219 52479
rect 57069 52445 57103 52479
rect 57529 52445 57563 52479
rect 57713 52445 57747 52479
rect 25697 52309 25731 52343
rect 29561 52309 29595 52343
rect 34253 52309 34287 52343
rect 35725 52309 35759 52343
rect 36093 52309 36127 52343
rect 25973 52105 26007 52139
rect 26617 52105 26651 52139
rect 33057 52105 33091 52139
rect 36277 52105 36311 52139
rect 57253 52105 57287 52139
rect 32137 52037 32171 52071
rect 58173 52037 58207 52071
rect 21557 51969 21591 52003
rect 23949 51969 23983 52003
rect 28917 51969 28951 52003
rect 33609 51969 33643 52003
rect 1409 51901 1443 51935
rect 21281 51901 21315 51935
rect 21465 51901 21499 51935
rect 23121 51901 23155 51935
rect 23305 51901 23339 51935
rect 23397 51901 23431 51935
rect 26801 51901 26835 51935
rect 27997 51901 28031 51935
rect 28181 51901 28215 51935
rect 28273 51901 28307 51935
rect 29101 51901 29135 51935
rect 29561 51901 29595 51935
rect 30021 51901 30055 51935
rect 30277 51901 30311 51935
rect 31953 51901 31987 51935
rect 33425 51901 33459 51935
rect 34345 51901 34379 51935
rect 34612 51901 34646 51935
rect 36185 51901 36219 51935
rect 36369 51901 36403 51935
rect 56609 51901 56643 51935
rect 57437 51901 57471 51935
rect 24216 51833 24250 51867
rect 25789 51833 25823 51867
rect 29193 51833 29227 51867
rect 29285 51833 29319 51867
rect 29423 51833 29457 51867
rect 57989 51833 58023 51867
rect 21097 51765 21131 51799
rect 22937 51765 22971 51799
rect 25329 51765 25363 51799
rect 25994 51765 26028 51799
rect 26157 51765 26191 51799
rect 27813 51765 27847 51799
rect 31401 51765 31435 51799
rect 33517 51765 33551 51799
rect 35725 51765 35759 51799
rect 23673 51561 23707 51595
rect 24225 51561 24259 51595
rect 26801 51561 26835 51595
rect 28641 51561 28675 51595
rect 29101 51561 29135 51595
rect 31125 51561 31159 51595
rect 33425 51561 33459 51595
rect 20720 51493 20754 51527
rect 22560 51493 22594 51527
rect 25688 51493 25722 51527
rect 27528 51493 27562 51527
rect 33977 51493 34011 51527
rect 1409 51425 1443 51459
rect 22293 51425 22327 51459
rect 24133 51425 24167 51459
rect 24317 51425 24351 51459
rect 29285 51425 29319 51459
rect 31033 51425 31067 51459
rect 32312 51425 32346 51459
rect 33885 51425 33919 51459
rect 57989 51425 58023 51459
rect 20453 51357 20487 51391
rect 25421 51357 25455 51391
rect 27261 51357 27295 51391
rect 29561 51357 29595 51391
rect 32045 51357 32079 51391
rect 58173 51289 58207 51323
rect 21833 51221 21867 51255
rect 29469 51221 29503 51255
rect 57437 51221 57471 51255
rect 20913 51017 20947 51051
rect 21557 51017 21591 51051
rect 25053 51017 25087 51051
rect 26157 51017 26191 51051
rect 28273 51017 28307 51051
rect 28917 51017 28951 51051
rect 29561 51017 29595 51051
rect 30573 51017 30607 51051
rect 35817 51017 35851 51051
rect 57989 51017 58023 51051
rect 56885 50949 56919 50983
rect 25605 50881 25639 50915
rect 31769 50881 31803 50915
rect 34621 50881 34655 50915
rect 57529 50881 57563 50915
rect 57713 50881 57747 50915
rect 20821 50813 20855 50847
rect 21005 50813 21039 50847
rect 21465 50813 21499 50847
rect 22845 50813 22879 50847
rect 25234 50813 25268 50847
rect 25697 50813 25731 50847
rect 26157 50813 26191 50847
rect 26433 50813 26467 50847
rect 28181 50813 28215 50847
rect 28825 50813 28859 50847
rect 29009 50813 29043 50847
rect 29469 50813 29503 50847
rect 30481 50813 30515 50847
rect 30665 50813 30699 50847
rect 31585 50813 31619 50847
rect 31861 50813 31895 50847
rect 33057 50813 33091 50847
rect 33241 50813 33275 50847
rect 34345 50813 34379 50847
rect 34529 50813 34563 50847
rect 35081 50813 35115 50847
rect 35265 50813 35299 50847
rect 35725 50813 35759 50847
rect 57069 50813 57103 50847
rect 26341 50745 26375 50779
rect 33149 50745 33183 50779
rect 35173 50745 35207 50779
rect 22661 50677 22695 50711
rect 25237 50677 25271 50711
rect 31401 50677 31435 50711
rect 34161 50677 34195 50711
rect 23949 50473 23983 50507
rect 31861 50473 31895 50507
rect 32321 50473 32355 50507
rect 34805 50473 34839 50507
rect 28917 50405 28951 50439
rect 30748 50405 30782 50439
rect 32689 50405 32723 50439
rect 32827 50405 32861 50439
rect 33692 50405 33726 50439
rect 58173 50405 58207 50439
rect 1409 50337 1443 50371
rect 20361 50337 20395 50371
rect 21456 50337 21490 50371
rect 24133 50337 24167 50371
rect 25789 50337 25823 50371
rect 25973 50337 26007 50371
rect 28089 50337 28123 50371
rect 28825 50337 28859 50371
rect 29009 50337 29043 50371
rect 30481 50337 30515 50371
rect 32505 50337 32539 50371
rect 32597 50337 32631 50371
rect 32965 50337 32999 50371
rect 57253 50337 57287 50371
rect 57989 50337 58023 50371
rect 20637 50269 20671 50303
rect 21189 50269 21223 50303
rect 28365 50269 28399 50303
rect 33425 50269 33459 50303
rect 20177 50133 20211 50167
rect 20545 50133 20579 50167
rect 22569 50133 22603 50167
rect 25789 50133 25823 50167
rect 27905 50133 27939 50167
rect 28273 50133 28307 50167
rect 20821 49929 20855 49963
rect 21373 49929 21407 49963
rect 29193 49929 29227 49963
rect 31125 49929 31159 49963
rect 33149 49929 33183 49963
rect 33701 49929 33735 49963
rect 19441 49793 19475 49827
rect 23581 49793 23615 49827
rect 30113 49793 30147 49827
rect 31769 49793 31803 49827
rect 19708 49725 19742 49759
rect 21281 49725 21315 49759
rect 21465 49725 21499 49759
rect 22569 49725 22603 49759
rect 23848 49725 23882 49759
rect 25513 49725 25547 49759
rect 25780 49725 25814 49759
rect 27813 49725 27847 49759
rect 28069 49725 28103 49759
rect 30021 49725 30055 49759
rect 30205 49725 30239 49759
rect 31033 49725 31067 49759
rect 31677 49725 31711 49759
rect 31861 49725 31895 49759
rect 33057 49725 33091 49759
rect 33885 49725 33919 49759
rect 34529 49725 34563 49759
rect 34713 49725 34747 49759
rect 57437 49725 57471 49759
rect 58173 49725 58207 49759
rect 57989 49657 58023 49691
rect 22661 49589 22695 49623
rect 24961 49589 24995 49623
rect 26893 49589 26927 49623
rect 34621 49589 34655 49623
rect 57253 49589 57287 49623
rect 21465 49385 21499 49419
rect 25237 49385 25271 49419
rect 25421 49385 25455 49419
rect 26709 49385 26743 49419
rect 33517 49385 33551 49419
rect 34805 49385 34839 49419
rect 58173 49385 58207 49419
rect 22477 49317 22511 49351
rect 26341 49317 26375 49351
rect 26546 49317 26580 49351
rect 27712 49317 27746 49351
rect 29377 49317 29411 49351
rect 34463 49317 34497 49351
rect 34653 49317 34687 49351
rect 1409 49249 1443 49283
rect 21649 49249 21683 49283
rect 21833 49249 21867 49283
rect 22385 49249 22419 49283
rect 22569 49249 22603 49283
rect 25362 49249 25396 49283
rect 25881 49249 25915 49283
rect 29285 49249 29319 49283
rect 29469 49249 29503 49283
rect 31300 49249 31334 49283
rect 33514 49249 33548 49283
rect 33977 49249 34011 49283
rect 56885 49249 56919 49283
rect 57713 49249 57747 49283
rect 21925 49181 21959 49215
rect 25789 49181 25823 49215
rect 27445 49181 27479 49215
rect 31033 49181 31067 49215
rect 33885 49181 33919 49215
rect 57529 49181 57563 49215
rect 57069 49113 57103 49147
rect 26525 49045 26559 49079
rect 28825 49045 28859 49079
rect 32413 49045 32447 49079
rect 33333 49045 33367 49079
rect 34621 49045 34655 49079
rect 20453 48841 20487 48875
rect 20637 48841 20671 48875
rect 25513 48841 25547 48875
rect 30481 48841 30515 48875
rect 31309 48841 31343 48875
rect 31953 48841 31987 48875
rect 34437 48841 34471 48875
rect 36277 48841 36311 48875
rect 57437 48841 57471 48875
rect 24961 48705 24995 48739
rect 29101 48705 29135 48739
rect 31401 48705 31435 48739
rect 34897 48705 34931 48739
rect 18153 48637 18187 48671
rect 21097 48637 21131 48671
rect 21281 48637 21315 48671
rect 24869 48637 24903 48671
rect 25697 48637 25731 48671
rect 25789 48637 25823 48671
rect 26709 48637 26743 48671
rect 27813 48637 27847 48671
rect 28457 48637 28491 48671
rect 31125 48637 31159 48671
rect 31861 48637 31895 48671
rect 33057 48637 33091 48671
rect 33324 48637 33358 48671
rect 56609 48637 56643 48671
rect 18420 48569 18454 48603
rect 20269 48569 20303 48603
rect 20485 48569 20519 48603
rect 25513 48569 25547 48603
rect 29368 48569 29402 48603
rect 30941 48569 30975 48603
rect 35142 48569 35176 48603
rect 57989 48569 58023 48603
rect 19533 48501 19567 48535
rect 21189 48501 21223 48535
rect 26801 48501 26835 48535
rect 27905 48501 27939 48535
rect 28549 48501 28583 48535
rect 58081 48501 58115 48535
rect 15209 48297 15243 48331
rect 18429 48297 18463 48331
rect 18613 48297 18647 48331
rect 31309 48297 31343 48331
rect 33701 48297 33735 48331
rect 34437 48297 34471 48331
rect 58173 48297 58207 48331
rect 16221 48229 16255 48263
rect 16437 48229 16471 48263
rect 20812 48229 20846 48263
rect 28641 48229 28675 48263
rect 32321 48229 32355 48263
rect 34253 48229 34287 48263
rect 1409 48161 1443 48195
rect 15206 48161 15240 48195
rect 17049 48161 17083 48195
rect 17233 48161 17267 48195
rect 18610 48161 18644 48195
rect 19073 48161 19107 48195
rect 23673 48161 23707 48195
rect 24133 48161 24167 48195
rect 24317 48161 24351 48195
rect 25605 48161 25639 48195
rect 25872 48161 25906 48195
rect 27905 48161 27939 48195
rect 28825 48161 28859 48195
rect 30481 48161 30515 48195
rect 31493 48161 31527 48195
rect 31677 48161 31711 48195
rect 31769 48161 31803 48195
rect 32229 48161 32263 48195
rect 33057 48161 33091 48195
rect 33609 48161 33643 48195
rect 34529 48161 34563 48195
rect 15577 48093 15611 48127
rect 15669 48093 15703 48127
rect 20545 48093 20579 48127
rect 28181 48093 28215 48127
rect 57069 48093 57103 48127
rect 57529 48093 57563 48127
rect 57713 48093 57747 48127
rect 16589 48025 16623 48059
rect 18981 48025 19015 48059
rect 23489 48025 23523 48059
rect 26985 48025 27019 48059
rect 34253 48025 34287 48059
rect 15025 47957 15059 47991
rect 16405 47957 16439 47991
rect 17049 47957 17083 47991
rect 21925 47957 21959 47991
rect 24225 47957 24259 47991
rect 27721 47957 27755 47991
rect 28089 47957 28123 47991
rect 29009 47957 29043 47991
rect 30573 47957 30607 47991
rect 32873 47957 32907 47991
rect 18705 47753 18739 47787
rect 20177 47753 20211 47787
rect 25329 47753 25363 47787
rect 26341 47753 26375 47787
rect 26801 47753 26835 47787
rect 29929 47753 29963 47787
rect 57253 47753 57287 47787
rect 19257 47617 19291 47651
rect 28273 47617 28307 47651
rect 1409 47549 1443 47583
rect 14381 47549 14415 47583
rect 14648 47549 14682 47583
rect 17325 47549 17359 47583
rect 17581 47549 17615 47583
rect 19165 47549 19199 47583
rect 19349 47549 19383 47583
rect 20361 47549 20395 47583
rect 20453 47549 20487 47583
rect 20913 47549 20947 47583
rect 23949 47549 23983 47583
rect 26525 47549 26559 47583
rect 26617 47549 26651 47583
rect 26893 47549 26927 47583
rect 27813 47549 27847 47583
rect 27905 47549 27939 47583
rect 28089 47549 28123 47583
rect 29745 47549 29779 47583
rect 30021 47549 30055 47583
rect 30665 47549 30699 47583
rect 33333 47549 33367 47583
rect 33517 47549 33551 47583
rect 33609 47549 33643 47583
rect 57437 47549 57471 47583
rect 20177 47481 20211 47515
rect 21005 47481 21039 47515
rect 24216 47481 24250 47515
rect 30932 47481 30966 47515
rect 57989 47481 58023 47515
rect 58173 47481 58207 47515
rect 15761 47413 15795 47447
rect 29561 47413 29595 47447
rect 32045 47413 32079 47447
rect 33149 47413 33183 47447
rect 16313 47209 16347 47243
rect 24225 47209 24259 47243
rect 25237 47209 25271 47243
rect 28273 47209 28307 47243
rect 29561 47209 29595 47243
rect 31033 47209 31067 47243
rect 33701 47209 33735 47243
rect 34253 47209 34287 47243
rect 57713 47209 57747 47243
rect 16129 47141 16163 47175
rect 32588 47141 32622 47175
rect 14933 47073 14967 47107
rect 16405 47073 16439 47107
rect 16865 47073 16899 47107
rect 17049 47073 17083 47107
rect 18797 47073 18831 47107
rect 18981 47073 19015 47107
rect 19993 47073 20027 47107
rect 21180 47073 21214 47107
rect 22937 47073 22971 47107
rect 23673 47073 23707 47107
rect 24133 47073 24167 47107
rect 25421 47073 25455 47107
rect 25697 47073 25731 47107
rect 26801 47073 26835 47107
rect 27813 47073 27847 47107
rect 27997 47073 28031 47107
rect 28273 47073 28307 47107
rect 28457 47073 28491 47107
rect 29377 47073 29411 47107
rect 29561 47073 29595 47107
rect 31217 47073 31251 47107
rect 31493 47073 31527 47107
rect 34161 47073 34195 47107
rect 34345 47073 34379 47107
rect 56885 47073 56919 47107
rect 57529 47073 57563 47107
rect 15209 47005 15243 47039
rect 19073 47005 19107 47039
rect 20913 47005 20947 47039
rect 25605 47005 25639 47039
rect 27077 47005 27111 47039
rect 32321 47005 32355 47039
rect 16129 46937 16163 46971
rect 22753 46937 22787 46971
rect 23489 46937 23523 46971
rect 26985 46937 27019 46971
rect 31401 46937 31435 46971
rect 14749 46869 14783 46903
rect 15117 46869 15151 46903
rect 16957 46869 16991 46903
rect 18613 46869 18647 46903
rect 20085 46869 20119 46903
rect 22293 46869 22327 46903
rect 26617 46869 26651 46903
rect 14841 46665 14875 46699
rect 15393 46665 15427 46699
rect 16037 46665 16071 46699
rect 18981 46665 19015 46699
rect 20821 46665 20855 46699
rect 22753 46665 22787 46699
rect 27813 46665 27847 46699
rect 30297 46665 30331 46699
rect 32045 46665 32079 46699
rect 31217 46597 31251 46631
rect 19441 46529 19475 46563
rect 25513 46529 25547 46563
rect 33057 46529 33091 46563
rect 58173 46529 58207 46563
rect 1409 46461 1443 46495
rect 13461 46461 13495 46495
rect 13728 46461 13762 46495
rect 15301 46461 15335 46495
rect 15485 46461 15519 46495
rect 15945 46461 15979 46495
rect 17601 46461 17635 46495
rect 17868 46461 17902 46495
rect 19708 46461 19742 46495
rect 21465 46461 21499 46495
rect 23397 46461 23431 46495
rect 23581 46461 23615 46495
rect 24777 46461 24811 46495
rect 24961 46461 24995 46495
rect 25053 46461 25087 46495
rect 25780 46461 25814 46495
rect 27813 46461 27847 46495
rect 27997 46461 28031 46495
rect 28917 46461 28951 46495
rect 31493 46461 31527 46495
rect 31953 46461 31987 46495
rect 32137 46461 32171 46495
rect 22569 46393 22603 46427
rect 22785 46393 22819 46427
rect 29184 46393 29218 46427
rect 31217 46393 31251 46427
rect 33324 46393 33358 46427
rect 57989 46393 58023 46427
rect 21557 46325 21591 46359
rect 22937 46325 22971 46359
rect 23489 46325 23523 46359
rect 24593 46325 24627 46359
rect 26893 46325 26927 46359
rect 31401 46325 31435 46359
rect 34437 46325 34471 46359
rect 17141 46121 17175 46155
rect 20637 46121 20671 46155
rect 21465 46121 21499 46155
rect 21649 46121 21683 46155
rect 26617 46121 26651 46155
rect 30481 46121 30515 46155
rect 32505 46121 32539 46155
rect 33517 46121 33551 46155
rect 58173 46121 58207 46155
rect 23020 46053 23054 46087
rect 25482 46053 25516 46087
rect 14749 45985 14783 46019
rect 16028 45985 16062 46019
rect 17601 45985 17635 46019
rect 17785 45985 17819 46019
rect 18521 45985 18555 46019
rect 19993 45985 20027 46019
rect 20177 45985 20211 46019
rect 20821 45985 20855 46019
rect 21646 45985 21680 46019
rect 22109 45985 22143 46019
rect 27077 45985 27111 46019
rect 27261 45985 27295 46019
rect 27721 45985 27755 46019
rect 27977 45985 28011 46019
rect 30665 45985 30699 46019
rect 31392 45985 31426 46019
rect 33425 45985 33459 46019
rect 15761 45917 15795 45951
rect 18061 45917 18095 45951
rect 22017 45917 22051 45951
rect 22753 45917 22787 45951
rect 25237 45917 25271 45951
rect 31125 45917 31159 45951
rect 57069 45917 57103 45951
rect 57529 45917 57563 45951
rect 57713 45917 57747 45951
rect 17969 45849 18003 45883
rect 14841 45781 14875 45815
rect 18613 45781 18647 45815
rect 20085 45781 20119 45815
rect 24133 45781 24167 45815
rect 27169 45781 27203 45815
rect 29101 45781 29135 45815
rect 15393 45577 15427 45611
rect 22569 45577 22603 45611
rect 25145 45577 25179 45611
rect 27813 45577 27847 45611
rect 31493 45577 31527 45611
rect 57253 45577 57287 45611
rect 17785 45509 17819 45543
rect 31677 45509 31711 45543
rect 58173 45509 58207 45543
rect 14013 45441 14047 45475
rect 29285 45441 29319 45475
rect 33149 45441 33183 45475
rect 1409 45373 1443 45407
rect 14280 45373 14314 45407
rect 17601 45373 17635 45407
rect 17877 45373 17911 45407
rect 18613 45373 18647 45407
rect 20913 45373 20947 45407
rect 21097 45373 21131 45407
rect 21189 45373 21223 45407
rect 22569 45373 22603 45407
rect 22845 45373 22879 45407
rect 23305 45373 23339 45407
rect 23489 45373 23523 45407
rect 24409 45373 24443 45407
rect 24593 45373 24627 45407
rect 25053 45373 25087 45407
rect 26065 45373 26099 45407
rect 26249 45373 26283 45407
rect 27813 45373 27847 45407
rect 28089 45373 28123 45407
rect 28641 45373 28675 45407
rect 33057 45373 33091 45407
rect 33241 45373 33275 45407
rect 56609 45373 56643 45407
rect 57437 45373 57471 45407
rect 18858 45305 18892 45339
rect 22753 45305 22787 45339
rect 26433 45305 26467 45339
rect 27997 45305 28031 45339
rect 28733 45305 28767 45339
rect 29552 45305 29586 45339
rect 31309 45305 31343 45339
rect 31514 45305 31548 45339
rect 57989 45305 58023 45339
rect 17417 45237 17451 45271
rect 19993 45237 20027 45271
rect 20729 45237 20763 45271
rect 23397 45237 23431 45271
rect 24501 45237 24535 45271
rect 30665 45237 30699 45271
rect 18153 45033 18187 45067
rect 18613 45033 18647 45067
rect 21649 45033 21683 45067
rect 27905 45033 27939 45067
rect 30481 45033 30515 45067
rect 30665 45033 30699 45067
rect 17040 44965 17074 44999
rect 20536 44965 20570 44999
rect 25596 44965 25630 44999
rect 32045 44965 32079 44999
rect 1409 44897 1443 44931
rect 16773 44897 16807 44931
rect 18797 44897 18831 44931
rect 19073 44897 19107 44931
rect 22753 44897 22787 44931
rect 24041 44897 24075 44931
rect 25329 44897 25363 44931
rect 27169 44897 27203 44931
rect 27813 44897 27847 44931
rect 28641 44897 28675 44931
rect 29101 44897 29135 44931
rect 29285 44897 29319 44931
rect 30662 44897 30696 44931
rect 31125 44897 31159 44931
rect 32229 44897 32263 44931
rect 32321 44897 32355 44931
rect 57253 44897 57287 44931
rect 57989 44897 58023 44931
rect 58173 44897 58207 44931
rect 20269 44829 20303 44863
rect 22937 44829 22971 44863
rect 23029 44829 23063 44863
rect 24317 44829 24351 44863
rect 18981 44761 19015 44795
rect 26709 44761 26743 44795
rect 28457 44761 28491 44795
rect 31033 44761 31067 44795
rect 22569 44693 22603 44727
rect 23857 44693 23891 44727
rect 24225 44693 24259 44727
rect 27261 44693 27295 44727
rect 29101 44693 29135 44727
rect 32045 44693 32079 44727
rect 57437 44693 57471 44727
rect 17785 44489 17819 44523
rect 18613 44489 18647 44523
rect 21097 44489 21131 44523
rect 23949 44489 23983 44523
rect 25789 44489 25823 44523
rect 28457 44489 28491 44523
rect 31953 44489 31987 44523
rect 32137 44489 32171 44523
rect 57989 44489 58023 44523
rect 26893 44421 26927 44455
rect 28135 44421 28169 44455
rect 28273 44421 28307 44455
rect 33057 44421 33091 44455
rect 56885 44421 56919 44455
rect 28365 44353 28399 44387
rect 56425 44353 56459 44387
rect 57529 44353 57563 44387
rect 57713 44353 57747 44387
rect 17693 44285 17727 44319
rect 17877 44285 17911 44319
rect 18521 44285 18555 44319
rect 20361 44285 20395 44319
rect 20453 44285 20487 44319
rect 21005 44285 21039 44319
rect 21189 44285 21223 44319
rect 22569 44285 22603 44319
rect 22825 44285 22859 44319
rect 24409 44285 24443 44319
rect 24665 44285 24699 44319
rect 26525 44285 26559 44319
rect 29285 44285 29319 44319
rect 33057 44285 33091 44319
rect 33241 44285 33275 44319
rect 57069 44285 57103 44319
rect 26709 44217 26743 44251
rect 27997 44217 28031 44251
rect 29530 44217 29564 44251
rect 31769 44217 31803 44251
rect 30665 44149 30699 44183
rect 31974 44149 32008 44183
rect 23765 43945 23799 43979
rect 25237 43945 25271 43979
rect 26157 43945 26191 43979
rect 29469 43945 29503 43979
rect 30573 43945 30607 43979
rect 31585 43945 31619 43979
rect 33977 43945 34011 43979
rect 21097 43877 21131 43911
rect 21302 43877 21336 43911
rect 27537 43877 27571 43911
rect 32864 43877 32898 43911
rect 58173 43877 58207 43911
rect 1409 43809 1443 43843
rect 20453 43809 20487 43843
rect 20637 43809 20671 43843
rect 23673 43809 23707 43843
rect 25421 43809 25455 43843
rect 26341 43809 26375 43843
rect 27445 43809 27479 43843
rect 28089 43809 28123 43843
rect 28181 43809 28215 43843
rect 28365 43809 28399 43843
rect 29285 43809 29319 43843
rect 29561 43809 29595 43843
rect 30481 43809 30515 43843
rect 31582 43809 31616 43843
rect 32597 43809 32631 43843
rect 57989 43809 58023 43843
rect 26617 43741 26651 43775
rect 28549 43741 28583 43775
rect 32045 43741 32079 43775
rect 21465 43673 21499 43707
rect 26525 43673 26559 43707
rect 29285 43673 29319 43707
rect 20453 43605 20487 43639
rect 21281 43605 21315 43639
rect 31401 43605 31435 43639
rect 31953 43605 31987 43639
rect 57437 43605 57471 43639
rect 26341 43401 26375 43435
rect 32045 43401 32079 43435
rect 23121 43333 23155 43367
rect 58173 43333 58207 43367
rect 30665 43265 30699 43299
rect 20177 43197 20211 43231
rect 20444 43197 20478 43231
rect 22750 43197 22784 43231
rect 23213 43197 23247 43231
rect 23765 43197 23799 43231
rect 26065 43197 26099 43231
rect 26157 43197 26191 43231
rect 26433 43197 26467 43231
rect 27813 43197 27847 43231
rect 29653 43197 29687 43231
rect 29837 43197 29871 43231
rect 30932 43197 30966 43231
rect 56609 43197 56643 43231
rect 57437 43197 57471 43231
rect 24032 43129 24066 43163
rect 28058 43129 28092 43163
rect 30021 43129 30055 43163
rect 57989 43129 58023 43163
rect 21557 43061 21591 43095
rect 22569 43061 22603 43095
rect 22753 43061 22787 43095
rect 25145 43061 25179 43095
rect 25881 43061 25915 43095
rect 29193 43061 29227 43095
rect 57253 43061 57287 43095
rect 20453 42857 20487 42891
rect 23305 42857 23339 42891
rect 23970 42857 24004 42891
rect 26617 42857 26651 42891
rect 27169 42857 27203 42891
rect 27997 42857 28031 42891
rect 58173 42857 58207 42891
rect 22192 42789 22226 42823
rect 23765 42789 23799 42823
rect 25504 42789 25538 42823
rect 1409 42721 1443 42755
rect 20450 42721 20484 42755
rect 20913 42721 20947 42755
rect 21925 42721 21959 42755
rect 25237 42721 25271 42755
rect 27077 42721 27111 42755
rect 28181 42721 28215 42755
rect 28365 42721 28399 42755
rect 29193 42721 29227 42755
rect 29377 42721 29411 42755
rect 30481 42721 30515 42755
rect 31309 42721 31343 42755
rect 31953 42721 31987 42755
rect 32505 42721 32539 42755
rect 32689 42721 32723 42755
rect 56885 42721 56919 42755
rect 57069 42721 57103 42755
rect 57529 42721 57563 42755
rect 57713 42721 57747 42755
rect 20821 42653 20855 42687
rect 28457 42653 28491 42687
rect 20269 42517 20303 42551
rect 23949 42517 23983 42551
rect 24133 42517 24167 42551
rect 29561 42517 29595 42551
rect 30573 42517 30607 42551
rect 31125 42517 31159 42551
rect 31769 42517 31803 42551
rect 32505 42517 32539 42551
rect 21373 42313 21407 42347
rect 24317 42313 24351 42347
rect 25881 42313 25915 42347
rect 26617 42313 26651 42347
rect 28070 42313 28104 42347
rect 30481 42313 30515 42347
rect 23581 42245 23615 42279
rect 28181 42245 28215 42279
rect 28273 42177 28307 42211
rect 32045 42177 32079 42211
rect 33057 42177 33091 42211
rect 1409 42109 1443 42143
rect 19533 42109 19567 42143
rect 19800 42109 19834 42143
rect 21373 42109 21407 42143
rect 21649 42109 21683 42143
rect 23765 42109 23799 42143
rect 23857 42109 23891 42143
rect 24317 42109 24351 42143
rect 24501 42109 24535 42143
rect 24961 42109 24995 42143
rect 26065 42109 26099 42143
rect 26525 42109 26559 42143
rect 28641 42109 28675 42143
rect 29101 42109 29135 42143
rect 29368 42109 29402 42143
rect 31674 42109 31708 42143
rect 32137 42109 32171 42143
rect 33313 42109 33347 42143
rect 56609 42109 56643 42143
rect 57437 42109 57471 42143
rect 23581 42041 23615 42075
rect 27905 42041 27939 42075
rect 57989 42041 58023 42075
rect 58173 42041 58207 42075
rect 20913 41973 20947 42007
rect 21557 41973 21591 42007
rect 25053 41973 25087 42007
rect 31493 41973 31527 42007
rect 31677 41973 31711 42007
rect 34437 41973 34471 42007
rect 20913 41769 20947 41803
rect 27721 41769 27755 41803
rect 32045 41769 32079 41803
rect 33517 41769 33551 41803
rect 58173 41769 58207 41803
rect 30932 41701 30966 41735
rect 32505 41701 32539 41735
rect 32710 41701 32744 41735
rect 33333 41701 33367 41735
rect 20821 41633 20855 41667
rect 21721 41633 21755 41667
rect 23857 41633 23891 41667
rect 24041 41633 24075 41667
rect 25513 41633 25547 41667
rect 25697 41633 25731 41667
rect 26341 41633 26375 41667
rect 26608 41633 26642 41667
rect 28181 41633 28215 41667
rect 28457 41633 28491 41667
rect 29377 41633 29411 41667
rect 30665 41633 30699 41667
rect 33609 41633 33643 41667
rect 57069 41633 57103 41667
rect 57529 41633 57563 41667
rect 21465 41565 21499 41599
rect 24133 41565 24167 41599
rect 25789 41565 25823 41599
rect 28917 41565 28951 41599
rect 29469 41565 29503 41599
rect 57713 41565 57747 41599
rect 28273 41497 28307 41531
rect 32873 41497 32907 41531
rect 33333 41497 33367 41531
rect 56885 41497 56919 41531
rect 22845 41429 22879 41463
rect 23673 41429 23707 41463
rect 25329 41429 25363 41463
rect 32689 41429 32723 41463
rect 21189 41225 21223 41259
rect 24501 41225 24535 41259
rect 26341 41225 26375 41259
rect 27813 41225 27847 41259
rect 30665 41225 30699 41259
rect 57345 41225 57379 41259
rect 23121 41089 23155 41123
rect 28825 41089 28859 41123
rect 31033 41089 31067 41123
rect 1409 41021 1443 41055
rect 21373 41021 21407 41055
rect 21557 41021 21591 41055
rect 21649 41021 21683 41055
rect 23388 41021 23422 41055
rect 24961 41021 24995 41055
rect 25228 41021 25262 41055
rect 28089 41021 28123 41055
rect 30849 41021 30883 41055
rect 31125 41021 31159 41055
rect 31861 41021 31895 41055
rect 33057 41021 33091 41055
rect 33241 41021 33275 41055
rect 56517 41021 56551 41055
rect 27813 40953 27847 40987
rect 27997 40953 28031 40987
rect 29070 40953 29104 40987
rect 57253 40953 57287 40987
rect 57989 40953 58023 40987
rect 58173 40953 58207 40987
rect 30205 40885 30239 40919
rect 31953 40885 31987 40919
rect 33149 40885 33183 40919
rect 21649 40681 21683 40715
rect 22293 40681 22327 40715
rect 24225 40681 24259 40715
rect 29009 40681 29043 40715
rect 32597 40681 32631 40715
rect 58173 40681 58207 40715
rect 20085 40613 20119 40647
rect 33517 40613 33551 40647
rect 15117 40545 15151 40579
rect 15301 40545 15335 40579
rect 18797 40545 18831 40579
rect 18981 40545 19015 40579
rect 19993 40545 20027 40579
rect 20177 40545 20211 40579
rect 20821 40545 20855 40579
rect 21557 40545 21591 40579
rect 22201 40545 22235 40579
rect 22385 40545 22419 40579
rect 24041 40545 24075 40579
rect 24225 40545 24259 40579
rect 25697 40545 25731 40579
rect 25881 40545 25915 40579
rect 26893 40545 26927 40579
rect 27077 40545 27111 40579
rect 27721 40545 27755 40579
rect 29193 40545 29227 40579
rect 29285 40545 29319 40579
rect 29561 40545 29595 40579
rect 30481 40545 30515 40579
rect 31493 40545 31527 40579
rect 31585 40545 31619 40579
rect 31861 40545 31895 40579
rect 32781 40545 32815 40579
rect 33701 40545 33735 40579
rect 57069 40545 57103 40579
rect 19073 40477 19107 40511
rect 21097 40477 21131 40511
rect 27997 40477 28031 40511
rect 30573 40477 30607 40511
rect 33057 40477 33091 40511
rect 57529 40477 57563 40511
rect 57713 40477 57747 40511
rect 25697 40409 25731 40443
rect 26893 40409 26927 40443
rect 27905 40409 27939 40443
rect 29469 40409 29503 40443
rect 56885 40409 56919 40443
rect 15117 40341 15151 40375
rect 18613 40341 18647 40375
rect 20637 40341 20671 40375
rect 21005 40341 21039 40375
rect 27537 40341 27571 40375
rect 31309 40341 31343 40375
rect 31769 40341 31803 40375
rect 32965 40341 32999 40375
rect 33885 40341 33919 40375
rect 19717 40137 19751 40171
rect 21557 40137 21591 40171
rect 29745 40137 29779 40171
rect 31861 40137 31895 40171
rect 57437 40137 57471 40171
rect 14749 40069 14783 40103
rect 15853 40001 15887 40035
rect 34989 40001 35023 40035
rect 1409 39933 1443 39967
rect 12449 39933 12483 39967
rect 12633 39933 12667 39967
rect 12725 39933 12759 39967
rect 13369 39933 13403 39967
rect 15347 39933 15381 39967
rect 15761 39933 15795 39967
rect 18337 39933 18371 39967
rect 18604 39933 18638 39967
rect 20177 39933 20211 39967
rect 20444 39933 20478 39967
rect 25973 39933 26007 39967
rect 27813 39933 27847 39967
rect 29653 39933 29687 39967
rect 30481 39933 30515 39967
rect 30748 39933 30782 39967
rect 33057 39933 33091 39967
rect 33313 39933 33347 39967
rect 34897 39933 34931 39967
rect 57989 39933 58023 39967
rect 13636 39865 13670 39899
rect 28058 39865 28092 39899
rect 58173 39865 58207 39899
rect 12265 39797 12299 39831
rect 15209 39797 15243 39831
rect 15393 39797 15427 39831
rect 26065 39797 26099 39831
rect 29193 39797 29227 39831
rect 34437 39797 34471 39831
rect 12909 39593 12943 39627
rect 13461 39593 13495 39627
rect 17325 39593 17359 39627
rect 20913 39593 20947 39627
rect 26893 39593 26927 39627
rect 28181 39593 28215 39627
rect 31309 39593 31343 39627
rect 33057 39593 33091 39627
rect 11796 39525 11830 39559
rect 15454 39525 15488 39559
rect 25780 39525 25814 39559
rect 11529 39457 11563 39491
rect 13369 39457 13403 39491
rect 13553 39457 13587 39491
rect 17509 39457 17543 39491
rect 20177 39457 20211 39491
rect 20269 39457 20303 39491
rect 20821 39457 20855 39491
rect 21005 39457 21039 39491
rect 27353 39457 27387 39491
rect 28089 39457 28123 39491
rect 31217 39457 31251 39491
rect 31861 39457 31895 39491
rect 32597 39457 32631 39491
rect 32781 39457 32815 39491
rect 33057 39457 33091 39491
rect 33149 39457 33183 39491
rect 57989 39457 58023 39491
rect 15209 39389 15243 39423
rect 25513 39389 25547 39423
rect 31953 39389 31987 39423
rect 16589 39253 16623 39287
rect 27445 39253 27479 39287
rect 13461 39049 13495 39083
rect 14933 39049 14967 39083
rect 15577 39049 15611 39083
rect 20545 39049 20579 39083
rect 15117 38981 15151 39015
rect 25881 38981 25915 39015
rect 26709 38981 26743 39015
rect 32045 38981 32079 39015
rect 33057 38981 33091 39015
rect 17693 38913 17727 38947
rect 26801 38913 26835 38947
rect 32137 38913 32171 38947
rect 1409 38845 1443 38879
rect 12449 38845 12483 38879
rect 13369 38845 13403 38879
rect 15577 38845 15611 38879
rect 15761 38845 15795 38879
rect 15853 38845 15887 38879
rect 19717 38845 19751 38879
rect 19901 38845 19935 38879
rect 19993 38845 20027 38879
rect 20453 38845 20487 38879
rect 24501 38845 24535 38879
rect 26525 38845 26559 38879
rect 28365 38845 28399 38879
rect 31861 38845 31895 38879
rect 33057 38845 33091 38879
rect 33241 38845 33275 38879
rect 33701 38845 33735 38879
rect 14749 38777 14783 38811
rect 14965 38777 14999 38811
rect 17960 38777 17994 38811
rect 24768 38777 24802 38811
rect 26341 38777 26375 38811
rect 28632 38777 28666 38811
rect 33968 38777 34002 38811
rect 57989 38777 58023 38811
rect 58173 38777 58207 38811
rect 12541 38709 12575 38743
rect 19073 38709 19107 38743
rect 19533 38709 19567 38743
rect 29745 38709 29779 38743
rect 31677 38709 31711 38743
rect 35081 38709 35115 38743
rect 13277 38505 13311 38539
rect 17325 38505 17359 38539
rect 18981 38505 19015 38539
rect 21373 38505 21407 38539
rect 26065 38505 26099 38539
rect 27905 38505 27939 38539
rect 29377 38505 29411 38539
rect 32321 38505 32355 38539
rect 33241 38505 33275 38539
rect 58173 38505 58207 38539
rect 12164 38437 12198 38471
rect 18061 38437 18095 38471
rect 18277 38437 18311 38471
rect 20238 38437 20272 38471
rect 28365 38437 28399 38471
rect 28581 38437 28615 38471
rect 29193 38437 29227 38471
rect 31208 38437 31242 38471
rect 33977 38437 34011 38471
rect 1409 38369 1443 38403
rect 11897 38369 11931 38403
rect 14933 38369 14967 38403
rect 15945 38369 15979 38403
rect 16212 38369 16246 38403
rect 18889 38369 18923 38403
rect 19073 38369 19107 38403
rect 19993 38369 20027 38403
rect 25881 38369 25915 38403
rect 26065 38369 26099 38403
rect 26792 38369 26826 38403
rect 29469 38369 29503 38403
rect 30941 38369 30975 38403
rect 32781 38369 32815 38403
rect 32873 38369 32907 38403
rect 33057 38369 33091 38403
rect 34161 38369 34195 38403
rect 34253 38369 34287 38403
rect 15209 38301 15243 38335
rect 26525 38301 26559 38335
rect 57069 38301 57103 38335
rect 57529 38301 57563 38335
rect 57713 38301 57747 38335
rect 18429 38233 18463 38267
rect 33977 38233 34011 38267
rect 14749 38165 14783 38199
rect 15117 38165 15151 38199
rect 18245 38165 18279 38199
rect 28549 38165 28583 38199
rect 28733 38165 28767 38199
rect 29193 38165 29227 38199
rect 15117 37961 15151 37995
rect 15669 37961 15703 37995
rect 17325 37961 17359 37995
rect 18429 37961 18463 37995
rect 27813 37961 27847 37995
rect 28365 37961 28399 37995
rect 28917 37961 28951 37995
rect 35173 37961 35207 37995
rect 57253 37961 57287 37995
rect 17877 37893 17911 37927
rect 58173 37893 58207 37927
rect 17969 37825 18003 37859
rect 28457 37825 28491 37859
rect 13737 37757 13771 37791
rect 14004 37757 14038 37791
rect 15577 37757 15611 37791
rect 15761 37757 15795 37791
rect 16405 37757 16439 37791
rect 17506 37757 17540 37791
rect 18429 37757 18463 37791
rect 18613 37757 18647 37791
rect 18705 37757 18739 37791
rect 27994 37757 28028 37791
rect 28917 37757 28951 37791
rect 29101 37757 29135 37791
rect 33333 37757 33367 37791
rect 34437 37757 34471 37791
rect 35081 37757 35115 37791
rect 56609 37757 56643 37791
rect 57437 37757 57471 37791
rect 19717 37689 19751 37723
rect 33149 37689 33183 37723
rect 33517 37689 33551 37723
rect 57989 37689 58023 37723
rect 16221 37621 16255 37655
rect 17509 37621 17543 37655
rect 21005 37621 21039 37655
rect 27997 37621 28031 37655
rect 34529 37621 34563 37655
rect 18797 37417 18831 37451
rect 20177 37417 20211 37451
rect 20637 37417 20671 37451
rect 34805 37417 34839 37451
rect 58081 37417 58115 37451
rect 15761 37349 15795 37383
rect 18153 37349 18187 37383
rect 28457 37349 28491 37383
rect 33670 37349 33704 37383
rect 1409 37281 1443 37315
rect 14933 37281 14967 37315
rect 15117 37281 15151 37315
rect 15669 37281 15703 37315
rect 16313 37281 16347 37315
rect 16405 37281 16439 37315
rect 16957 37281 16991 37315
rect 17141 37281 17175 37315
rect 18061 37281 18095 37315
rect 18245 37281 18279 37315
rect 18705 37281 18739 37315
rect 19993 37281 20027 37315
rect 20177 37281 20211 37315
rect 20821 37281 20855 37315
rect 28365 37281 28399 37315
rect 28549 37281 28583 37315
rect 29009 37281 29043 37315
rect 29101 37281 29135 37315
rect 30481 37281 30515 37315
rect 30665 37281 30699 37315
rect 31125 37281 31159 37315
rect 31392 37281 31426 37315
rect 33425 37281 33459 37315
rect 57253 37281 57287 37315
rect 57989 37281 58023 37315
rect 15209 37213 15243 37247
rect 14749 37077 14783 37111
rect 17049 37077 17083 37111
rect 30573 37077 30607 37111
rect 32505 37077 32539 37111
rect 57437 37077 57471 37111
rect 15301 36873 15335 36907
rect 15853 36873 15887 36907
rect 18981 36873 19015 36907
rect 28273 36873 28307 36907
rect 31217 36873 31251 36907
rect 57989 36873 58023 36907
rect 30389 36805 30423 36839
rect 33241 36805 33275 36839
rect 17601 36737 17635 36771
rect 31309 36737 31343 36771
rect 13921 36669 13955 36703
rect 14188 36669 14222 36703
rect 15761 36669 15795 36703
rect 15945 36669 15979 36703
rect 28089 36669 28123 36703
rect 28365 36669 28399 36703
rect 29009 36669 29043 36703
rect 31033 36669 31067 36703
rect 31953 36669 31987 36703
rect 33149 36669 33183 36703
rect 33425 36669 33459 36703
rect 56333 36669 56367 36703
rect 57529 36669 57563 36703
rect 57713 36669 57747 36703
rect 17868 36601 17902 36635
rect 29276 36601 29310 36635
rect 30849 36601 30883 36635
rect 56885 36601 56919 36635
rect 57069 36601 57103 36635
rect 27905 36533 27939 36567
rect 32045 36533 32079 36567
rect 33609 36533 33643 36567
rect 17049 36329 17083 36363
rect 18429 36329 18463 36363
rect 28641 36329 28675 36363
rect 32229 36329 32263 36363
rect 33241 36329 33275 36363
rect 57253 36329 57287 36363
rect 27528 36261 27562 36295
rect 1409 36193 1443 36227
rect 15669 36193 15703 36227
rect 15936 36193 15970 36227
rect 17509 36193 17543 36227
rect 17693 36193 17727 36227
rect 17969 36193 18003 36227
rect 18613 36193 18647 36227
rect 18889 36193 18923 36227
rect 30481 36193 30515 36227
rect 32413 36193 32447 36227
rect 32505 36193 32539 36227
rect 32781 36193 32815 36227
rect 33425 36193 33459 36227
rect 34161 36193 34195 36227
rect 57437 36193 57471 36227
rect 57989 36193 58023 36227
rect 17877 36125 17911 36159
rect 27261 36125 27295 36159
rect 33701 36125 33735 36159
rect 34253 36057 34287 36091
rect 18797 35989 18831 36023
rect 30573 35989 30607 36023
rect 32689 35989 32723 36023
rect 33609 35989 33643 36023
rect 58081 35989 58115 36023
rect 17601 35785 17635 35819
rect 31125 35785 31159 35819
rect 57989 35785 58023 35819
rect 18153 35717 18187 35751
rect 33149 35649 33183 35683
rect 1409 35581 1443 35615
rect 17509 35581 17543 35615
rect 18337 35581 18371 35615
rect 30941 35581 30975 35615
rect 31217 35581 31251 35615
rect 31677 35581 31711 35615
rect 31861 35581 31895 35615
rect 34989 35581 35023 35615
rect 35173 35581 35207 35615
rect 56241 35581 56275 35615
rect 57069 35581 57103 35615
rect 57529 35581 57563 35615
rect 57713 35581 57747 35615
rect 33416 35513 33450 35547
rect 35081 35513 35115 35547
rect 30757 35445 30791 35479
rect 31769 35445 31803 35479
rect 34529 35445 34563 35479
rect 31861 35241 31895 35275
rect 32321 35241 32355 35275
rect 57253 35241 57287 35275
rect 30748 35173 30782 35207
rect 20177 35105 20211 35139
rect 32505 35105 32539 35139
rect 32689 35105 32723 35139
rect 33241 35105 33275 35139
rect 33517 35105 33551 35139
rect 34437 35105 34471 35139
rect 57437 35105 57471 35139
rect 57989 35105 58023 35139
rect 30481 35037 30515 35071
rect 32781 35037 32815 35071
rect 33701 35037 33735 35071
rect 33333 34969 33367 35003
rect 34529 34969 34563 35003
rect 58173 34969 58207 35003
rect 19993 34901 20027 34935
rect 17693 34697 17727 34731
rect 22569 34697 22603 34731
rect 33517 34697 33551 34731
rect 34805 34629 34839 34663
rect 31861 34561 31895 34595
rect 56149 34561 56183 34595
rect 1409 34493 1443 34527
rect 17877 34493 17911 34527
rect 22753 34493 22787 34527
rect 31033 34493 31067 34527
rect 31217 34493 31251 34527
rect 31309 34493 31343 34527
rect 31769 34493 31803 34527
rect 33241 34493 33275 34527
rect 33333 34493 33367 34527
rect 33609 34493 33643 34527
rect 34069 34493 34103 34527
rect 34253 34493 34287 34527
rect 34713 34493 34747 34527
rect 55321 34493 55355 34527
rect 56793 34493 56827 34527
rect 57437 34493 57471 34527
rect 58173 34493 58207 34527
rect 57989 34425 58023 34459
rect 30849 34357 30883 34391
rect 33057 34357 33091 34391
rect 34161 34357 34195 34391
rect 57253 34357 57287 34391
rect 22385 34153 22419 34187
rect 31861 34153 31895 34187
rect 33701 34153 33735 34187
rect 58173 34153 58207 34187
rect 30748 34085 30782 34119
rect 32588 34085 32622 34119
rect 34253 34085 34287 34119
rect 21261 34017 21295 34051
rect 23029 34017 23063 34051
rect 23397 34017 23431 34051
rect 34161 34017 34195 34051
rect 35725 34017 35759 34051
rect 54953 34017 54987 34051
rect 55781 34017 55815 34051
rect 57069 34017 57103 34051
rect 57529 34017 57563 34051
rect 21005 33949 21039 33983
rect 23121 33949 23155 33983
rect 30481 33949 30515 33983
rect 32321 33949 32355 33983
rect 57713 33949 57747 33983
rect 23029 33881 23063 33915
rect 56885 33881 56919 33915
rect 35817 33813 35851 33847
rect 55597 33813 55631 33847
rect 20637 33609 20671 33643
rect 22753 33609 22787 33643
rect 54125 33609 54159 33643
rect 31309 33541 31343 33575
rect 33057 33541 33091 33575
rect 35357 33541 35391 33575
rect 26065 33473 26099 33507
rect 54401 33473 54435 33507
rect 55045 33473 55079 33507
rect 57069 33473 57103 33507
rect 57713 33473 57747 33507
rect 1409 33405 1443 33439
rect 20637 33405 20671 33439
rect 20821 33405 20855 33439
rect 21281 33405 21315 33439
rect 22661 33405 22695 33439
rect 23489 33405 23523 33439
rect 25329 33405 25363 33439
rect 25789 33405 25823 33439
rect 31217 33405 31251 33439
rect 31401 33405 31435 33439
rect 33057 33405 33091 33439
rect 33241 33405 33275 33439
rect 33977 33405 34011 33439
rect 34244 33405 34278 33439
rect 35817 33405 35851 33439
rect 36001 33405 36035 33439
rect 56333 33405 56367 33439
rect 57529 33405 57563 33439
rect 23756 33337 23790 33371
rect 54493 33337 54527 33371
rect 55689 33337 55723 33371
rect 55781 33337 55815 33371
rect 56885 33337 56919 33371
rect 21373 33269 21407 33303
rect 24869 33269 24903 33303
rect 36185 33269 36219 33303
rect 58173 33269 58207 33303
rect 21373 33065 21407 33099
rect 23397 33065 23431 33099
rect 23949 33065 23983 33099
rect 33333 33065 33367 33099
rect 35725 33065 35759 33099
rect 53665 33065 53699 33099
rect 55781 33065 55815 33099
rect 23029 32997 23063 33031
rect 31585 32997 31619 33031
rect 34069 32997 34103 33031
rect 54493 32997 54527 33031
rect 57345 32997 57379 33031
rect 57897 32997 57931 33031
rect 1409 32929 1443 32963
rect 20260 32929 20294 32963
rect 22017 32929 22051 32963
rect 22109 32929 22143 32963
rect 22385 32929 22419 32963
rect 22845 32929 22879 32963
rect 23121 32929 23155 32963
rect 23213 32929 23247 32963
rect 23857 32929 23891 32963
rect 24041 32929 24075 32963
rect 25237 32929 25271 32963
rect 25789 32929 25823 32963
rect 31769 32929 31803 32963
rect 31861 32929 31895 32963
rect 32873 32929 32907 32963
rect 33119 32929 33153 32963
rect 34216 32929 34250 32963
rect 35909 32929 35943 32963
rect 36093 32929 36127 32963
rect 53849 32929 53883 32963
rect 55597 32929 55631 32963
rect 19993 32861 20027 32895
rect 25973 32861 26007 32895
rect 34437 32861 34471 32895
rect 36185 32861 36219 32895
rect 54401 32861 54435 32895
rect 57253 32861 57287 32895
rect 32965 32793 32999 32827
rect 34345 32793 34379 32827
rect 54953 32793 54987 32827
rect 21833 32725 21867 32759
rect 22293 32725 22327 32759
rect 31585 32725 31619 32759
rect 34529 32725 34563 32759
rect 54401 32521 54435 32555
rect 23489 32453 23523 32487
rect 33149 32453 33183 32487
rect 55965 32453 55999 32487
rect 58173 32453 58207 32487
rect 13737 32385 13771 32419
rect 25697 32385 25731 32419
rect 30573 32385 30607 32419
rect 56241 32385 56275 32419
rect 57161 32385 57195 32419
rect 13369 32317 13403 32351
rect 14657 32317 14691 32351
rect 14841 32317 14875 32351
rect 15485 32317 15519 32351
rect 17969 32317 18003 32351
rect 18153 32317 18187 32351
rect 19441 32317 19475 32351
rect 20809 32317 20843 32351
rect 21005 32317 21039 32351
rect 21465 32317 21499 32351
rect 22937 32317 22971 32351
rect 23305 32317 23339 32351
rect 23949 32317 23983 32351
rect 24961 32317 24995 32351
rect 25421 32317 25455 32351
rect 26157 32317 26191 32351
rect 30840 32317 30874 32351
rect 33057 32317 33091 32351
rect 33885 32317 33919 32351
rect 54585 32317 54619 32351
rect 55505 32317 55539 32351
rect 57989 32317 58023 32351
rect 13185 32249 13219 32283
rect 23121 32249 23155 32283
rect 23213 32249 23247 32283
rect 24041 32249 24075 32283
rect 34152 32249 34186 32283
rect 56333 32249 56367 32283
rect 14749 32181 14783 32215
rect 15301 32181 15335 32215
rect 18061 32181 18095 32215
rect 19533 32181 19567 32215
rect 20913 32181 20947 32215
rect 21557 32181 21591 32215
rect 26249 32181 26283 32215
rect 31953 32181 31987 32215
rect 35265 32181 35299 32215
rect 55689 32181 55723 32215
rect 16865 31977 16899 32011
rect 19073 31977 19107 32011
rect 21189 31977 21223 32011
rect 32045 31977 32079 32011
rect 34253 31977 34287 32011
rect 12449 31909 12483 31943
rect 17960 31909 17994 31943
rect 20729 31909 20763 31943
rect 22293 31909 22327 31943
rect 26525 31909 26559 31943
rect 55137 31909 55171 31943
rect 55229 31909 55263 31943
rect 55781 31909 55815 31943
rect 57621 31909 57655 31943
rect 58173 31909 58207 31943
rect 1409 31841 1443 31875
rect 13645 31841 13679 31875
rect 14933 31841 14967 31875
rect 15117 31841 15151 31875
rect 15577 31841 15611 31875
rect 15761 31841 15795 31875
rect 16221 31841 16255 31875
rect 16405 31841 16439 31875
rect 17049 31841 17083 31875
rect 19993 31841 20027 31875
rect 20453 31841 20487 31875
rect 21465 31841 21499 31875
rect 21557 31841 21591 31875
rect 21649 31841 21683 31875
rect 21833 31841 21867 31875
rect 22477 31841 22511 31875
rect 23121 31841 23155 31875
rect 23305 31841 23339 31875
rect 25237 31841 25271 31875
rect 25697 31841 25731 31875
rect 26433 31841 26467 31875
rect 27344 31841 27378 31875
rect 32045 31841 32079 31875
rect 32137 31841 32171 31875
rect 32404 31841 32438 31875
rect 34437 31841 34471 31875
rect 34529 31841 34563 31875
rect 34805 31841 34839 31875
rect 35725 31841 35759 31875
rect 53941 31841 53975 31875
rect 54585 31841 54619 31875
rect 56793 31841 56827 31875
rect 56977 31841 57011 31875
rect 12596 31773 12630 31807
rect 12817 31773 12851 31807
rect 15669 31773 15703 31807
rect 16313 31773 16347 31807
rect 17693 31773 17727 31807
rect 22661 31773 22695 31807
rect 25973 31773 26007 31807
rect 27077 31773 27111 31807
rect 34713 31773 34747 31807
rect 35817 31773 35851 31807
rect 57345 31773 57379 31807
rect 57529 31773 57563 31807
rect 13829 31705 13863 31739
rect 53757 31705 53791 31739
rect 54401 31705 54435 31739
rect 12725 31637 12759 31671
rect 13093 31637 13127 31671
rect 14933 31637 14967 31671
rect 23121 31637 23155 31671
rect 28457 31637 28491 31671
rect 33517 31637 33551 31671
rect 12725 31433 12759 31467
rect 19533 31433 19567 31467
rect 21649 31433 21683 31467
rect 27813 31433 27847 31467
rect 33057 31433 33091 31467
rect 33425 31433 33459 31467
rect 34069 31433 34103 31467
rect 34713 31433 34747 31467
rect 12614 31365 12648 31399
rect 13737 31365 13771 31399
rect 12817 31297 12851 31331
rect 15761 31297 15795 31331
rect 20177 31297 20211 31331
rect 23029 31297 23063 31331
rect 23581 31297 23615 31331
rect 24133 31297 24167 31331
rect 25145 31297 25179 31331
rect 33517 31297 33551 31331
rect 58173 31297 58207 31331
rect 12449 31229 12483 31263
rect 13645 31229 13679 31263
rect 14473 31229 14507 31263
rect 15485 31229 15519 31263
rect 17877 31229 17911 31263
rect 17969 31229 18003 31263
rect 18061 31229 18095 31263
rect 18245 31229 18279 31263
rect 19257 31229 19291 31263
rect 19349 31229 19383 31263
rect 19625 31229 19659 31263
rect 20085 31229 20119 31263
rect 21005 31229 21039 31263
rect 21153 31229 21187 31263
rect 21373 31229 21407 31263
rect 21470 31229 21504 31263
rect 22569 31229 22603 31263
rect 22753 31229 22787 31263
rect 22845 31229 22879 31263
rect 23121 31229 23155 31263
rect 23765 31229 23799 31263
rect 27813 31229 27847 31263
rect 27997 31229 28031 31263
rect 33241 31229 33275 31263
rect 33977 31229 34011 31263
rect 34621 31229 34655 31263
rect 52929 31229 52963 31263
rect 55597 31229 55631 31263
rect 56241 31229 56275 31263
rect 13185 31161 13219 31195
rect 21281 31161 21315 31195
rect 24041 31161 24075 31195
rect 25412 31161 25446 31195
rect 54493 31161 54527 31195
rect 54585 31161 54619 31195
rect 55137 31161 55171 31195
rect 57161 31161 57195 31195
rect 57253 31161 57287 31195
rect 14565 31093 14599 31127
rect 17601 31093 17635 31127
rect 19073 31093 19107 31127
rect 23949 31093 23983 31127
rect 26525 31093 26559 31127
rect 55781 31093 55815 31127
rect 56425 31093 56459 31127
rect 56885 31093 56919 31127
rect 13645 30889 13679 30923
rect 15393 30889 15427 30923
rect 18429 30889 18463 30923
rect 21373 30889 21407 30923
rect 21925 30889 21959 30923
rect 25973 30889 26007 30923
rect 28825 30889 28859 30923
rect 54309 30889 54343 30923
rect 54953 30889 54987 30923
rect 12449 30821 12483 30855
rect 16212 30821 16246 30855
rect 18061 30821 18095 30855
rect 18981 30821 19015 30855
rect 56885 30821 56919 30855
rect 57805 30821 57839 30855
rect 1409 30753 1443 30787
rect 10517 30753 10551 30787
rect 10977 30753 11011 30787
rect 11161 30753 11195 30787
rect 11805 30753 11839 30787
rect 13829 30753 13863 30787
rect 15209 30753 15243 30787
rect 15301 30753 15335 30787
rect 17785 30753 17819 30787
rect 17933 30753 17967 30787
rect 18153 30753 18187 30787
rect 18291 30753 18325 30787
rect 18889 30753 18923 30787
rect 19993 30753 20027 30787
rect 20260 30753 20294 30787
rect 21833 30753 21867 30787
rect 23029 30753 23063 30787
rect 23213 30753 23247 30787
rect 23305 30753 23339 30787
rect 23581 30753 23615 30787
rect 25237 30753 25271 30787
rect 25421 30753 25455 30787
rect 25516 30753 25550 30787
rect 25789 30753 25823 30787
rect 26617 30753 26651 30787
rect 26709 30753 26743 30787
rect 26985 30753 27019 30787
rect 27712 30753 27746 30787
rect 29285 30753 29319 30787
rect 54493 30753 54527 30787
rect 55137 30753 55171 30787
rect 55597 30753 55631 30787
rect 11897 30685 11931 30719
rect 12817 30685 12851 30719
rect 12725 30617 12759 30651
rect 15945 30685 15979 30719
rect 23397 30685 23431 30719
rect 25605 30685 25639 30719
rect 27445 30685 27479 30719
rect 56793 30685 56827 30719
rect 53849 30617 53883 30651
rect 55781 30617 55815 30651
rect 10333 30549 10367 30583
rect 10977 30549 11011 30583
rect 12614 30549 12648 30583
rect 13093 30549 13127 30583
rect 15209 30549 15243 30583
rect 17325 30549 17359 30583
rect 23765 30549 23799 30583
rect 26433 30549 26467 30583
rect 26893 30549 26927 30583
rect 29377 30549 29411 30583
rect 56609 30549 56643 30583
rect 10333 30345 10367 30379
rect 12725 30345 12759 30379
rect 13829 30345 13863 30379
rect 18337 30345 18371 30379
rect 20177 30345 20211 30379
rect 25513 30345 25547 30379
rect 28457 30345 28491 30379
rect 31125 30345 31159 30379
rect 12587 30277 12621 30311
rect 16037 30277 16071 30311
rect 17785 30277 17819 30311
rect 20729 30277 20763 30311
rect 21465 30277 21499 30311
rect 24869 30277 24903 30311
rect 25973 30277 26007 30311
rect 26709 30277 26743 30311
rect 12817 30209 12851 30243
rect 14105 30209 14139 30243
rect 16238 30209 16272 30243
rect 17877 30209 17911 30243
rect 18797 30209 18831 30243
rect 19717 30209 19751 30243
rect 19809 30209 19843 30243
rect 1409 30141 1443 30175
rect 9689 30141 9723 30175
rect 10517 30141 10551 30175
rect 10977 30141 11011 30175
rect 12449 30141 12483 30175
rect 13645 30141 13679 30175
rect 15117 30141 15151 30175
rect 15945 30141 15979 30175
rect 16129 30141 16163 30175
rect 16405 30141 16439 30175
rect 17325 30141 17359 30175
rect 17509 30141 17543 30175
rect 18521 30141 18555 30175
rect 18613 30141 18647 30175
rect 18889 30141 18923 30175
rect 19441 30141 19475 30175
rect 19625 30141 19659 30175
rect 19993 30141 20027 30175
rect 20637 30141 20671 30175
rect 21373 30141 21407 30175
rect 22845 30141 22879 30175
rect 23489 30141 23523 30175
rect 23756 30141 23790 30175
rect 25697 30141 25731 30175
rect 25789 30141 25823 30175
rect 26065 30141 26099 30175
rect 26617 30141 26651 30175
rect 27805 30141 27839 30175
rect 29837 30277 29871 30311
rect 57069 30277 57103 30311
rect 30573 30209 30607 30243
rect 36553 30209 36587 30243
rect 57529 30209 57563 30243
rect 28549 30141 28583 30175
rect 29193 30141 29227 30175
rect 29837 30141 29871 30175
rect 30021 30141 30055 30175
rect 30481 30141 30515 30175
rect 30665 30141 30699 30175
rect 31125 30141 31159 30175
rect 31309 30141 31343 30175
rect 35449 30141 35483 30175
rect 35541 30141 35575 30175
rect 36185 30141 36219 30175
rect 36369 30141 36403 30175
rect 54769 30141 54803 30175
rect 57713 30141 57747 30175
rect 29285 30073 29319 30107
rect 35725 30073 35759 30107
rect 55321 30073 55355 30107
rect 55413 30073 55447 30107
rect 55965 30073 55999 30107
rect 56885 30073 56919 30107
rect 58173 30073 58207 30107
rect 9505 30005 9539 30039
rect 11069 30005 11103 30039
rect 13093 30005 13127 30039
rect 15209 30005 15243 30039
rect 15761 30005 15795 30039
rect 22937 30005 22971 30039
rect 27905 30005 27939 30039
rect 28457 30005 28491 30039
rect 28641 30005 28675 30039
rect 54585 30005 54619 30039
rect 16129 29801 16163 29835
rect 16681 29801 16715 29835
rect 54401 29801 54435 29835
rect 12357 29733 12391 29767
rect 14994 29733 15028 29767
rect 17969 29733 18003 29767
rect 20085 29733 20119 29767
rect 21158 29733 21192 29767
rect 30748 29733 30782 29767
rect 55229 29733 55263 29767
rect 55781 29733 55815 29767
rect 56885 29733 56919 29767
rect 57437 29733 57471 29767
rect 1869 29665 1903 29699
rect 6469 29665 6503 29699
rect 7113 29665 7147 29699
rect 7297 29665 7331 29699
rect 8125 29665 8159 29699
rect 9505 29665 9539 29699
rect 9689 29665 9723 29699
rect 10784 29665 10818 29699
rect 12504 29665 12538 29699
rect 13645 29665 13679 29699
rect 13829 29665 13863 29699
rect 16589 29665 16623 29699
rect 16773 29665 16807 29699
rect 17233 29665 17267 29699
rect 17693 29665 17727 29699
rect 18613 29665 18647 29699
rect 18705 29665 18739 29699
rect 18889 29665 18923 29699
rect 19993 29665 20027 29699
rect 22753 29665 22787 29699
rect 22845 29665 22879 29699
rect 23857 29665 23891 29699
rect 24041 29665 24075 29699
rect 25237 29665 25271 29699
rect 26341 29665 26375 29699
rect 26433 29665 26467 29699
rect 26617 29665 26651 29699
rect 26709 29665 26743 29699
rect 27353 29665 27387 29699
rect 27997 29665 28031 29699
rect 28181 29665 28215 29699
rect 28273 29665 28307 29699
rect 28549 29665 28583 29699
rect 29009 29665 29043 29699
rect 32321 29665 32355 29699
rect 53757 29665 53791 29699
rect 54585 29665 54619 29699
rect 57989 29665 58023 29699
rect 10517 29597 10551 29631
rect 12725 29597 12759 29631
rect 14749 29597 14783 29631
rect 20913 29597 20947 29631
rect 23029 29597 23063 29631
rect 24317 29597 24351 29631
rect 28457 29597 28491 29631
rect 30481 29597 30515 29631
rect 55137 29597 55171 29631
rect 56793 29597 56827 29631
rect 12633 29529 12667 29563
rect 18797 29529 18831 29563
rect 22293 29529 22327 29563
rect 29101 29529 29135 29563
rect 31861 29529 31895 29563
rect 58173 29529 58207 29563
rect 1961 29461 1995 29495
rect 6561 29461 6595 29495
rect 7113 29461 7147 29495
rect 8217 29461 8251 29495
rect 9505 29461 9539 29495
rect 11897 29461 11931 29495
rect 13001 29461 13035 29495
rect 13645 29461 13679 29495
rect 18429 29461 18463 29495
rect 22937 29461 22971 29495
rect 24225 29461 24259 29495
rect 25329 29461 25363 29495
rect 26157 29461 26191 29495
rect 27445 29461 27479 29495
rect 32413 29461 32447 29495
rect 8217 29257 8251 29291
rect 12173 29257 12207 29291
rect 13185 29257 13219 29291
rect 18889 29257 18923 29291
rect 20453 29257 20487 29291
rect 24409 29257 24443 29291
rect 25053 29257 25087 29291
rect 27813 29257 27847 29291
rect 30205 29257 30239 29291
rect 54861 29257 54895 29291
rect 56149 29257 56183 29291
rect 57989 29257 58023 29291
rect 10149 29189 10183 29223
rect 15117 29189 15151 29223
rect 19349 29189 19383 29223
rect 23007 29189 23041 29223
rect 24225 29189 24259 29223
rect 35725 29189 35759 29223
rect 55689 29189 55723 29223
rect 57069 29189 57103 29223
rect 8769 29121 8803 29155
rect 13553 29121 13587 29155
rect 16405 29121 16439 29155
rect 23121 29121 23155 29155
rect 23213 29121 23247 29155
rect 24317 29121 24351 29155
rect 26617 29121 26651 29155
rect 28273 29121 28307 29155
rect 32137 29121 32171 29155
rect 36645 29121 36679 29155
rect 54401 29121 54435 29155
rect 57529 29121 57563 29155
rect 1869 29053 1903 29087
rect 5733 29053 5767 29087
rect 5917 29053 5951 29087
rect 6837 29053 6871 29087
rect 7104 29053 7138 29087
rect 9036 29053 9070 29087
rect 10609 29053 10643 29087
rect 12081 29053 12115 29087
rect 13093 29053 13127 29087
rect 14289 29053 14323 29087
rect 15025 29053 15059 29087
rect 15669 29053 15703 29087
rect 16129 29053 16163 29087
rect 17325 29053 17359 29087
rect 17785 29053 17819 29087
rect 19073 29053 19107 29087
rect 19165 29053 19199 29087
rect 19441 29053 19475 29087
rect 20709 29053 20743 29087
rect 20818 29053 20852 29087
rect 20913 29053 20947 29087
rect 21097 29053 21131 29087
rect 23305 29053 23339 29087
rect 24133 29053 24167 29087
rect 24501 29053 24535 29087
rect 25053 29053 25087 29087
rect 25237 29053 25271 29087
rect 25881 29053 25915 29087
rect 26065 29053 26099 29087
rect 26157 29053 26191 29087
rect 26295 29053 26329 29087
rect 26433 29053 26467 29087
rect 27997 29053 28031 29087
rect 28089 29053 28123 29087
rect 28365 29053 28399 29087
rect 28825 29053 28859 29087
rect 30941 29053 30975 29087
rect 31585 29053 31619 29087
rect 31769 29053 31803 29087
rect 33287 29053 33321 29087
rect 33425 29053 33459 29087
rect 33517 29053 33551 29087
rect 33701 29053 33735 29087
rect 35449 29053 35483 29087
rect 35633 29053 35667 29087
rect 36277 29053 36311 29087
rect 36461 29053 36495 29087
rect 55045 29053 55079 29087
rect 55505 29053 55539 29087
rect 56333 29053 56367 29087
rect 57713 29053 57747 29087
rect 2053 28985 2087 29019
rect 14105 28985 14139 29019
rect 14473 28985 14507 29019
rect 18061 28985 18095 29019
rect 22937 28985 22971 29019
rect 29070 28985 29104 29019
rect 33057 28985 33091 29019
rect 56885 28985 56919 29019
rect 5825 28917 5859 28951
rect 10701 28917 10735 28951
rect 23857 28917 23891 28951
rect 31033 28917 31067 28951
rect 32045 28917 32079 28951
rect 6561 28713 6595 28747
rect 7665 28713 7699 28747
rect 21373 28713 21407 28747
rect 21833 28713 21867 28747
rect 22937 28713 22971 28747
rect 26157 28713 26191 28747
rect 28089 28713 28123 28747
rect 28549 28713 28583 28747
rect 32321 28713 32355 28747
rect 34437 28713 34471 28747
rect 5448 28645 5482 28679
rect 10885 28645 10919 28679
rect 13553 28645 13587 28679
rect 14994 28645 15028 28679
rect 20260 28645 20294 28679
rect 27353 28645 27387 28679
rect 27813 28645 27847 28679
rect 31217 28645 31251 28679
rect 33302 28645 33336 28679
rect 55229 28645 55263 28679
rect 55781 28645 55815 28679
rect 56885 28645 56919 28679
rect 58173 28645 58207 28679
rect 1501 28577 1535 28611
rect 2789 28577 2823 28611
rect 4537 28577 4571 28611
rect 4721 28577 4755 28611
rect 5181 28577 5215 28611
rect 7021 28577 7055 28611
rect 7205 28577 7239 28611
rect 7849 28577 7883 28611
rect 7941 28577 7975 28611
rect 8217 28577 8251 28611
rect 9689 28577 9723 28611
rect 9781 28577 9815 28611
rect 10057 28577 10091 28611
rect 11161 28577 11195 28611
rect 11529 28577 11563 28611
rect 12541 28577 12575 28611
rect 12725 28577 12759 28611
rect 13001 28577 13035 28611
rect 16589 28577 16623 28611
rect 16773 28577 16807 28611
rect 17233 28577 17267 28611
rect 17785 28577 17819 28611
rect 18705 28577 18739 28611
rect 18797 28577 18831 28611
rect 18889 28577 18923 28611
rect 19073 28577 19107 28611
rect 19993 28577 20027 28611
rect 22017 28577 22051 28611
rect 22109 28577 22143 28611
rect 22385 28577 22419 28611
rect 23121 28577 23155 28611
rect 23213 28577 23247 28611
rect 23489 28577 23523 28611
rect 23949 28577 23983 28611
rect 25513 28577 25547 28611
rect 26709 28577 26743 28611
rect 26893 28577 26927 28611
rect 1685 28509 1719 28543
rect 10701 28509 10735 28543
rect 11253 28509 11287 28543
rect 11437 28509 11471 28543
rect 12633 28509 12667 28543
rect 12817 28509 12851 28543
rect 14749 28509 14783 28543
rect 17877 28509 17911 28543
rect 22293 28509 22327 28543
rect 24041 28509 24075 28543
rect 25881 28509 25915 28543
rect 1869 28441 1903 28475
rect 4537 28441 4571 28475
rect 12357 28441 12391 28475
rect 25789 28441 25823 28475
rect 27445 28577 27479 28611
rect 27583 28577 27617 28611
rect 27721 28577 27755 28611
rect 27910 28577 27944 28611
rect 28779 28577 28813 28611
rect 28917 28577 28951 28611
rect 29009 28577 29043 28611
rect 29193 28577 29227 28611
rect 30941 28577 30975 28611
rect 31125 28577 31159 28611
rect 31666 28577 31700 28611
rect 31770 28577 31804 28611
rect 31953 28577 31987 28611
rect 32045 28577 32079 28611
rect 32183 28577 32217 28611
rect 35725 28577 35759 28611
rect 54401 28577 54435 28611
rect 57989 28577 58023 28611
rect 33057 28509 33091 28543
rect 55137 28509 55171 28543
rect 56793 28509 56827 28543
rect 57437 28509 57471 28543
rect 7021 28373 7055 28407
rect 8125 28373 8159 28407
rect 9505 28373 9539 28407
rect 9965 28373 9999 28407
rect 13645 28373 13679 28407
rect 16129 28373 16163 28407
rect 16681 28373 16715 28407
rect 18429 28373 18463 28407
rect 23397 28373 23431 28407
rect 25651 28373 25685 28407
rect 26709 28373 26743 28407
rect 27353 28373 27387 28407
rect 35909 28373 35943 28407
rect 2973 28169 3007 28203
rect 7113 28169 7147 28203
rect 19993 28169 20027 28203
rect 21281 28169 21315 28203
rect 23397 28169 23431 28203
rect 25973 28169 26007 28203
rect 28365 28169 28399 28203
rect 55321 28169 55355 28203
rect 56241 28169 56275 28203
rect 57253 28169 57287 28203
rect 11161 28101 11195 28135
rect 19349 28101 19383 28135
rect 23949 28101 23983 28135
rect 24777 28101 24811 28135
rect 2605 28033 2639 28067
rect 7573 28033 7607 28067
rect 13001 28033 13035 28067
rect 15761 28033 15795 28067
rect 17417 28033 17451 28067
rect 19901 28033 19935 28067
rect 20085 28033 20119 28067
rect 24501 28033 24535 28067
rect 31309 28033 31343 28067
rect 31401 28033 31435 28067
rect 33793 28033 33827 28067
rect 35725 28033 35759 28067
rect 2789 27965 2823 27999
rect 4445 27965 4479 27999
rect 4629 27965 4663 27999
rect 5089 27965 5123 27999
rect 5273 27965 5307 27999
rect 7297 27965 7331 27999
rect 7389 27965 7423 27999
rect 7665 27965 7699 27999
rect 8585 27965 8619 27999
rect 10977 27965 11011 27999
rect 12081 27965 12115 27999
rect 12725 27965 12759 27999
rect 13737 27965 13771 27999
rect 14473 27965 14507 27999
rect 15117 27965 15151 27999
rect 15301 27965 15335 27999
rect 15945 27965 15979 27999
rect 16313 27965 16347 27999
rect 17325 27965 17359 27999
rect 17969 27965 18003 27999
rect 18236 27965 18270 27999
rect 19809 27965 19843 27999
rect 20637 27965 20671 27999
rect 20730 27965 20764 27999
rect 21102 27965 21136 27999
rect 22845 27965 22879 27999
rect 23213 27965 23247 27999
rect 23857 27965 23891 27999
rect 24685 27965 24719 27999
rect 25053 27965 25087 27999
rect 26157 27965 26191 27999
rect 26249 27965 26283 27999
rect 26433 27965 26467 27999
rect 26525 27965 26559 27999
rect 27813 27965 27847 27999
rect 28089 27965 28123 27999
rect 28181 27965 28215 27999
rect 29101 27965 29135 27999
rect 31125 27965 31159 27999
rect 31217 27965 31251 27999
rect 31585 27965 31619 27999
rect 33057 27965 33091 27999
rect 33701 27965 33735 27999
rect 34345 27965 34379 27999
rect 34529 27965 34563 27999
rect 35449 27965 35483 27999
rect 35541 27965 35575 27999
rect 36277 27965 36311 27999
rect 36369 27965 36403 27999
rect 55505 27965 55539 27999
rect 56425 27965 56459 27999
rect 57437 27965 57471 27999
rect 1869 27897 1903 27931
rect 8830 27897 8864 27931
rect 13921 27897 13955 27931
rect 14565 27897 14599 27931
rect 20913 27897 20947 27931
rect 21005 27897 21039 27931
rect 23029 27897 23063 27931
rect 23121 27897 23155 27931
rect 24961 27897 24995 27931
rect 27997 27897 28031 27931
rect 29368 27897 29402 27931
rect 34437 27897 34471 27931
rect 36553 27897 36587 27931
rect 57989 27897 58023 27931
rect 58173 27897 58207 27931
rect 1961 27829 1995 27863
rect 4537 27829 4571 27863
rect 5181 27829 5215 27863
rect 9965 27829 9999 27863
rect 12173 27829 12207 27863
rect 15209 27829 15243 27863
rect 16221 27829 16255 27863
rect 30481 27829 30515 27863
rect 30941 27829 30975 27863
rect 33149 27829 33183 27863
rect 2513 27625 2547 27659
rect 3157 27625 3191 27659
rect 7205 27625 7239 27659
rect 16497 27625 16531 27659
rect 29101 27625 29135 27659
rect 58173 27625 58207 27659
rect 5457 27557 5491 27591
rect 20269 27557 20303 27591
rect 22477 27557 22511 27591
rect 23581 27557 23615 27591
rect 24225 27557 24259 27591
rect 26065 27557 26099 27591
rect 1869 27489 1903 27523
rect 2697 27489 2731 27523
rect 3341 27489 3375 27523
rect 4629 27489 4663 27523
rect 7389 27489 7423 27523
rect 7481 27489 7515 27523
rect 7757 27489 7791 27523
rect 8309 27489 8343 27523
rect 9689 27489 9723 27523
rect 9781 27489 9815 27523
rect 10057 27489 10091 27523
rect 11069 27489 11103 27523
rect 11325 27489 11359 27523
rect 13461 27489 13495 27523
rect 15393 27489 15427 27523
rect 15577 27489 15611 27523
rect 15853 27489 15887 27523
rect 16313 27489 16347 27523
rect 16589 27489 16623 27523
rect 17233 27489 17267 27523
rect 17371 27489 17405 27523
rect 17601 27489 17635 27523
rect 18245 27489 18279 27523
rect 18429 27489 18463 27523
rect 19993 27489 20027 27523
rect 20086 27489 20120 27523
rect 20361 27489 20395 27523
rect 20458 27489 20492 27523
rect 21189 27489 21223 27523
rect 21373 27489 21407 27523
rect 21833 27489 21867 27523
rect 22661 27489 22695 27523
rect 22753 27489 22787 27523
rect 23029 27489 23063 27523
rect 23489 27489 23523 27523
rect 24133 27489 24167 27523
rect 25697 27489 25731 27523
rect 25881 27489 25915 27523
rect 26525 27489 26559 27523
rect 26617 27489 26651 27523
rect 27436 27489 27470 27523
rect 29009 27489 29043 27523
rect 30849 27489 30883 27523
rect 31585 27489 31619 27523
rect 32597 27489 32631 27523
rect 33681 27489 33715 27523
rect 35725 27489 35759 27523
rect 55597 27489 55631 27523
rect 56885 27489 56919 27523
rect 5365 27421 5399 27455
rect 6377 27421 6411 27455
rect 7665 27421 7699 27455
rect 9965 27421 9999 27455
rect 13737 27421 13771 27455
rect 15209 27421 15243 27455
rect 15669 27421 15703 27455
rect 18337 27421 18371 27455
rect 18521 27421 18555 27455
rect 21281 27421 21315 27455
rect 21925 27421 21959 27455
rect 22937 27421 22971 27455
rect 27169 27421 27203 27455
rect 31125 27421 31159 27455
rect 33425 27421 33459 27455
rect 57529 27421 57563 27455
rect 57713 27421 57747 27455
rect 13645 27353 13679 27387
rect 15485 27353 15519 27387
rect 16313 27353 16347 27387
rect 17509 27353 17543 27387
rect 25697 27353 25731 27387
rect 31033 27353 31067 27387
rect 1961 27285 1995 27319
rect 4813 27285 4847 27319
rect 8401 27285 8435 27319
rect 9505 27285 9539 27319
rect 12449 27285 12483 27319
rect 13553 27285 13587 27319
rect 17049 27285 17083 27319
rect 18061 27285 18095 27319
rect 20637 27285 20671 27319
rect 28549 27285 28583 27319
rect 30941 27285 30975 27319
rect 31677 27285 31711 27319
rect 32689 27285 32723 27319
rect 34805 27285 34839 27319
rect 35909 27285 35943 27319
rect 56977 27285 57011 27319
rect 1869 27081 1903 27115
rect 5457 27081 5491 27115
rect 11161 27081 11195 27115
rect 21097 27081 21131 27115
rect 24041 27081 24075 27115
rect 24685 27081 24719 27115
rect 26065 27081 26099 27115
rect 27813 27081 27847 27115
rect 33057 27081 33091 27115
rect 56793 27081 56827 27115
rect 57253 27081 57287 27115
rect 2605 27013 2639 27047
rect 8953 27013 8987 27047
rect 12909 27013 12943 27047
rect 14289 27013 14323 27047
rect 15117 27013 15151 27047
rect 16313 27013 16347 27047
rect 17785 27013 17819 27047
rect 28181 27013 28215 27047
rect 29193 27013 29227 27047
rect 1685 26945 1719 26979
rect 6837 26945 6871 26979
rect 10701 26945 10735 26979
rect 13001 26945 13035 26979
rect 13740 26945 13774 26979
rect 14473 26945 14507 26979
rect 17325 26945 17359 26979
rect 21281 26945 21315 26979
rect 26525 26945 26559 26979
rect 28273 26945 28307 26979
rect 29285 26945 29319 26979
rect 34805 26945 34839 26979
rect 56057 26945 56091 26979
rect 1501 26877 1535 26911
rect 2789 26877 2823 26911
rect 3433 26877 3467 26911
rect 4077 26877 4111 26911
rect 4537 26877 4571 26911
rect 4721 26877 4755 26911
rect 5273 26877 5307 26911
rect 7104 26877 7138 26911
rect 10425 26877 10459 26911
rect 10609 26877 10643 26911
rect 10793 26877 10827 26911
rect 10977 26877 11011 26911
rect 12081 26877 12115 26911
rect 12725 26877 12759 26911
rect 12817 26877 12851 26911
rect 13461 26877 13495 26911
rect 13553 26877 13587 26911
rect 14197 26877 14231 26911
rect 14933 26877 14967 26911
rect 15577 26877 15611 26911
rect 15669 26877 15703 26911
rect 16221 26877 16255 26911
rect 17509 26877 17543 26911
rect 17601 26877 17635 26911
rect 17877 26877 17911 26911
rect 18337 26877 18371 26911
rect 18981 26877 19015 26911
rect 21005 26877 21039 26911
rect 22661 26877 22695 26911
rect 25421 26877 25455 26911
rect 26249 26877 26283 26911
rect 26341 26877 26375 26911
rect 26617 26877 26651 26911
rect 27997 26877 28031 26911
rect 29101 26877 29135 26911
rect 29377 26877 29411 26911
rect 29561 26877 29595 26911
rect 30021 26877 30055 26911
rect 30205 26877 30239 26911
rect 30389 26877 30423 26911
rect 31677 26877 31711 26911
rect 33333 26877 33367 26911
rect 33425 26877 33459 26911
rect 33517 26877 33551 26911
rect 33701 26877 33735 26911
rect 34161 26877 34195 26911
rect 57437 26877 57471 26911
rect 8769 26809 8803 26843
rect 9781 26809 9815 26843
rect 9965 26809 9999 26843
rect 13737 26809 13771 26843
rect 14473 26809 14507 26843
rect 18429 26809 18463 26843
rect 19248 26809 19282 26843
rect 22928 26809 22962 26843
rect 24593 26809 24627 26843
rect 25237 26809 25271 26843
rect 25605 26809 25639 26843
rect 30297 26809 30331 26843
rect 31493 26809 31527 26843
rect 35072 26809 35106 26843
rect 55413 26809 55447 26843
rect 55505 26809 55539 26843
rect 57989 26809 58023 26843
rect 3249 26741 3283 26775
rect 3893 26741 3927 26775
rect 4629 26741 4663 26775
rect 8217 26741 8251 26775
rect 12265 26741 12299 26775
rect 20361 26741 20395 26775
rect 21281 26741 21315 26775
rect 28917 26741 28951 26775
rect 30573 26741 30607 26775
rect 31861 26741 31895 26775
rect 34253 26741 34287 26775
rect 36185 26741 36219 26775
rect 58081 26741 58115 26775
rect 2513 26537 2547 26571
rect 7573 26537 7607 26571
rect 8493 26537 8527 26571
rect 16129 26537 16163 26571
rect 25697 26537 25731 26571
rect 27169 26537 27203 26571
rect 29561 26537 29595 26571
rect 31309 26537 31343 26571
rect 32137 26537 32171 26571
rect 33241 26537 33275 26571
rect 37197 26537 37231 26571
rect 55781 26537 55815 26571
rect 58173 26537 58207 26571
rect 4629 26469 4663 26503
rect 13829 26469 13863 26503
rect 15016 26469 15050 26503
rect 23489 26469 23523 26503
rect 31125 26469 31159 26503
rect 32965 26469 32999 26503
rect 1869 26401 1903 26435
rect 2053 26401 2087 26435
rect 3065 26401 3099 26435
rect 4537 26401 4571 26435
rect 4721 26401 4755 26435
rect 5365 26401 5399 26435
rect 6193 26401 6227 26435
rect 6837 26401 6871 26435
rect 7021 26401 7055 26435
rect 7481 26401 7515 26435
rect 8401 26401 8435 26435
rect 8585 26401 8619 26435
rect 9781 26401 9815 26435
rect 9965 26401 9999 26435
rect 10057 26401 10091 26435
rect 10333 26401 10367 26435
rect 10977 26401 11011 26435
rect 11161 26401 11195 26435
rect 11262 26401 11296 26435
rect 11529 26401 11563 26435
rect 12173 26401 12207 26435
rect 12357 26401 12391 26435
rect 12449 26401 12483 26435
rect 12725 26401 12759 26435
rect 13553 26401 13587 26435
rect 16773 26401 16807 26435
rect 16865 26401 16899 26435
rect 17141 26401 17175 26435
rect 17693 26401 17727 26435
rect 20821 26401 20855 26435
rect 21465 26401 21499 26435
rect 21658 26401 21692 26435
rect 21925 26401 21959 26435
rect 22477 26401 22511 26435
rect 23305 26401 23339 26435
rect 23949 26401 23983 26435
rect 25421 26401 25455 26435
rect 26617 26401 26651 26435
rect 26801 26401 26835 26435
rect 26893 26401 26927 26435
rect 27031 26401 27065 26435
rect 28448 26401 28482 26435
rect 30941 26401 30975 26435
rect 31769 26401 31803 26435
rect 31953 26401 31987 26435
rect 32597 26401 32631 26435
rect 32745 26401 32779 26435
rect 32873 26401 32907 26435
rect 33062 26401 33096 26435
rect 33701 26401 33735 26435
rect 33886 26401 33920 26435
rect 33977 26401 34011 26435
rect 34253 26401 34287 26435
rect 36369 26401 36403 26435
rect 36461 26401 36495 26435
rect 37105 26401 37139 26435
rect 37289 26401 37323 26435
rect 55137 26401 55171 26435
rect 10149 26333 10183 26367
rect 11345 26333 11379 26367
rect 12541 26333 12575 26367
rect 13829 26333 13863 26367
rect 14749 26333 14783 26367
rect 17877 26333 17911 26367
rect 18337 26333 18371 26367
rect 20177 26333 20211 26367
rect 21557 26333 21591 26367
rect 21741 26333 21775 26367
rect 25237 26333 25271 26367
rect 25789 26333 25823 26367
rect 28181 26333 28215 26367
rect 55321 26333 55355 26367
rect 57069 26333 57103 26367
rect 57529 26333 57563 26367
rect 57713 26333 57747 26367
rect 6837 26265 6871 26299
rect 13645 26265 13679 26299
rect 16589 26265 16623 26299
rect 18981 26265 19015 26299
rect 22661 26265 22695 26299
rect 34161 26265 34195 26299
rect 36553 26265 36587 26299
rect 3157 26197 3191 26231
rect 6285 26197 6319 26231
rect 10517 26197 10551 26231
rect 11713 26197 11747 26231
rect 12909 26197 12943 26231
rect 17049 26197 17083 26231
rect 21281 26197 21315 26231
rect 24133 26197 24167 26231
rect 25513 26197 25547 26231
rect 2605 25993 2639 26027
rect 5917 25993 5951 26027
rect 29377 25993 29411 26027
rect 30113 25993 30147 26027
rect 31953 25993 31987 26027
rect 33057 25993 33091 26027
rect 34897 25993 34931 26027
rect 55321 25993 55355 26027
rect 55965 25993 55999 26027
rect 8309 25925 8343 25959
rect 10701 25925 10735 25959
rect 15669 25925 15703 25959
rect 19625 25925 19659 25959
rect 23213 25925 23247 25959
rect 25513 25925 25547 25959
rect 30757 25925 30791 25959
rect 31125 25925 31159 25959
rect 33517 25925 33551 25959
rect 34161 25925 34195 25959
rect 1961 25857 1995 25891
rect 2145 25857 2179 25891
rect 6929 25857 6963 25891
rect 15025 25857 15059 25891
rect 19257 25857 19291 25891
rect 20545 25857 20579 25891
rect 22569 25857 22603 25891
rect 26341 25857 26375 25891
rect 34345 25857 34379 25891
rect 36645 25857 36679 25891
rect 3617 25789 3651 25823
rect 3709 25789 3743 25823
rect 4537 25789 4571 25823
rect 8769 25789 8803 25823
rect 9036 25789 9070 25823
rect 10609 25789 10643 25823
rect 12081 25789 12115 25823
rect 12348 25789 12382 25823
rect 14933 25789 14967 25823
rect 15117 25789 15151 25823
rect 15577 25789 15611 25823
rect 16221 25789 16255 25823
rect 17877 25789 17911 25823
rect 18877 25789 18911 25823
rect 19077 25789 19111 25823
rect 19165 25789 19199 25823
rect 19441 25789 19475 25823
rect 20361 25789 20395 25823
rect 21097 25789 21131 25823
rect 24133 25789 24167 25823
rect 25973 25789 26007 25823
rect 26157 25789 26191 25823
rect 26249 25789 26283 25823
rect 26525 25789 26559 25823
rect 29285 25789 29319 25823
rect 30021 25789 30055 25823
rect 30941 25789 30975 25823
rect 31033 25789 31067 25823
rect 31217 25789 31251 25823
rect 31769 25789 31803 25823
rect 31953 25789 31987 25823
rect 33241 25789 33275 25823
rect 33333 25789 33367 25823
rect 33609 25789 33643 25823
rect 34069 25789 34103 25823
rect 34805 25789 34839 25823
rect 35633 25789 35667 25823
rect 36369 25789 36403 25823
rect 36461 25789 36495 25823
rect 55505 25789 55539 25823
rect 56149 25789 56183 25823
rect 56609 25789 56643 25823
rect 57253 25789 57287 25823
rect 57989 25789 58023 25823
rect 4804 25721 4838 25755
rect 7196 25721 7230 25755
rect 14013 25721 14047 25755
rect 14197 25721 14231 25755
rect 24400 25721 24434 25755
rect 26709 25721 26743 25755
rect 27905 25721 27939 25755
rect 28641 25721 28675 25755
rect 28825 25721 28859 25755
rect 58173 25721 58207 25755
rect 3893 25653 3927 25687
rect 10149 25653 10183 25687
rect 13461 25653 13495 25687
rect 16313 25653 16347 25687
rect 18429 25653 18463 25687
rect 21649 25653 21683 25687
rect 27997 25653 28031 25687
rect 32137 25653 32171 25687
rect 34345 25653 34379 25687
rect 35725 25653 35759 25687
rect 57437 25653 57471 25687
rect 5181 25449 5215 25483
rect 7481 25449 7515 25483
rect 17969 25449 18003 25483
rect 21373 25449 21407 25483
rect 23213 25449 23247 25483
rect 28273 25449 28307 25483
rect 31861 25449 31895 25483
rect 32321 25449 32355 25483
rect 34345 25449 34379 25483
rect 57989 25449 58023 25483
rect 9781 25381 9815 25415
rect 11060 25381 11094 25415
rect 13645 25381 13679 25415
rect 16497 25381 16531 25415
rect 20260 25381 20294 25415
rect 22078 25381 22112 25415
rect 24133 25381 24167 25415
rect 27160 25381 27194 25415
rect 57161 25381 57195 25415
rect 1869 25313 1903 25347
rect 3157 25313 3191 25347
rect 4261 25313 4295 25347
rect 4445 25313 4479 25347
rect 5089 25313 5123 25347
rect 5273 25313 5307 25347
rect 5917 25313 5951 25347
rect 6009 25313 6043 25347
rect 6285 25313 6319 25347
rect 6837 25313 6871 25347
rect 7665 25313 7699 25347
rect 7757 25313 7791 25347
rect 8033 25313 8067 25347
rect 9597 25313 9631 25347
rect 12909 25313 12943 25347
rect 14933 25313 14967 25347
rect 15853 25313 15887 25347
rect 16681 25313 16715 25347
rect 16773 25313 16807 25347
rect 17325 25313 17359 25347
rect 18245 25313 18279 25347
rect 18337 25313 18371 25347
rect 18434 25313 18468 25347
rect 18613 25313 18647 25347
rect 23949 25313 23983 25347
rect 25237 25313 25271 25347
rect 25421 25313 25455 25347
rect 25513 25313 25547 25347
rect 25789 25313 25823 25347
rect 28825 25313 28859 25347
rect 29009 25313 29043 25347
rect 29377 25313 29411 25347
rect 30481 25313 30515 25347
rect 31125 25313 31159 25347
rect 31309 25313 31343 25347
rect 31677 25313 31711 25347
rect 32505 25313 32539 25347
rect 32781 25313 32815 25347
rect 33793 25313 33827 25347
rect 33977 25313 34011 25347
rect 34069 25313 34103 25347
rect 34207 25313 34241 25347
rect 35725 25313 35759 25347
rect 36461 25313 36495 25347
rect 36553 25313 36587 25347
rect 37197 25313 37231 25347
rect 37381 25313 37415 25347
rect 55597 25313 55631 25347
rect 58173 25313 58207 25347
rect 2973 25245 3007 25279
rect 5733 25245 5767 25279
rect 7021 25245 7055 25279
rect 10793 25245 10827 25279
rect 13001 25245 13035 25279
rect 19993 25245 20027 25279
rect 21833 25245 21867 25279
rect 25605 25245 25639 25279
rect 26893 25245 26927 25279
rect 29101 25245 29135 25279
rect 29193 25245 29227 25279
rect 31401 25245 31435 25279
rect 31493 25245 31527 25279
rect 32597 25245 32631 25279
rect 32689 25245 32723 25279
rect 36737 25245 36771 25279
rect 15945 25177 15979 25211
rect 1961 25109 1995 25143
rect 3341 25109 3375 25143
rect 4629 25109 4663 25143
rect 6193 25109 6227 25143
rect 7941 25109 7975 25143
rect 12173 25109 12207 25143
rect 13737 25109 13771 25143
rect 15209 25109 15243 25143
rect 16497 25109 16531 25143
rect 17417 25109 17451 25143
rect 25973 25109 26007 25143
rect 29561 25109 29595 25143
rect 30573 25109 30607 25143
rect 35817 25109 35851 25143
rect 37197 25109 37231 25143
rect 55413 25109 55447 25143
rect 57253 25109 57287 25143
rect 2329 24905 2363 24939
rect 13645 24905 13679 24939
rect 26893 24905 26927 24939
rect 30481 24905 30515 24939
rect 32045 24905 32079 24939
rect 17693 24837 17727 24871
rect 24133 24837 24167 24871
rect 33701 24837 33735 24871
rect 1961 24769 1995 24803
rect 3525 24769 3559 24803
rect 10517 24769 10551 24803
rect 20545 24769 20579 24803
rect 21097 24769 21131 24803
rect 24869 24769 24903 24803
rect 31585 24769 31619 24803
rect 54677 24769 54711 24803
rect 56241 24769 56275 24803
rect 2145 24701 2179 24735
rect 3709 24701 3743 24735
rect 4721 24701 4755 24735
rect 4905 24701 4939 24735
rect 5365 24701 5399 24735
rect 7389 24701 7423 24735
rect 8033 24701 8067 24735
rect 8309 24701 8343 24735
rect 9321 24701 9355 24735
rect 10149 24701 10183 24735
rect 10333 24701 10367 24735
rect 10425 24701 10459 24735
rect 10701 24701 10735 24735
rect 12633 24701 12667 24735
rect 13461 24701 13495 24735
rect 14565 24701 14599 24735
rect 17325 24701 17359 24735
rect 17509 24701 17543 24735
rect 18344 24701 18378 24735
rect 18604 24701 18638 24735
rect 20361 24701 20395 24735
rect 21649 24701 21683 24735
rect 22753 24701 22787 24735
rect 25513 24701 25547 24735
rect 25780 24701 25814 24735
rect 29009 24701 29043 24735
rect 29101 24701 29135 24735
rect 29368 24701 29402 24735
rect 30941 24701 30975 24735
rect 31769 24701 31803 24735
rect 31861 24701 31895 24735
rect 32137 24701 32171 24735
rect 33425 24701 33459 24735
rect 33563 24701 33597 24735
rect 33793 24701 33827 24735
rect 34621 24701 34655 24735
rect 34888 24701 34922 24735
rect 36461 24701 36495 24735
rect 36645 24701 36679 24735
rect 54493 24701 54527 24735
rect 55137 24701 55171 24735
rect 55597 24701 55631 24735
rect 55781 24701 55815 24735
rect 57069 24701 57103 24735
rect 57529 24701 57563 24735
rect 57713 24701 57747 24735
rect 13277 24633 13311 24667
rect 14810 24633 14844 24667
rect 23397 24633 23431 24667
rect 23949 24633 23983 24667
rect 24685 24633 24719 24667
rect 27905 24633 27939 24667
rect 3893 24565 3927 24599
rect 4813 24565 4847 24599
rect 5457 24565 5491 24599
rect 7481 24565 7515 24599
rect 9505 24565 9539 24599
rect 10885 24565 10919 24599
rect 12817 24565 12851 24599
rect 15945 24565 15979 24599
rect 19717 24565 19751 24599
rect 27997 24565 28031 24599
rect 29009 24565 29043 24599
rect 31033 24565 31067 24599
rect 33241 24565 33275 24599
rect 36001 24565 36035 24599
rect 36737 24565 36771 24599
rect 56885 24565 56919 24599
rect 58173 24565 58207 24599
rect 5641 24361 5675 24395
rect 6101 24361 6135 24395
rect 8493 24361 8527 24395
rect 13645 24361 13679 24395
rect 17233 24361 17267 24395
rect 21741 24361 21775 24395
rect 22845 24361 22879 24395
rect 29561 24361 29595 24395
rect 31585 24361 31619 24395
rect 32505 24361 32539 24395
rect 35909 24361 35943 24395
rect 55505 24361 55539 24395
rect 4528 24293 4562 24327
rect 9772 24293 9806 24327
rect 16120 24293 16154 24327
rect 19073 24293 19107 24327
rect 20913 24293 20947 24327
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 6285 24225 6319 24259
rect 6377 24225 6411 24259
rect 6653 24225 6687 24259
rect 7481 24225 7515 24259
rect 7573 24225 7607 24259
rect 7849 24225 7883 24259
rect 8401 24225 8435 24259
rect 11345 24225 11379 24259
rect 11529 24225 11563 24259
rect 11713 24225 11747 24259
rect 11897 24225 11931 24259
rect 12725 24225 12759 24259
rect 13369 24225 13403 24259
rect 14841 24225 14875 24259
rect 17877 24225 17911 24259
rect 17969 24225 18003 24259
rect 18337 24225 18371 24259
rect 18889 24225 18923 24259
rect 22017 24293 22051 24327
rect 23489 24293 23523 24327
rect 26617 24293 26651 24327
rect 26801 24293 26835 24327
rect 57989 24293 58023 24327
rect 58173 24293 58207 24327
rect 22753 24225 22787 24259
rect 24133 24225 24167 24259
rect 25513 24225 25547 24259
rect 25697 24225 25731 24259
rect 25789 24225 25823 24259
rect 25881 24225 25915 24259
rect 30665 24225 30699 24259
rect 31309 24225 31343 24259
rect 31401 24225 31435 24259
rect 32413 24225 32447 24259
rect 33313 24225 33347 24259
rect 35817 24225 35851 24259
rect 55689 24225 55723 24259
rect 57437 24225 57471 24259
rect 1593 24157 1627 24191
rect 2697 24157 2731 24191
rect 4261 24157 4295 24191
rect 9505 24157 9539 24191
rect 11621 24157 11655 24191
rect 12081 24157 12115 24191
rect 13645 24157 13679 24191
rect 15853 24157 15887 24191
rect 18061 24157 18095 24191
rect 18153 24157 18187 24191
rect 20361 24157 20395 24191
rect 21741 24157 21775 24191
rect 27905 24157 27939 24191
rect 28917 24157 28951 24191
rect 30481 24157 30515 24191
rect 31585 24157 31619 24191
rect 33057 24157 33091 24191
rect 7757 24089 7791 24123
rect 12909 24089 12943 24123
rect 24317 24089 24351 24123
rect 1869 24021 1903 24055
rect 2881 24021 2915 24055
rect 6561 24021 6595 24055
rect 7297 24021 7331 24055
rect 10885 24021 10919 24055
rect 13461 24021 13495 24055
rect 15025 24021 15059 24055
rect 17693 24021 17727 24055
rect 22109 24021 22143 24055
rect 23581 24021 23615 24055
rect 26065 24021 26099 24055
rect 28457 24021 28491 24055
rect 30849 24021 30883 24055
rect 34437 24021 34471 24055
rect 5825 23817 5859 23851
rect 8861 23817 8895 23851
rect 9781 23817 9815 23851
rect 13461 23817 13495 23851
rect 14013 23817 14047 23851
rect 20361 23817 20395 23851
rect 29193 23817 29227 23851
rect 30481 23817 30515 23851
rect 32045 23817 32079 23851
rect 33057 23817 33091 23851
rect 56057 23817 56091 23851
rect 3617 23749 3651 23783
rect 10885 23749 10919 23783
rect 25053 23749 25087 23783
rect 34253 23749 34287 23783
rect 58173 23749 58207 23783
rect 2145 23681 2179 23715
rect 3249 23681 3283 23715
rect 5365 23681 5399 23715
rect 14197 23681 14231 23715
rect 15209 23681 15243 23715
rect 16313 23681 16347 23715
rect 18981 23681 19015 23715
rect 19625 23681 19659 23715
rect 27813 23681 27847 23715
rect 34805 23681 34839 23715
rect 1501 23613 1535 23647
rect 2329 23613 2363 23647
rect 3433 23613 3467 23647
rect 4721 23613 4755 23647
rect 4905 23613 4939 23647
rect 5549 23613 5583 23647
rect 5641 23613 5675 23647
rect 5917 23613 5951 23647
rect 6837 23613 6871 23647
rect 8769 23613 8803 23647
rect 9597 23613 9631 23647
rect 10609 23613 10643 23647
rect 12081 23613 12115 23647
rect 12348 23613 12382 23647
rect 13922 23613 13956 23647
rect 14933 23613 14967 23647
rect 15025 23613 15059 23647
rect 15301 23613 15335 23647
rect 16221 23613 16255 23647
rect 16405 23613 16439 23647
rect 17877 23613 17911 23647
rect 20085 23613 20119 23647
rect 22845 23613 22879 23647
rect 23673 23613 23707 23647
rect 23929 23613 23963 23647
rect 25513 23613 25547 23647
rect 26709 23613 26743 23647
rect 28080 23613 28114 23647
rect 30113 23613 30147 23647
rect 31125 23613 31159 23647
rect 31217 23613 31251 23647
rect 31401 23613 31435 23647
rect 31493 23613 31527 23647
rect 31953 23613 31987 23647
rect 33333 23613 33367 23647
rect 33425 23613 33459 23647
rect 33517 23613 33551 23647
rect 33701 23613 33735 23647
rect 34161 23613 34195 23647
rect 36645 23613 36679 23647
rect 55413 23613 55447 23647
rect 55597 23613 55631 23647
rect 56609 23613 56643 23647
rect 57253 23613 57287 23647
rect 7082 23545 7116 23579
rect 20269 23545 20303 23579
rect 21281 23545 21315 23579
rect 21465 23545 21499 23579
rect 22661 23545 22695 23579
rect 30297 23545 30331 23579
rect 35072 23545 35106 23579
rect 57989 23545 58023 23579
rect 1593 23477 1627 23511
rect 2789 23477 2823 23511
rect 4813 23477 4847 23511
rect 8217 23477 8251 23511
rect 14197 23477 14231 23511
rect 14749 23477 14783 23511
rect 18521 23477 18555 23511
rect 21649 23477 21683 23511
rect 26157 23477 26191 23511
rect 26801 23477 26835 23511
rect 30941 23477 30975 23511
rect 36185 23477 36219 23511
rect 36737 23477 36771 23511
rect 55229 23477 55263 23511
rect 3157 23273 3191 23307
rect 7021 23273 7055 23307
rect 10333 23273 10367 23307
rect 12357 23273 12391 23307
rect 13185 23273 13219 23307
rect 54677 23273 54711 23307
rect 1869 23205 1903 23239
rect 4874 23205 4908 23239
rect 2513 23137 2547 23171
rect 3341 23137 3375 23171
rect 4629 23137 4663 23171
rect 6929 23137 6963 23171
rect 7113 23137 7147 23171
rect 7849 23137 7883 23171
rect 9505 23137 9539 23171
rect 10149 23137 10183 23171
rect 10977 23137 11011 23171
rect 11161 23137 11195 23171
rect 11345 23137 11379 23171
rect 11529 23137 11563 23171
rect 12173 23137 12207 23171
rect 17960 23205 17994 23239
rect 25329 23205 25363 23239
rect 25513 23205 25547 23239
rect 26240 23205 26274 23239
rect 31769 23205 31803 23239
rect 32597 23205 32631 23239
rect 13277 23137 13311 23171
rect 14749 23137 14783 23171
rect 15016 23137 15050 23171
rect 17049 23137 17083 23171
rect 17693 23137 17727 23171
rect 20177 23137 20211 23171
rect 20637 23137 20671 23171
rect 21905 23137 21939 23171
rect 23857 23137 23891 23171
rect 24133 23137 24167 23171
rect 24317 23137 24351 23171
rect 27813 23137 27847 23171
rect 28917 23137 28951 23171
rect 29101 23137 29135 23171
rect 29377 23137 29411 23171
rect 31033 23137 31067 23171
rect 31217 23137 31251 23171
rect 31585 23137 31619 23171
rect 32229 23137 32263 23171
rect 32377 23137 32411 23171
rect 32505 23137 32539 23171
rect 32735 23137 32769 23171
rect 33333 23137 33367 23171
rect 33977 23137 34011 23171
rect 34161 23137 34195 23171
rect 34253 23137 34287 23171
rect 34529 23137 34563 23171
rect 36001 23137 36035 23171
rect 36093 23137 36127 23171
rect 54861 23137 54895 23171
rect 55321 23137 55355 23171
rect 57989 23137 58023 23171
rect 11253 23069 11287 23103
rect 13185 23069 13219 23103
rect 13553 23069 13587 23103
rect 20361 23069 20395 23103
rect 20470 23069 20504 23103
rect 21649 23069 21683 23103
rect 23673 23069 23707 23103
rect 24041 23069 24075 23103
rect 25973 23069 26007 23103
rect 29193 23069 29227 23103
rect 31309 23069 31343 23103
rect 31401 23069 31435 23103
rect 2697 23001 2731 23035
rect 9689 23001 9723 23035
rect 13461 23001 13495 23035
rect 20269 23001 20303 23035
rect 23949 23001 23983 23035
rect 27353 23001 27387 23035
rect 29009 23001 29043 23035
rect 32873 23001 32907 23035
rect 34437 23001 34471 23035
rect 55505 23001 55539 23035
rect 58173 23001 58207 23035
rect 1961 22933 1995 22967
rect 6009 22933 6043 22967
rect 7941 22933 7975 22967
rect 11713 22933 11747 22967
rect 13369 22933 13403 22967
rect 16129 22933 16163 22967
rect 17141 22933 17175 22967
rect 19073 22933 19107 22967
rect 19993 22933 20027 22967
rect 23029 22933 23063 22967
rect 27905 22933 27939 22967
rect 28733 22933 28767 22967
rect 33425 22933 33459 22967
rect 57437 22933 57471 22967
rect 14749 22729 14783 22763
rect 15669 22729 15703 22763
rect 19993 22729 20027 22763
rect 20361 22729 20395 22763
rect 21649 22729 21683 22763
rect 24133 22729 24167 22763
rect 28457 22729 28491 22763
rect 31217 22729 31251 22763
rect 31677 22729 31711 22763
rect 36001 22729 36035 22763
rect 57989 22729 58023 22763
rect 2145 22661 2179 22695
rect 3709 22661 3743 22695
rect 9873 22661 9907 22695
rect 14013 22661 14047 22695
rect 16313 22661 16347 22695
rect 19533 22661 19567 22695
rect 25237 22661 25271 22695
rect 29653 22661 29687 22695
rect 30205 22661 30239 22695
rect 30297 22661 30331 22695
rect 34253 22661 34287 22695
rect 54861 22661 54895 22695
rect 1777 22593 1811 22627
rect 3341 22593 3375 22627
rect 8493 22593 8527 22627
rect 10609 22593 10643 22627
rect 10701 22593 10735 22627
rect 12081 22593 12115 22627
rect 14197 22593 14231 22627
rect 14933 22593 14967 22627
rect 30389 22593 30423 22627
rect 55689 22593 55723 22627
rect 57529 22593 57563 22627
rect 1961 22525 1995 22559
rect 3525 22525 3559 22559
rect 5733 22525 5767 22559
rect 7481 22525 7515 22559
rect 7573 22525 7607 22559
rect 10333 22525 10367 22559
rect 10517 22525 10551 22559
rect 10885 22525 10919 22559
rect 12337 22525 12371 22559
rect 13921 22525 13955 22559
rect 14657 22525 14691 22559
rect 15577 22525 15611 22559
rect 16221 22525 16255 22559
rect 17601 22525 17635 22559
rect 18981 22525 19015 22559
rect 19257 22525 19291 22559
rect 19349 22525 19383 22559
rect 20177 22525 20211 22559
rect 20453 22525 20487 22559
rect 21005 22525 21039 22559
rect 21098 22525 21132 22559
rect 21511 22525 21545 22559
rect 22661 22525 22695 22559
rect 23765 22525 23799 22559
rect 23949 22525 23983 22559
rect 24593 22525 24627 22559
rect 24686 22525 24720 22559
rect 25099 22525 25133 22559
rect 25973 22525 26007 22559
rect 26062 22525 26096 22559
rect 26157 22525 26191 22559
rect 26341 22525 26375 22559
rect 27813 22525 27847 22559
rect 28457 22525 28491 22559
rect 28641 22525 28675 22559
rect 29101 22525 29135 22559
rect 29285 22525 29319 22559
rect 29469 22525 29503 22559
rect 30113 22525 30147 22559
rect 30849 22525 30883 22559
rect 31677 22525 31711 22559
rect 31861 22525 31895 22559
rect 33057 22525 33091 22559
rect 34161 22525 34195 22559
rect 35357 22525 35391 22559
rect 36001 22525 36035 22559
rect 36185 22525 36219 22559
rect 55045 22525 55079 22559
rect 55505 22525 55539 22559
rect 57713 22525 57747 22559
rect 4629 22457 4663 22491
rect 4997 22457 5031 22491
rect 8760 22457 8794 22491
rect 11069 22457 11103 22491
rect 18337 22457 18371 22491
rect 19165 22457 19199 22491
rect 21281 22457 21315 22491
rect 21373 22457 21407 22491
rect 24869 22457 24903 22491
rect 24961 22457 24995 22491
rect 29377 22457 29411 22491
rect 31033 22457 31067 22491
rect 56149 22457 56183 22491
rect 56885 22457 56919 22491
rect 57069 22457 57103 22491
rect 5825 22389 5859 22423
rect 7757 22389 7791 22423
rect 13461 22389 13495 22423
rect 14197 22389 14231 22423
rect 14933 22389 14967 22423
rect 17693 22389 17727 22423
rect 18429 22389 18463 22423
rect 22753 22389 22787 22423
rect 25697 22389 25731 22423
rect 27905 22389 27939 22423
rect 32045 22389 32079 22423
rect 33149 22389 33183 22423
rect 35449 22389 35483 22423
rect 7849 22185 7883 22219
rect 36369 22185 36403 22219
rect 4353 22117 4387 22151
rect 4445 22117 4479 22151
rect 11437 22117 11471 22151
rect 11989 22117 12023 22151
rect 12725 22117 12759 22151
rect 13369 22117 13403 22151
rect 14841 22117 14875 22151
rect 21005 22117 21039 22151
rect 23949 22117 23983 22151
rect 24133 22117 24167 22151
rect 25329 22117 25363 22151
rect 26494 22117 26528 22151
rect 32321 22117 32355 22151
rect 32413 22117 32447 22151
rect 37289 22117 37323 22151
rect 3249 22049 3283 22083
rect 5549 22049 5583 22083
rect 6009 22049 6043 22083
rect 6653 22049 6687 22083
rect 6837 22049 6871 22083
rect 7573 22049 7607 22083
rect 7665 22049 7699 22083
rect 8309 22049 8343 22083
rect 9965 22049 9999 22083
rect 10149 22049 10183 22083
rect 10333 22049 10367 22083
rect 10517 22049 10551 22083
rect 11253 22049 11287 22083
rect 12633 22049 12667 22083
rect 15485 22049 15519 22083
rect 15669 22049 15703 22083
rect 16385 22049 16419 22083
rect 18136 22049 18170 22083
rect 18245 22049 18279 22083
rect 18521 22049 18555 22083
rect 20085 22049 20119 22083
rect 21649 22049 21683 22083
rect 22569 22049 22603 22083
rect 25513 22049 25547 22083
rect 26249 22049 26283 22083
rect 28448 22049 28482 22083
rect 30757 22049 30791 22083
rect 30941 22049 30975 22083
rect 31033 22049 31067 22083
rect 31217 22049 31251 22083
rect 32045 22049 32079 22083
rect 32193 22049 32227 22083
rect 32510 22049 32544 22083
rect 33425 22049 33459 22083
rect 33517 22049 33551 22083
rect 33609 22049 33643 22083
rect 33793 22049 33827 22083
rect 34253 22049 34287 22083
rect 36093 22049 36127 22083
rect 36277 22049 36311 22083
rect 36921 22049 36955 22083
rect 37105 22049 37139 22083
rect 55137 22049 55171 22083
rect 55781 22049 55815 22083
rect 57989 22049 58023 22083
rect 1961 21981 1995 22015
rect 2145 21981 2179 22015
rect 10241 21981 10275 22015
rect 16129 21981 16163 22015
rect 18429 21981 18463 22015
rect 20177 21981 20211 22015
rect 21741 21981 21775 22015
rect 22845 21981 22879 22015
rect 28181 21981 28215 22015
rect 56701 21981 56735 22015
rect 56885 21981 56919 22015
rect 57345 21981 57379 22015
rect 3065 21913 3099 21947
rect 4905 21913 4939 21947
rect 12173 21913 12207 21947
rect 15485 21913 15519 21947
rect 27629 21913 27663 21947
rect 31125 21913 31159 21947
rect 32689 21913 32723 21947
rect 54953 21913 54987 21947
rect 58173 21913 58207 21947
rect 2329 21845 2363 21879
rect 7021 21845 7055 21879
rect 8493 21845 8527 21879
rect 10701 21845 10735 21879
rect 13461 21845 13495 21879
rect 14933 21845 14967 21879
rect 17509 21845 17543 21879
rect 17969 21845 18003 21879
rect 20085 21845 20119 21879
rect 20453 21845 20487 21879
rect 21097 21845 21131 21879
rect 24317 21845 24351 21879
rect 29561 21845 29595 21879
rect 33149 21845 33183 21879
rect 34345 21845 34379 21879
rect 55597 21845 55631 21879
rect 1961 21641 1995 21675
rect 2513 21641 2547 21675
rect 4997 21641 5031 21675
rect 6837 21641 6871 21675
rect 14657 21641 14691 21675
rect 19165 21641 19199 21675
rect 21557 21641 21591 21675
rect 24225 21641 24259 21675
rect 29193 21641 29227 21675
rect 29837 21641 29871 21675
rect 30849 21641 30883 21675
rect 33149 21641 33183 21675
rect 33609 21641 33643 21675
rect 35541 21641 35575 21675
rect 55045 21641 55079 21675
rect 57989 21641 58023 21675
rect 4721 21573 4755 21607
rect 13461 21573 13495 21607
rect 15761 21573 15795 21607
rect 56333 21573 56367 21607
rect 7573 21505 7607 21539
rect 10793 21505 10827 21539
rect 12357 21505 12391 21539
rect 13645 21505 13679 21539
rect 20085 21505 20119 21539
rect 23305 21505 23339 21539
rect 24409 21505 24443 21539
rect 28273 21505 28307 21539
rect 55873 21505 55907 21539
rect 2697 21437 2731 21471
rect 4721 21437 4755 21471
rect 4813 21437 4847 21471
rect 5641 21437 5675 21471
rect 7021 21437 7055 21471
rect 7757 21437 7791 21471
rect 8585 21437 8619 21471
rect 8852 21437 8886 21471
rect 10425 21437 10459 21471
rect 10609 21437 10643 21471
rect 10701 21437 10735 21471
rect 10977 21437 11011 21471
rect 12081 21437 12115 21471
rect 12265 21437 12299 21471
rect 12449 21437 12483 21471
rect 12633 21437 12667 21471
rect 13277 21437 13311 21471
rect 13369 21437 13403 21471
rect 13553 21437 13587 21471
rect 14657 21437 14691 21471
rect 14841 21437 14875 21471
rect 15301 21437 15335 21471
rect 15485 21437 15519 21471
rect 15577 21437 15611 21471
rect 15853 21437 15887 21471
rect 17785 21437 17819 21471
rect 19809 21437 19843 21471
rect 19947 21437 19981 21471
rect 20177 21437 20211 21471
rect 20821 21437 20855 21471
rect 21465 21437 21499 21471
rect 22937 21437 22971 21471
rect 23121 21437 23155 21471
rect 23216 21437 23250 21471
rect 23489 21437 23523 21471
rect 24133 21437 24167 21471
rect 25145 21437 25179 21471
rect 26525 21437 26559 21471
rect 26617 21437 26651 21471
rect 26813 21437 26847 21471
rect 26903 21437 26937 21471
rect 27997 21437 28031 21471
rect 28089 21437 28123 21471
rect 28365 21437 28399 21471
rect 29101 21437 29135 21471
rect 29745 21437 29779 21471
rect 30573 21437 30607 21471
rect 30665 21437 30699 21471
rect 30941 21437 30975 21471
rect 31677 21437 31711 21471
rect 33333 21437 33367 21471
rect 33425 21437 33459 21471
rect 33701 21437 33735 21471
rect 34161 21437 34195 21471
rect 36093 21437 36127 21471
rect 36277 21437 36311 21471
rect 55229 21437 55263 21471
rect 55689 21437 55723 21471
rect 56885 21437 56919 21471
rect 57529 21437 57563 21471
rect 57713 21437 57747 21471
rect 1869 21369 1903 21403
rect 3433 21369 3467 21403
rect 3525 21369 3559 21403
rect 4077 21369 4111 21403
rect 18030 21369 18064 21403
rect 25329 21369 25363 21403
rect 27813 21369 27847 21403
rect 31493 21369 31527 21403
rect 34428 21369 34462 21403
rect 36461 21369 36495 21403
rect 5457 21301 5491 21335
rect 7941 21301 7975 21335
rect 9965 21301 9999 21335
rect 11161 21301 11195 21335
rect 12817 21301 12851 21335
rect 19625 21301 19659 21335
rect 20913 21301 20947 21335
rect 23673 21301 23707 21335
rect 24409 21301 24443 21335
rect 25513 21301 25547 21335
rect 26341 21301 26375 21335
rect 30389 21301 30423 21335
rect 57069 21301 57103 21335
rect 3157 21097 3191 21131
rect 4261 21097 4295 21131
rect 6193 21097 6227 21131
rect 8585 21097 8619 21131
rect 17877 21097 17911 21131
rect 18981 21097 19015 21131
rect 20269 21097 20303 21131
rect 22109 21097 22143 21131
rect 23949 21097 23983 21131
rect 25421 21097 25455 21131
rect 26157 21097 26191 21131
rect 33885 21097 33919 21131
rect 34437 21097 34471 21131
rect 55597 21097 55631 21131
rect 1869 21029 1903 21063
rect 7113 21029 7147 21063
rect 7205 21029 7239 21063
rect 9772 21029 9806 21063
rect 11888 21029 11922 21063
rect 22836 21029 22870 21063
rect 32873 21029 32907 21063
rect 2513 20961 2547 20995
rect 3341 20961 3375 20995
rect 4445 20961 4479 20995
rect 5089 20961 5123 20995
rect 5549 20961 5583 20995
rect 6377 20961 6411 20995
rect 8217 20961 8251 20995
rect 8401 20961 8435 20995
rect 9505 20961 9539 20995
rect 11621 20961 11655 20995
rect 13645 20961 13679 20995
rect 13829 20961 13863 20995
rect 15005 20961 15039 20995
rect 17049 20961 17083 20995
rect 17785 20961 17819 20995
rect 17969 20961 18003 20995
rect 18889 20961 18923 20995
rect 19993 20961 20027 20995
rect 20729 20961 20763 20995
rect 20985 20961 21019 20995
rect 22569 20961 22603 20995
rect 25329 20961 25363 20995
rect 26387 20961 26421 20995
rect 26525 20961 26559 20995
rect 26617 20961 26651 20995
rect 27353 20961 27387 20995
rect 28181 20961 28215 20995
rect 28825 20961 28859 20995
rect 29009 20961 29043 20995
rect 29101 20961 29135 20995
rect 29377 20961 29411 20995
rect 31217 20961 31251 20995
rect 31309 20961 31343 20995
rect 31585 20961 31619 20995
rect 32597 20961 32631 20995
rect 32781 20961 32815 20995
rect 32989 20961 33023 20995
rect 33609 20961 33643 20995
rect 34345 20961 34379 20995
rect 36093 20961 36127 20995
rect 36277 20961 36311 20995
rect 36921 20961 36955 20995
rect 55137 20961 55171 20995
rect 55781 20961 55815 20995
rect 56885 20961 56919 20995
rect 57345 20961 57379 20995
rect 57989 20961 58023 20995
rect 58173 20961 58207 20995
rect 7389 20893 7423 20927
rect 13737 20893 13771 20927
rect 14749 20893 14783 20927
rect 20269 20893 20303 20927
rect 26893 20893 26927 20927
rect 29193 20893 29227 20927
rect 33701 20893 33735 20927
rect 33885 20893 33919 20927
rect 56609 20893 56643 20927
rect 56701 20893 56735 20927
rect 4905 20825 4939 20859
rect 20085 20825 20119 20859
rect 27445 20825 27479 20859
rect 31033 20825 31067 20859
rect 33149 20825 33183 20859
rect 36369 20825 36403 20859
rect 1961 20757 1995 20791
rect 2697 20757 2731 20791
rect 5733 20757 5767 20791
rect 10885 20757 10919 20791
rect 13001 20757 13035 20791
rect 16129 20757 16163 20791
rect 17141 20757 17175 20791
rect 26801 20757 26835 20791
rect 28273 20757 28307 20791
rect 29561 20757 29595 20791
rect 31493 20757 31527 20791
rect 37105 20757 37139 20791
rect 1961 20553 1995 20587
rect 8033 20553 8067 20587
rect 12265 20553 12299 20587
rect 13277 20553 13311 20587
rect 14013 20553 14047 20587
rect 14841 20553 14875 20587
rect 23029 20553 23063 20587
rect 24225 20553 24259 20587
rect 25402 20553 25436 20587
rect 25881 20553 25915 20587
rect 26801 20553 26835 20587
rect 29193 20553 29227 20587
rect 31493 20553 31527 20587
rect 34437 20553 34471 20587
rect 34897 20553 34931 20587
rect 55045 20553 55079 20587
rect 56885 20553 56919 20587
rect 4445 20485 4479 20519
rect 13369 20485 13403 20519
rect 19073 20485 19107 20519
rect 24501 20485 24535 20519
rect 25513 20485 25547 20519
rect 31033 20485 31067 20519
rect 5273 20417 5307 20451
rect 6929 20417 6963 20451
rect 8769 20417 8803 20451
rect 10425 20417 10459 20451
rect 10517 20417 10551 20451
rect 13461 20417 13495 20451
rect 14197 20417 14231 20451
rect 16313 20417 16347 20451
rect 19901 20417 19935 20451
rect 21189 20417 21223 20451
rect 23489 20417 23523 20451
rect 25605 20417 25639 20451
rect 27813 20417 27847 20451
rect 31953 20417 31987 20451
rect 36461 20417 36495 20451
rect 2145 20349 2179 20383
rect 4629 20349 4663 20383
rect 5089 20349 5123 20383
rect 8217 20349 8251 20383
rect 8677 20349 8711 20383
rect 8861 20349 8895 20383
rect 9505 20349 9539 20383
rect 10149 20349 10183 20383
rect 10333 20349 10367 20383
rect 10701 20349 10735 20383
rect 12081 20349 12115 20383
rect 13185 20349 13219 20383
rect 13921 20349 13955 20383
rect 14841 20349 14875 20383
rect 15025 20349 15059 20383
rect 15577 20349 15611 20383
rect 16221 20349 16255 20383
rect 17693 20349 17727 20383
rect 19533 20349 19567 20383
rect 19717 20349 19751 20383
rect 19818 20349 19852 20383
rect 20085 20349 20119 20383
rect 20913 20349 20947 20383
rect 21005 20349 21039 20383
rect 21281 20349 21315 20383
rect 23213 20349 23247 20383
rect 23305 20349 23339 20383
rect 23581 20349 23615 20383
rect 24409 20349 24443 20383
rect 24593 20349 24627 20383
rect 24685 20349 24719 20383
rect 26617 20349 26651 20383
rect 29653 20349 29687 20383
rect 29909 20349 29943 20383
rect 31677 20349 31711 20383
rect 31769 20349 31803 20383
rect 32045 20349 32079 20383
rect 33057 20349 33091 20383
rect 33313 20349 33347 20383
rect 34897 20349 34931 20383
rect 35081 20349 35115 20383
rect 36093 20349 36127 20383
rect 36277 20349 36311 20383
rect 54401 20349 54435 20383
rect 55229 20349 55263 20383
rect 55689 20349 55723 20383
rect 57529 20349 57563 20383
rect 57713 20349 57747 20383
rect 2973 20281 3007 20315
rect 3065 20281 3099 20315
rect 3617 20281 3651 20315
rect 7021 20281 7055 20315
rect 7573 20281 7607 20315
rect 17960 20281 17994 20315
rect 20269 20281 20303 20315
rect 25237 20281 25271 20315
rect 26433 20281 26467 20315
rect 28080 20281 28114 20315
rect 56793 20281 56827 20315
rect 5733 20213 5767 20247
rect 9689 20213 9723 20247
rect 10885 20213 10919 20247
rect 14197 20213 14231 20247
rect 15669 20213 15703 20247
rect 20729 20213 20763 20247
rect 55873 20213 55907 20247
rect 58173 20213 58207 20247
rect 8309 20009 8343 20043
rect 1685 19941 1719 19975
rect 2513 19941 2547 19975
rect 4445 19941 4479 19975
rect 7297 19941 7331 19975
rect 9772 19941 9806 19975
rect 15853 19941 15887 19975
rect 16650 19941 16684 19975
rect 18337 19941 18371 19975
rect 25605 19941 25639 19975
rect 26617 19941 26651 19975
rect 27721 19941 27755 19975
rect 28365 19941 28399 19975
rect 54953 19941 54987 19975
rect 55321 19941 55355 19975
rect 57989 19941 58023 19975
rect 5457 19873 5491 19907
rect 8493 19873 8527 19907
rect 9505 19873 9539 19907
rect 11621 19873 11655 19907
rect 11805 19873 11839 19907
rect 11897 19873 11931 19907
rect 12173 19873 12207 19907
rect 12817 19873 12851 19907
rect 13001 19873 13035 19907
rect 13369 19873 13403 19907
rect 14841 19873 14875 19907
rect 15025 19873 15059 19907
rect 15761 19873 15795 19907
rect 15945 19873 15979 19907
rect 18245 19873 18279 19907
rect 18889 19873 18923 19907
rect 20545 19873 20579 19907
rect 20729 19873 20763 19907
rect 21005 19873 21039 19907
rect 21557 19873 21591 19907
rect 21650 19873 21684 19907
rect 21787 19873 21821 19907
rect 21925 19873 21959 19907
rect 22063 19873 22097 19907
rect 22891 19873 22925 19907
rect 23029 19873 23063 19907
rect 23121 19873 23155 19907
rect 23305 19873 23339 19907
rect 23949 19873 23983 19907
rect 24041 19873 24075 19907
rect 24317 19873 24351 19907
rect 25237 19873 25271 19907
rect 25330 19873 25364 19907
rect 25513 19873 25547 19907
rect 25702 19873 25736 19907
rect 26801 19873 26835 19907
rect 26893 19873 26927 19907
rect 27169 19873 27203 19907
rect 27629 19873 27663 19907
rect 28273 19873 28307 19907
rect 28457 19873 28491 19907
rect 28917 19873 28951 19907
rect 31197 19873 31231 19907
rect 32781 19873 32815 19907
rect 32873 19873 32907 19907
rect 53757 19873 53791 19907
rect 58173 19873 58207 19907
rect 2421 19805 2455 19839
rect 4353 19805 4387 19839
rect 4813 19805 4847 19839
rect 5641 19805 5675 19839
rect 7205 19805 7239 19839
rect 7481 19805 7515 19839
rect 11989 19805 12023 19839
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 16405 19805 16439 19839
rect 23765 19805 23799 19839
rect 27077 19805 27111 19839
rect 30941 19805 30975 19839
rect 54309 19805 54343 19839
rect 56701 19805 56735 19839
rect 56885 19805 56919 19839
rect 1869 19737 1903 19771
rect 2973 19737 3007 19771
rect 20825 19737 20859 19771
rect 20913 19737 20947 19771
rect 22201 19737 22235 19771
rect 29009 19737 29043 19771
rect 32321 19737 32355 19771
rect 5825 19669 5859 19703
rect 10885 19669 10919 19703
rect 12357 19669 12391 19703
rect 13553 19669 13587 19703
rect 14841 19669 14875 19703
rect 17785 19669 17819 19703
rect 18981 19669 19015 19703
rect 22661 19669 22695 19703
rect 24225 19669 24259 19703
rect 25881 19669 25915 19703
rect 57345 19669 57379 19703
rect 1961 19465 1995 19499
rect 4537 19465 4571 19499
rect 6837 19465 6871 19499
rect 14197 19465 14231 19499
rect 15117 19465 15151 19499
rect 17325 19465 17359 19499
rect 19073 19465 19107 19499
rect 19533 19465 19567 19499
rect 20177 19465 20211 19499
rect 21281 19465 21315 19499
rect 24225 19465 24259 19499
rect 24685 19465 24719 19499
rect 26709 19465 26743 19499
rect 28733 19465 28767 19499
rect 29929 19465 29963 19499
rect 56793 19465 56827 19499
rect 57253 19465 57287 19499
rect 14105 19397 14139 19431
rect 16129 19397 16163 19431
rect 9781 19329 9815 19363
rect 10609 19329 10643 19363
rect 14289 19329 14323 19363
rect 15577 19329 15611 19363
rect 16773 19329 16807 19363
rect 17785 19329 17819 19363
rect 2145 19261 2179 19295
rect 2605 19261 2639 19295
rect 3801 19261 3835 19295
rect 4537 19261 4571 19295
rect 4721 19261 4755 19295
rect 5365 19261 5399 19295
rect 7021 19261 7055 19295
rect 9965 19261 9999 19295
rect 10793 19261 10827 19295
rect 12173 19261 12207 19295
rect 12440 19261 12474 19295
rect 14013 19261 14047 19295
rect 15301 19261 15335 19295
rect 15393 19261 15427 19295
rect 15669 19261 15703 19295
rect 16129 19261 16163 19295
rect 16313 19261 16347 19295
rect 7941 19193 7975 19227
rect 8033 19193 8067 19227
rect 8953 19193 8987 19227
rect 17509 19261 17543 19295
rect 17601 19261 17635 19295
rect 17877 19261 17911 19295
rect 18429 19261 18463 19295
rect 18521 19261 18555 19295
rect 19257 19261 19291 19295
rect 19379 19261 19413 19295
rect 19625 19261 19659 19295
rect 20085 19261 20119 19295
rect 21189 19261 21223 19295
rect 23029 19261 23063 19295
rect 23489 19261 23523 19295
rect 24409 19261 24443 19295
rect 24501 19261 24535 19295
rect 24777 19261 24811 19295
rect 25605 19261 25639 19295
rect 25973 19261 26007 19295
rect 26617 19261 26651 19295
rect 27813 19261 27847 19295
rect 28641 19261 28675 19295
rect 29285 19261 29319 19295
rect 29377 19261 29411 19295
rect 29929 19261 29963 19295
rect 30113 19261 30147 19295
rect 30665 19261 30699 19295
rect 31493 19261 31527 19295
rect 56149 19261 56183 19295
rect 57437 19261 57471 19295
rect 57989 19261 58023 19295
rect 58173 19261 58207 19295
rect 23765 19193 23799 19227
rect 25789 19193 25823 19227
rect 25881 19193 25915 19227
rect 30757 19193 30791 19227
rect 2789 19125 2823 19159
rect 3617 19125 3651 19159
rect 5181 19125 5215 19159
rect 10149 19125 10183 19159
rect 10977 19125 11011 19159
rect 13553 19125 13587 19159
rect 16773 19125 16807 19159
rect 26157 19125 26191 19159
rect 27905 19125 27939 19159
rect 31585 19125 31619 19159
rect 55965 19125 55999 19159
rect 2881 18921 2915 18955
rect 5825 18921 5859 18955
rect 6377 18921 6411 18955
rect 7021 18921 7055 18955
rect 7757 18921 7791 18955
rect 10241 18921 10275 18955
rect 12541 18921 12575 18955
rect 16129 18921 16163 18955
rect 16681 18921 16715 18955
rect 19073 18921 19107 18955
rect 20085 18921 20119 18955
rect 20637 18921 20671 18955
rect 28917 18921 28951 18955
rect 29469 18921 29503 18955
rect 31033 18921 31067 18955
rect 2053 18853 2087 18887
rect 11428 18853 11462 18887
rect 14994 18853 15028 18887
rect 22284 18853 22318 18887
rect 1869 18785 1903 18819
rect 3065 18785 3099 18819
rect 5641 18785 5675 18819
rect 6285 18785 6319 18819
rect 6469 18785 6503 18819
rect 6929 18785 6963 18819
rect 7113 18785 7147 18819
rect 7573 18785 7607 18819
rect 8217 18785 8251 18819
rect 9873 18785 9907 18819
rect 10057 18785 10091 18819
rect 13001 18785 13035 18819
rect 13185 18785 13219 18819
rect 13645 18785 13679 18819
rect 14749 18785 14783 18819
rect 16589 18785 16623 18819
rect 17693 18785 17727 18819
rect 17960 18785 17994 18819
rect 19993 18785 20027 18819
rect 20821 18785 20855 18819
rect 21281 18785 21315 18819
rect 24041 18785 24075 18819
rect 25743 18785 25777 18819
rect 25862 18785 25896 18819
rect 25994 18785 26028 18819
rect 26157 18785 26191 18819
rect 26617 18785 26651 18819
rect 26709 18785 26743 18819
rect 27804 18785 27838 18819
rect 29377 18785 29411 18819
rect 29561 18785 29595 18819
rect 30941 18785 30975 18819
rect 31125 18785 31159 18819
rect 55597 18785 55631 18819
rect 57989 18785 58023 18819
rect 11161 18717 11195 18751
rect 21005 18717 21039 18751
rect 21097 18717 21131 18751
rect 22017 18717 22051 18751
rect 26893 18717 26927 18751
rect 27537 18717 27571 18751
rect 20913 18649 20947 18683
rect 58173 18649 58207 18683
rect 8401 18581 8435 18615
rect 13001 18581 13035 18615
rect 13829 18581 13863 18615
rect 23397 18581 23431 18615
rect 24133 18581 24167 18615
rect 25513 18581 25547 18615
rect 26801 18581 26835 18615
rect 57437 18581 57471 18615
rect 5733 18377 5767 18411
rect 16129 18377 16163 18411
rect 17325 18377 17359 18411
rect 18981 18377 19015 18411
rect 26065 18377 26099 18411
rect 28457 18377 28491 18411
rect 29285 18377 29319 18411
rect 57989 18377 58023 18411
rect 21465 18309 21499 18343
rect 27905 18309 27939 18343
rect 56885 18309 56919 18343
rect 8677 18241 8711 18275
rect 9965 18241 9999 18275
rect 10793 18241 10827 18275
rect 21005 18241 21039 18275
rect 23397 18241 23431 18275
rect 57529 18241 57563 18275
rect 57713 18241 57747 18275
rect 5733 18173 5767 18207
rect 5917 18173 5951 18207
rect 10149 18173 10183 18207
rect 10977 18173 11011 18207
rect 12345 18173 12379 18207
rect 12541 18173 12575 18207
rect 13001 18173 13035 18207
rect 13185 18173 13219 18207
rect 15209 18173 15243 18207
rect 15393 18173 15427 18207
rect 16129 18173 16163 18207
rect 16313 18173 16347 18207
rect 17325 18173 17359 18207
rect 17509 18173 17543 18207
rect 18337 18173 18371 18207
rect 18981 18173 19015 18207
rect 19165 18173 19199 18207
rect 19717 18173 19751 18207
rect 19901 18173 19935 18207
rect 20361 18173 20395 18207
rect 20545 18173 20579 18207
rect 21189 18173 21223 18207
rect 21557 18173 21591 18207
rect 22845 18173 22879 18207
rect 23213 18173 23247 18207
rect 23949 18173 23983 18207
rect 26065 18173 26099 18207
rect 26249 18173 26283 18207
rect 27813 18173 27847 18207
rect 28457 18173 28491 18207
rect 28641 18173 28675 18207
rect 29285 18173 29319 18207
rect 29469 18173 29503 18207
rect 56241 18173 56275 18207
rect 57069 18173 57103 18207
rect 8401 18105 8435 18139
rect 8493 18105 8527 18139
rect 12449 18105 12483 18139
rect 13093 18105 13127 18139
rect 13737 18105 13771 18139
rect 13829 18105 13863 18139
rect 14749 18105 14783 18139
rect 18429 18105 18463 18139
rect 20453 18105 20487 18139
rect 24216 18105 24250 18139
rect 10333 18037 10367 18071
rect 11161 18037 11195 18071
rect 15301 18037 15335 18071
rect 19809 18037 19843 18071
rect 25329 18037 25363 18071
rect 1961 17833 1995 17867
rect 14841 17833 14875 17867
rect 16037 17833 16071 17867
rect 21373 17833 21407 17867
rect 21925 17833 21959 17867
rect 24133 17833 24167 17867
rect 25329 17833 25363 17867
rect 27261 17833 27295 17867
rect 1869 17765 1903 17799
rect 10609 17765 10643 17799
rect 20238 17765 20272 17799
rect 26126 17765 26160 17799
rect 56609 17765 56643 17799
rect 58173 17765 58207 17799
rect 12081 17697 12115 17731
rect 13829 17697 13863 17731
rect 14749 17697 14783 17731
rect 14933 17697 14967 17731
rect 15577 17697 15611 17731
rect 16221 17697 16255 17731
rect 19993 17697 20027 17731
rect 21833 17697 21867 17731
rect 22845 17697 22879 17731
rect 23305 17697 23339 17731
rect 24041 17697 24075 17731
rect 25237 17697 25271 17731
rect 56701 17697 56735 17731
rect 57345 17697 57379 17731
rect 57989 17697 58023 17731
rect 10517 17629 10551 17663
rect 10793 17629 10827 17663
rect 23581 17629 23615 17663
rect 25881 17629 25915 17663
rect 56885 17629 56919 17663
rect 15393 17561 15427 17595
rect 12265 17493 12299 17527
rect 13645 17493 13679 17527
rect 15025 17289 15059 17323
rect 21373 17289 21407 17323
rect 24777 17289 24811 17323
rect 55413 17289 55447 17323
rect 56333 17221 56367 17255
rect 56885 17221 56919 17255
rect 10333 17153 10367 17187
rect 10609 17153 10643 17187
rect 12173 17153 12207 17187
rect 13737 17153 13771 17187
rect 23397 17153 23431 17187
rect 57713 17153 57747 17187
rect 1869 17085 1903 17119
rect 9781 17085 9815 17119
rect 14841 17085 14875 17119
rect 21281 17085 21315 17119
rect 22845 17085 22879 17119
rect 23213 17085 23247 17119
rect 24133 17085 24167 17119
rect 55597 17085 55631 17119
rect 57069 17085 57103 17119
rect 57529 17085 57563 17119
rect 2053 17017 2087 17051
rect 10425 17017 10459 17051
rect 12265 17017 12299 17051
rect 13185 17017 13219 17051
rect 13829 17017 13863 17051
rect 14381 17017 14415 17051
rect 56149 17017 56183 17051
rect 9597 16949 9631 16983
rect 58173 16949 58207 16983
rect 10609 16745 10643 16779
rect 13829 16745 13863 16779
rect 24133 16745 24167 16779
rect 55597 16745 55631 16779
rect 23581 16677 23615 16711
rect 57989 16677 58023 16711
rect 58173 16677 58207 16711
rect 10793 16609 10827 16643
rect 13645 16609 13679 16643
rect 22845 16609 22879 16643
rect 23305 16609 23339 16643
rect 24041 16609 24075 16643
rect 24225 16609 24259 16643
rect 55781 16609 55815 16643
rect 56793 16609 56827 16643
rect 56977 16609 57011 16643
rect 57437 16609 57471 16643
rect 56977 16201 57011 16235
rect 55689 16133 55723 16167
rect 2053 16065 2087 16099
rect 1869 15997 1903 16031
rect 14749 15997 14783 16031
rect 54861 15997 54895 16031
rect 56149 15997 56183 16031
rect 15025 15929 15059 15963
rect 56885 15929 56919 15963
rect 57989 15929 58023 15963
rect 56333 15861 56367 15895
rect 58081 15861 58115 15895
rect 58173 15657 58207 15691
rect 55781 15521 55815 15555
rect 56885 15521 56919 15555
rect 55137 15453 55171 15487
rect 57529 15453 57563 15487
rect 57713 15453 57747 15487
rect 55597 15385 55631 15419
rect 56977 15317 57011 15351
rect 1961 15113 1995 15147
rect 56333 15113 56367 15147
rect 56425 15113 56459 15147
rect 56977 15113 57011 15147
rect 55965 15045 55999 15079
rect 58173 15045 58207 15079
rect 56793 14977 56827 15011
rect 1869 14909 1903 14943
rect 56149 14909 56183 14943
rect 56333 14909 56367 14943
rect 56609 14909 56643 14943
rect 57989 14909 58023 14943
rect 56793 14569 56827 14603
rect 1869 14501 1903 14535
rect 57621 14501 57655 14535
rect 55597 14433 55631 14467
rect 56977 14433 57011 14467
rect 57529 14365 57563 14399
rect 57805 14365 57839 14399
rect 1961 14229 1995 14263
rect 55781 14025 55815 14059
rect 56241 13957 56275 13991
rect 56885 13957 56919 13991
rect 57713 13889 57747 13923
rect 56425 13821 56459 13855
rect 57069 13821 57103 13855
rect 57529 13821 57563 13855
rect 58173 13685 58207 13719
rect 58081 13481 58115 13515
rect 1869 13413 1903 13447
rect 57989 13413 58023 13447
rect 55781 13345 55815 13379
rect 56885 13345 56919 13379
rect 56701 13277 56735 13311
rect 2053 13209 2087 13243
rect 56609 13209 56643 13243
rect 57253 13141 57287 13175
rect 56241 12937 56275 12971
rect 57345 12937 57379 12971
rect 55413 12733 55447 12767
rect 56057 12733 56091 12767
rect 57253 12733 57287 12767
rect 57989 12665 58023 12699
rect 58081 12597 58115 12631
rect 1961 12393 1995 12427
rect 58173 12393 58207 12427
rect 1869 12325 1903 12359
rect 56885 12257 56919 12291
rect 57529 12189 57563 12223
rect 57713 12189 57747 12223
rect 56977 12053 57011 12087
rect 55597 11849 55631 11883
rect 57713 11849 57747 11883
rect 56701 11781 56735 11815
rect 56241 11713 56275 11747
rect 57345 11713 57379 11747
rect 57529 11713 57563 11747
rect 1869 11645 1903 11679
rect 56885 11645 56919 11679
rect 1961 11509 1995 11543
rect 57253 11305 57287 11339
rect 55597 11169 55631 11203
rect 57437 11169 57471 11203
rect 57989 11169 58023 11203
rect 58173 11033 58207 11067
rect 57989 10761 58023 10795
rect 56425 10625 56459 10659
rect 57529 10625 57563 10659
rect 1869 10557 1903 10591
rect 57069 10557 57103 10591
rect 57713 10557 57747 10591
rect 2053 10489 2087 10523
rect 56885 10421 56919 10455
rect 57253 10217 57287 10251
rect 55597 10081 55631 10115
rect 57437 10081 57471 10115
rect 57989 10081 58023 10115
rect 58173 9945 58207 9979
rect 2053 9605 2087 9639
rect 57621 9605 57655 9639
rect 1869 9469 1903 9503
rect 55689 9469 55723 9503
rect 56517 9469 56551 9503
rect 56977 9469 57011 9503
rect 57161 9469 57195 9503
rect 56885 9129 56919 9163
rect 1869 9061 1903 9095
rect 55781 8993 55815 9027
rect 57069 8993 57103 9027
rect 57713 8993 57747 9027
rect 55137 8925 55171 8959
rect 57529 8925 57563 8959
rect 1961 8789 1995 8823
rect 57989 8789 58023 8823
rect 56149 8585 56183 8619
rect 55321 8517 55355 8551
rect 58173 8517 58207 8551
rect 54861 8449 54895 8483
rect 57437 8449 57471 8483
rect 55505 8381 55539 8415
rect 55965 8381 55999 8415
rect 57989 8381 58023 8415
rect 57253 8313 57287 8347
rect 1869 7973 1903 8007
rect 53665 7905 53699 7939
rect 57161 7905 57195 7939
rect 57345 7905 57379 7939
rect 2053 7769 2087 7803
rect 54493 7769 54527 7803
rect 57529 7769 57563 7803
rect 55137 7701 55171 7735
rect 55781 7701 55815 7735
rect 55781 7429 55815 7463
rect 56609 7361 56643 7395
rect 57529 7361 57563 7395
rect 52929 7293 52963 7327
rect 54677 7293 54711 7327
rect 55321 7293 55355 7327
rect 55965 7293 55999 7327
rect 56425 7293 56459 7327
rect 57713 7293 57747 7327
rect 57069 7157 57103 7191
rect 58173 7157 58207 7191
rect 1869 6817 1903 6851
rect 51733 6817 51767 6851
rect 52561 6817 52595 6851
rect 55137 6817 55171 6851
rect 55781 6817 55815 6851
rect 57989 6817 58023 6851
rect 58173 6817 58207 6851
rect 2053 6749 2087 6783
rect 53205 6749 53239 6783
rect 56793 6749 56827 6783
rect 56977 6749 57011 6783
rect 55597 6681 55631 6715
rect 53849 6613 53883 6647
rect 54493 6613 54527 6647
rect 54953 6613 54987 6647
rect 57161 6613 57195 6647
rect 55413 6409 55447 6443
rect 56333 6341 56367 6375
rect 56793 6273 56827 6307
rect 51641 6205 51675 6239
rect 52469 6205 52503 6239
rect 53113 6205 53147 6239
rect 54217 6205 54251 6239
rect 54953 6205 54987 6239
rect 55597 6205 55631 6239
rect 56149 6205 56183 6239
rect 56977 6205 57011 6239
rect 57437 6137 57471 6171
rect 57989 6137 58023 6171
rect 54769 6069 54803 6103
rect 58081 6069 58115 6103
rect 1961 5865 1995 5899
rect 54861 5865 54895 5899
rect 1869 5797 1903 5831
rect 55781 5797 55815 5831
rect 58173 5797 58207 5831
rect 52469 5729 52503 5763
rect 53757 5729 53791 5763
rect 54401 5729 54435 5763
rect 55045 5729 55079 5763
rect 55597 5729 55631 5763
rect 56701 5729 56735 5763
rect 57989 5729 58023 5763
rect 51825 5661 51859 5695
rect 56885 5661 56919 5695
rect 54217 5593 54251 5627
rect 53113 5525 53147 5559
rect 53573 5525 53607 5559
rect 57069 5525 57103 5559
rect 54217 5321 54251 5355
rect 54953 5185 54987 5219
rect 57529 5185 57563 5219
rect 1869 5117 1903 5151
rect 49801 5117 49835 5151
rect 50629 5117 50663 5151
rect 51641 5117 51675 5151
rect 52469 5117 52503 5151
rect 53113 5117 53147 5151
rect 54033 5117 54067 5151
rect 54769 5117 54803 5151
rect 56885 5117 56919 5151
rect 57713 5117 57747 5151
rect 55873 5049 55907 5083
rect 1961 4981 1995 5015
rect 52929 4981 52963 5015
rect 55965 4981 55999 5015
rect 56977 4981 57011 5015
rect 58173 4981 58207 5015
rect 53757 4709 53791 4743
rect 54493 4709 54527 4743
rect 56885 4709 56919 4743
rect 37933 4641 37967 4675
rect 48973 4641 49007 4675
rect 51917 4641 51951 4675
rect 52561 4641 52595 4675
rect 53205 4641 53239 4675
rect 55321 4641 55355 4675
rect 57713 4641 57747 4675
rect 55137 4573 55171 4607
rect 57529 4573 57563 4607
rect 46397 4505 46431 4539
rect 53021 4505 53055 4539
rect 32965 4437 32999 4471
rect 36093 4437 36127 4471
rect 37013 4437 37047 4471
rect 37749 4437 37783 4471
rect 38577 4437 38611 4471
rect 39221 4437 39255 4471
rect 39865 4437 39899 4471
rect 41521 4437 41555 4471
rect 42349 4437 42383 4471
rect 43453 4437 43487 4471
rect 47041 4437 47075 4471
rect 48053 4437 48087 4471
rect 48789 4437 48823 4471
rect 49617 4437 49651 4471
rect 50261 4437 50295 4471
rect 51733 4437 51767 4471
rect 52377 4437 52411 4471
rect 53849 4437 53883 4471
rect 54585 4437 54619 4471
rect 55597 4437 55631 4471
rect 56977 4437 57011 4471
rect 57989 4437 58023 4471
rect 34805 4165 34839 4199
rect 45109 4165 45143 4199
rect 45753 4165 45787 4199
rect 2053 4097 2087 4131
rect 49893 4097 49927 4131
rect 56425 4097 56459 4131
rect 56885 4097 56919 4131
rect 30297 4029 30331 4063
rect 32137 4029 32171 4063
rect 33241 4029 33275 4063
rect 34161 4029 34195 4063
rect 35449 4029 35483 4063
rect 36093 4029 36127 4063
rect 37381 4029 37415 4063
rect 38853 4029 38887 4063
rect 39957 4029 39991 4063
rect 40601 4029 40635 4063
rect 41245 4029 41279 4063
rect 42073 4029 42107 4063
rect 43729 4029 43763 4063
rect 44465 4029 44499 4063
rect 46949 4029 46983 4063
rect 47685 4029 47719 4063
rect 49157 4029 49191 4063
rect 50353 4029 50387 4063
rect 51181 4029 51215 4063
rect 51825 4029 51859 4063
rect 52469 4029 52503 4063
rect 53113 4029 53147 4063
rect 55781 4029 55815 4063
rect 56241 4029 56275 4063
rect 57989 4029 58023 4063
rect 1869 3961 1903 3995
rect 49709 3961 49743 3995
rect 54125 3961 54159 3995
rect 54953 3961 54987 3995
rect 58173 3961 58207 3995
rect 33057 3893 33091 3927
rect 33977 3893 34011 3927
rect 36277 3893 36311 3927
rect 37197 3893 37231 3927
rect 38669 3893 38703 3927
rect 39773 3893 39807 3927
rect 40417 3893 40451 3927
rect 41889 3893 41923 3927
rect 43545 3893 43579 3927
rect 44281 3893 44315 3927
rect 46765 3893 46799 3927
rect 47869 3893 47903 3927
rect 48973 3893 49007 3927
rect 50537 3893 50571 3927
rect 50997 3893 51031 3927
rect 51641 3893 51675 3927
rect 52285 3893 52319 3927
rect 52929 3893 52963 3927
rect 54217 3893 54251 3927
rect 55045 3893 55079 3927
rect 55597 3893 55631 3927
rect 12357 3689 12391 3723
rect 36921 3689 36955 3723
rect 43913 3689 43947 3723
rect 53757 3689 53791 3723
rect 56701 3689 56735 3723
rect 1869 3621 1903 3655
rect 11253 3621 11287 3655
rect 11345 3621 11379 3655
rect 55597 3621 55631 3655
rect 2881 3553 2915 3587
rect 12541 3553 12575 3587
rect 30665 3553 30699 3587
rect 32321 3553 32355 3587
rect 32873 3553 32907 3587
rect 33793 3553 33827 3587
rect 34805 3553 34839 3587
rect 35817 3553 35851 3587
rect 36737 3553 36771 3587
rect 37473 3553 37507 3587
rect 38393 3553 38427 3587
rect 39313 3553 39347 3587
rect 41061 3553 41095 3587
rect 42441 3553 42475 3587
rect 42993 3553 43027 3587
rect 43729 3553 43763 3587
rect 44741 3553 44775 3587
rect 46397 3553 46431 3587
rect 47041 3553 47075 3587
rect 47593 3553 47627 3587
rect 48513 3553 48547 3587
rect 49801 3553 49835 3587
rect 50353 3553 50387 3587
rect 51549 3553 51583 3587
rect 52285 3553 52319 3587
rect 53113 3553 53147 3587
rect 53297 3553 53331 3587
rect 54309 3553 54343 3587
rect 56885 3553 56919 3587
rect 57529 3553 57563 3587
rect 11529 3485 11563 3519
rect 57345 3485 57379 3519
rect 46213 3417 46247 3451
rect 55781 3417 55815 3451
rect 1961 3349 1995 3383
rect 29469 3349 29503 3383
rect 30481 3349 30515 3383
rect 31309 3349 31343 3383
rect 32137 3349 32171 3383
rect 32965 3349 32999 3383
rect 33885 3349 33919 3383
rect 34621 3349 34655 3383
rect 35909 3349 35943 3383
rect 37565 3349 37599 3383
rect 38485 3349 38519 3383
rect 39405 3349 39439 3383
rect 41153 3349 41187 3383
rect 42257 3349 42291 3383
rect 43085 3349 43119 3383
rect 44557 3349 44591 3383
rect 46857 3349 46891 3383
rect 47685 3349 47719 3383
rect 48605 3349 48639 3383
rect 49617 3349 49651 3383
rect 50445 3349 50479 3383
rect 51641 3349 51675 3383
rect 52377 3349 52411 3383
rect 54401 3349 54435 3383
rect 57989 3349 58023 3383
rect 1593 3145 1627 3179
rect 3065 3145 3099 3179
rect 33425 3145 33459 3179
rect 35449 3145 35483 3179
rect 38669 3145 38703 3179
rect 39773 3145 39807 3179
rect 47593 3145 47627 3179
rect 51457 3145 51491 3179
rect 52837 3145 52871 3179
rect 54677 3145 54711 3179
rect 55781 3145 55815 3179
rect 56701 3145 56735 3179
rect 57897 3077 57931 3111
rect 30021 3009 30055 3043
rect 30205 3009 30239 3043
rect 33241 3009 33275 3043
rect 34989 3009 35023 3043
rect 38301 3009 38335 3043
rect 39405 3009 39439 3043
rect 39589 3009 39623 3043
rect 40693 3009 40727 3043
rect 43545 3009 43579 3043
rect 43729 3009 43763 3043
rect 45661 3009 45695 3043
rect 47133 3009 47167 3043
rect 48973 3009 49007 3043
rect 50813 3009 50847 3043
rect 50997 3009 51031 3043
rect 52193 3009 52227 3043
rect 54033 3009 54067 3043
rect 54217 3009 54251 3043
rect 55137 3009 55171 3043
rect 56241 3009 56275 3043
rect 56425 3009 56459 3043
rect 57713 3009 57747 3043
rect 1409 2941 1443 2975
rect 2237 2941 2271 2975
rect 3617 2941 3651 2975
rect 4261 2941 4295 2975
rect 28089 2941 28123 2975
rect 28733 2941 28767 2975
rect 29561 2941 29595 2975
rect 31309 2941 31343 2975
rect 33057 2941 33091 2975
rect 34345 2941 34379 2975
rect 34805 2941 34839 2975
rect 36185 2941 36219 2975
rect 38485 2941 38519 2975
rect 40509 2941 40543 2975
rect 46949 2941 46983 2975
rect 48789 2941 48823 2975
rect 52377 2941 52411 2975
rect 55321 2941 55355 2975
rect 57529 2941 57563 2975
rect 2421 2873 2455 2907
rect 2973 2873 3007 2907
rect 30665 2873 30699 2907
rect 31953 2873 31987 2907
rect 36001 2873 36035 2907
rect 36737 2873 36771 2907
rect 41153 2873 41187 2907
rect 41705 2873 41739 2907
rect 42441 2873 42475 2907
rect 44189 2873 44223 2907
rect 44741 2873 44775 2907
rect 45477 2873 45511 2907
rect 46213 2873 46247 2907
rect 49433 2873 49467 2907
rect 49985 2873 50019 2907
rect 29377 2805 29411 2839
rect 31125 2805 31159 2839
rect 32045 2805 32079 2839
rect 34161 2805 34195 2839
rect 36829 2805 36863 2839
rect 41797 2805 41831 2839
rect 42533 2805 42567 2839
rect 44833 2805 44867 2839
rect 46305 2805 46339 2839
rect 50077 2805 50111 2839
rect 31585 2601 31619 2635
rect 35357 2601 35391 2635
rect 36921 2601 36955 2635
rect 40141 2601 40175 2635
rect 42257 2601 42291 2635
rect 44925 2601 44959 2635
rect 46029 2601 46063 2635
rect 48697 2601 48731 2635
rect 50261 2601 50295 2635
rect 56701 2601 56735 2635
rect 2789 2533 2823 2567
rect 28457 2533 28491 2567
rect 29745 2533 29779 2567
rect 32137 2533 32171 2567
rect 47593 2533 47627 2567
rect 50813 2533 50847 2567
rect 53849 2533 53883 2567
rect 54033 2533 54067 2567
rect 55413 2533 55447 2567
rect 57989 2533 58023 2567
rect 1685 2465 1719 2499
rect 4261 2465 4295 2499
rect 5089 2465 5123 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 7849 2465 7883 2499
rect 8493 2465 8527 2499
rect 9689 2465 9723 2499
rect 10609 2465 10643 2499
rect 12265 2465 12299 2499
rect 12909 2465 12943 2499
rect 13553 2465 13587 2499
rect 14933 2465 14967 2499
rect 15577 2465 15611 2499
rect 16221 2465 16255 2499
rect 17601 2465 17635 2499
rect 18245 2465 18279 2499
rect 18889 2465 18923 2499
rect 20269 2465 20303 2499
rect 20913 2465 20947 2499
rect 21649 2465 21683 2499
rect 22937 2465 22971 2499
rect 23581 2465 23615 2499
rect 24409 2465 24443 2499
rect 25605 2465 25639 2499
rect 26249 2465 26283 2499
rect 27169 2465 27203 2499
rect 29101 2465 29135 2499
rect 29285 2465 29319 2499
rect 30941 2465 30975 2499
rect 31125 2465 31159 2499
rect 33609 2465 33643 2499
rect 33793 2465 33827 2499
rect 34713 2465 34747 2499
rect 36461 2465 36495 2499
rect 37381 2465 37415 2499
rect 37565 2465 37599 2499
rect 39497 2465 39531 2499
rect 39681 2465 39715 2499
rect 41613 2465 41647 2499
rect 41797 2465 41831 2499
rect 42717 2465 42751 2499
rect 42901 2465 42935 2499
rect 44281 2465 44315 2499
rect 44465 2465 44499 2499
rect 45385 2465 45419 2499
rect 46949 2465 46983 2499
rect 47133 2465 47167 2499
rect 48053 2465 48087 2499
rect 49801 2465 49835 2499
rect 52285 2465 52319 2499
rect 56057 2465 56091 2499
rect 34897 2397 34931 2431
rect 36277 2397 36311 2431
rect 45569 2397 45603 2431
rect 48237 2397 48271 2431
rect 49617 2397 49651 2431
rect 52469 2397 52503 2431
rect 56241 2397 56275 2431
rect 2237 2329 2271 2363
rect 28641 2329 28675 2363
rect 33977 2329 34011 2363
rect 37749 2329 37783 2363
rect 43085 2329 43119 2363
rect 52653 2329 52687 2363
rect 55597 2329 55631 2363
rect 2881 2261 2915 2295
rect 32229 2261 32263 2295
rect 50905 2261 50939 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 55306 58624 55312 58676
rect 55364 58664 55370 58676
rect 56410 58664 56416 58676
rect 55364 58636 56416 58664
rect 55364 58624 55370 58636
rect 56410 58624 56416 58636
rect 56468 58624 56474 58676
rect 53742 58012 53748 58064
rect 53800 58052 53806 58064
rect 56502 58052 56508 58064
rect 53800 58024 56508 58052
rect 53800 58012 53806 58024
rect 56502 58012 56508 58024
rect 56560 58012 56566 58064
rect 27246 57876 27252 57928
rect 27304 57916 27310 57928
rect 34238 57916 34244 57928
rect 27304 57888 34244 57916
rect 27304 57876 27310 57888
rect 34238 57876 34244 57888
rect 34296 57876 34302 57928
rect 27982 57808 27988 57860
rect 28040 57848 28046 57860
rect 29822 57848 29828 57860
rect 28040 57820 29828 57848
rect 28040 57808 28046 57820
rect 29822 57808 29828 57820
rect 29880 57808 29886 57860
rect 30374 57808 30380 57860
rect 30432 57848 30438 57860
rect 37090 57848 37096 57860
rect 30432 57820 37096 57848
rect 30432 57808 30438 57820
rect 37090 57808 37096 57820
rect 37148 57808 37154 57860
rect 26418 57740 26424 57792
rect 26476 57780 26482 57792
rect 32306 57780 32312 57792
rect 26476 57752 32312 57780
rect 26476 57740 26482 57752
rect 32306 57740 32312 57752
rect 32364 57740 32370 57792
rect 33502 57740 33508 57792
rect 33560 57780 33566 57792
rect 36262 57780 36268 57792
rect 33560 57752 36268 57780
rect 33560 57740 33566 57752
rect 36262 57740 36268 57752
rect 36320 57740 36326 57792
rect 1104 57690 58880 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 58880 57690
rect 1104 57616 58880 57638
rect 3237 57579 3295 57585
rect 3237 57545 3249 57579
rect 3283 57576 3295 57579
rect 4062 57576 4068 57588
rect 3283 57548 4068 57576
rect 3283 57545 3295 57548
rect 3237 57539 3295 57545
rect 4062 57536 4068 57548
rect 4120 57536 4126 57588
rect 4614 57536 4620 57588
rect 4672 57576 4678 57588
rect 4672 57548 22094 57576
rect 4672 57536 4678 57548
rect 2041 57511 2099 57517
rect 2041 57477 2053 57511
rect 2087 57508 2099 57511
rect 2774 57508 2780 57520
rect 2087 57480 2780 57508
rect 2087 57477 2099 57480
rect 2041 57471 2099 57477
rect 2774 57468 2780 57480
rect 2832 57468 2838 57520
rect 10413 57511 10471 57517
rect 10413 57477 10425 57511
rect 10459 57508 10471 57511
rect 11974 57508 11980 57520
rect 10459 57480 11980 57508
rect 10459 57477 10471 57480
rect 10413 57471 10471 57477
rect 11974 57468 11980 57480
rect 12032 57468 12038 57520
rect 12158 57468 12164 57520
rect 12216 57508 12222 57520
rect 22066 57508 22094 57548
rect 24026 57536 24032 57588
rect 24084 57576 24090 57588
rect 24084 57548 27016 57576
rect 24084 57536 24090 57548
rect 26142 57508 26148 57520
rect 12216 57480 13492 57508
rect 22066 57480 26148 57508
rect 12216 57468 12222 57480
rect 6638 57400 6644 57452
rect 6696 57440 6702 57452
rect 11992 57440 12020 57468
rect 12713 57443 12771 57449
rect 12713 57440 12725 57443
rect 6696 57412 7604 57440
rect 11992 57412 12725 57440
rect 6696 57400 6702 57412
rect 4246 57372 4252 57384
rect 4207 57344 4252 57372
rect 4246 57332 4252 57344
rect 4304 57332 4310 57384
rect 4433 57375 4491 57381
rect 4433 57341 4445 57375
rect 4479 57372 4491 57375
rect 4798 57372 4804 57384
rect 4479 57344 4804 57372
rect 4479 57341 4491 57344
rect 4433 57335 4491 57341
rect 4798 57332 4804 57344
rect 4856 57332 4862 57384
rect 5074 57332 5080 57384
rect 5132 57372 5138 57384
rect 5353 57375 5411 57381
rect 5353 57372 5365 57375
rect 5132 57344 5365 57372
rect 5132 57332 5138 57344
rect 5353 57341 5365 57344
rect 5399 57341 5411 57375
rect 5353 57335 5411 57341
rect 5902 57332 5908 57384
rect 5960 57372 5966 57384
rect 7576 57381 7604 57412
rect 12713 57409 12725 57412
rect 12759 57409 12771 57443
rect 12713 57403 12771 57409
rect 6917 57375 6975 57381
rect 6917 57372 6929 57375
rect 5960 57344 6929 57372
rect 5960 57332 5966 57344
rect 6917 57341 6929 57344
rect 6963 57341 6975 57375
rect 6917 57335 6975 57341
rect 7561 57375 7619 57381
rect 7561 57341 7573 57375
rect 7607 57341 7619 57375
rect 7561 57335 7619 57341
rect 8205 57375 8263 57381
rect 8205 57341 8217 57375
rect 8251 57341 8263 57375
rect 8205 57335 8263 57341
rect 1854 57304 1860 57316
rect 1815 57276 1860 57304
rect 1854 57264 1860 57276
rect 1912 57264 1918 57316
rect 3145 57307 3203 57313
rect 3145 57273 3157 57307
rect 3191 57304 3203 57307
rect 4893 57307 4951 57313
rect 4893 57304 4905 57307
rect 3191 57276 4905 57304
rect 3191 57273 3203 57276
rect 3145 57267 3203 57273
rect 4893 57273 4905 57276
rect 4939 57273 4951 57307
rect 4893 57267 4951 57273
rect 7466 57264 7472 57316
rect 7524 57304 7530 57316
rect 8220 57304 8248 57335
rect 9030 57332 9036 57384
rect 9088 57372 9094 57384
rect 9585 57375 9643 57381
rect 9585 57372 9597 57375
rect 9088 57344 9597 57372
rect 9088 57332 9094 57344
rect 9585 57341 9597 57344
rect 9631 57341 9643 57375
rect 9585 57335 9643 57341
rect 9766 57332 9772 57384
rect 9824 57372 9830 57384
rect 10229 57375 10287 57381
rect 10229 57372 10241 57375
rect 9824 57344 10241 57372
rect 9824 57332 9830 57344
rect 10229 57341 10241 57344
rect 10275 57341 10287 57375
rect 10229 57335 10287 57341
rect 11057 57375 11115 57381
rect 11057 57341 11069 57375
rect 11103 57372 11115 57375
rect 11422 57372 11428 57384
rect 11103 57344 11428 57372
rect 11103 57341 11115 57344
rect 11057 57335 11115 57341
rect 11422 57332 11428 57344
rect 11480 57332 11486 57384
rect 12250 57372 12256 57384
rect 12211 57344 12256 57372
rect 12250 57332 12256 57344
rect 12308 57332 12314 57384
rect 13464 57381 13492 57480
rect 26142 57468 26148 57480
rect 26200 57468 26206 57520
rect 26694 57468 26700 57520
rect 26752 57517 26758 57520
rect 26752 57511 26801 57517
rect 26752 57477 26755 57511
rect 26789 57477 26801 57511
rect 26878 57508 26884 57520
rect 26839 57480 26884 57508
rect 26752 57471 26801 57477
rect 26752 57468 26758 57471
rect 26878 57468 26884 57480
rect 26936 57468 26942 57520
rect 26988 57508 27016 57548
rect 27062 57536 27068 57588
rect 27120 57576 27126 57588
rect 29733 57579 29791 57585
rect 29733 57576 29745 57579
rect 27120 57548 29745 57576
rect 27120 57536 27126 57548
rect 29733 57545 29745 57548
rect 29779 57545 29791 57579
rect 29733 57539 29791 57545
rect 29914 57536 29920 57588
rect 29972 57576 29978 57588
rect 32125 57579 32183 57585
rect 32125 57576 32137 57579
rect 29972 57548 32137 57576
rect 29972 57536 29978 57548
rect 32125 57545 32137 57548
rect 32171 57545 32183 57579
rect 36265 57579 36323 57585
rect 36265 57576 36277 57579
rect 32125 57539 32183 57545
rect 32232 57548 36277 57576
rect 32232 57508 32260 57548
rect 36265 57545 36277 57548
rect 36311 57545 36323 57579
rect 36265 57539 36323 57545
rect 26988 57480 28479 57508
rect 14550 57400 14556 57452
rect 14608 57440 14614 57452
rect 14608 57412 15240 57440
rect 14608 57400 14614 57412
rect 12805 57375 12863 57381
rect 12805 57341 12817 57375
rect 12851 57341 12863 57375
rect 12805 57335 12863 57341
rect 13449 57375 13507 57381
rect 13449 57341 13461 57375
rect 13495 57341 13507 57375
rect 13449 57335 13507 57341
rect 7524 57276 8248 57304
rect 7524 57264 7530 57276
rect 11790 57264 11796 57316
rect 11848 57304 11854 57316
rect 12820 57304 12848 57335
rect 13814 57332 13820 57384
rect 13872 57372 13878 57384
rect 15105 57375 15163 57381
rect 15105 57372 15117 57375
rect 13872 57344 15117 57372
rect 13872 57332 13878 57344
rect 15105 57341 15117 57344
rect 15151 57341 15163 57375
rect 15212 57372 15240 57412
rect 15378 57400 15384 57452
rect 15436 57440 15442 57452
rect 15436 57412 16436 57440
rect 15436 57400 15442 57412
rect 16408 57381 16436 57412
rect 20070 57400 20076 57452
rect 20128 57440 20134 57452
rect 20128 57412 20760 57440
rect 20128 57400 20134 57412
rect 15749 57375 15807 57381
rect 15749 57372 15761 57375
rect 15212 57344 15761 57372
rect 15105 57335 15163 57341
rect 15749 57341 15761 57344
rect 15795 57341 15807 57375
rect 15749 57335 15807 57341
rect 16393 57375 16451 57381
rect 16393 57341 16405 57375
rect 16439 57341 16451 57375
rect 16393 57335 16451 57341
rect 16942 57332 16948 57384
rect 17000 57372 17006 57384
rect 17773 57375 17831 57381
rect 17773 57372 17785 57375
rect 17000 57344 17785 57372
rect 17000 57332 17006 57344
rect 17773 57341 17785 57344
rect 17819 57341 17831 57375
rect 17773 57335 17831 57341
rect 17954 57332 17960 57384
rect 18012 57372 18018 57384
rect 18417 57375 18475 57381
rect 18417 57372 18429 57375
rect 18012 57344 18429 57372
rect 18012 57332 18018 57344
rect 18417 57341 18429 57344
rect 18463 57341 18475 57375
rect 18417 57335 18475 57341
rect 18506 57332 18512 57384
rect 18564 57372 18570 57384
rect 19061 57375 19119 57381
rect 19061 57372 19073 57375
rect 18564 57344 19073 57372
rect 18564 57332 18570 57344
rect 19061 57341 19073 57344
rect 19107 57341 19119 57375
rect 19061 57335 19119 57341
rect 19334 57332 19340 57384
rect 19392 57372 19398 57384
rect 20441 57375 20499 57381
rect 20441 57372 20453 57375
rect 19392 57344 20453 57372
rect 19392 57332 19398 57344
rect 20441 57341 20453 57344
rect 20487 57341 20499 57375
rect 20732 57372 20760 57412
rect 20898 57400 20904 57452
rect 20956 57440 20962 57452
rect 20956 57412 21772 57440
rect 20956 57400 20962 57412
rect 21744 57381 21772 57412
rect 24210 57400 24216 57452
rect 24268 57440 24274 57452
rect 24489 57443 24547 57449
rect 24489 57440 24501 57443
rect 24268 57412 24501 57440
rect 24268 57400 24274 57412
rect 24489 57409 24501 57412
rect 24535 57409 24547 57443
rect 24489 57403 24547 57409
rect 26973 57443 27031 57449
rect 26973 57409 26985 57443
rect 27019 57440 27031 57443
rect 28350 57440 28356 57452
rect 27019 57412 28356 57440
rect 27019 57409 27031 57412
rect 26973 57403 27031 57409
rect 28350 57400 28356 57412
rect 28408 57400 28414 57452
rect 21085 57375 21143 57381
rect 21085 57372 21097 57375
rect 20732 57344 21097 57372
rect 20441 57335 20499 57341
rect 21085 57341 21097 57344
rect 21131 57341 21143 57375
rect 21085 57335 21143 57341
rect 21729 57375 21787 57381
rect 21729 57341 21741 57375
rect 21775 57341 21787 57375
rect 21729 57335 21787 57341
rect 22094 57332 22100 57384
rect 22152 57372 22158 57384
rect 23109 57375 23167 57381
rect 23109 57372 23121 57375
rect 22152 57344 23121 57372
rect 22152 57332 22158 57344
rect 23109 57341 23121 57344
rect 23155 57341 23167 57375
rect 24302 57372 24308 57384
rect 24263 57344 24308 57372
rect 23109 57335 23167 57341
rect 24302 57332 24308 57344
rect 24360 57332 24366 57384
rect 24578 57332 24584 57384
rect 24636 57372 24642 57384
rect 25958 57372 25964 57384
rect 24636 57344 24681 57372
rect 25919 57344 25964 57372
rect 24636 57332 24642 57344
rect 25958 57332 25964 57344
rect 26016 57332 26022 57384
rect 26145 57375 26203 57381
rect 26145 57341 26157 57375
rect 26191 57372 26203 57375
rect 26326 57372 26332 57384
rect 26191 57344 26332 57372
rect 26191 57341 26203 57344
rect 26145 57335 26203 57341
rect 26326 57332 26332 57344
rect 26384 57332 26390 57384
rect 28451 57381 28479 57480
rect 29112 57480 32260 57508
rect 29112 57381 29140 57480
rect 33410 57468 33416 57520
rect 33468 57508 33474 57520
rect 37553 57511 37611 57517
rect 37553 57508 37565 57511
rect 33468 57480 37565 57508
rect 33468 57468 33474 57480
rect 37553 57477 37565 57480
rect 37599 57477 37611 57511
rect 37553 57471 37611 57477
rect 46934 57468 46940 57520
rect 46992 57468 46998 57520
rect 53285 57511 53343 57517
rect 53285 57477 53297 57511
rect 53331 57508 53343 57511
rect 55122 57508 55128 57520
rect 53331 57480 55128 57508
rect 53331 57477 53343 57480
rect 53285 57471 53343 57477
rect 55122 57468 55128 57480
rect 55180 57468 55186 57520
rect 55585 57511 55643 57517
rect 55585 57477 55597 57511
rect 55631 57508 55643 57511
rect 55674 57508 55680 57520
rect 55631 57480 55680 57508
rect 55631 57477 55643 57480
rect 55585 57471 55643 57477
rect 55674 57468 55680 57480
rect 55732 57468 55738 57520
rect 29181 57443 29239 57449
rect 29181 57409 29193 57443
rect 29227 57440 29239 57443
rect 29638 57440 29644 57452
rect 29227 57412 29644 57440
rect 29227 57409 29239 57412
rect 29181 57403 29239 57409
rect 29638 57400 29644 57412
rect 29696 57400 29702 57452
rect 29822 57400 29828 57452
rect 29880 57440 29886 57452
rect 29880 57412 34468 57440
rect 29880 57400 29886 57412
rect 28437 57375 28495 57381
rect 28437 57341 28449 57375
rect 28483 57341 28495 57375
rect 28437 57335 28495 57341
rect 29089 57375 29147 57381
rect 29089 57341 29101 57375
rect 29135 57341 29147 57375
rect 29089 57335 29147 57341
rect 29270 57332 29276 57384
rect 29328 57372 29334 57384
rect 29917 57375 29975 57381
rect 29917 57372 29929 57375
rect 29328 57344 29929 57372
rect 29328 57332 29334 57344
rect 29917 57341 29929 57344
rect 29963 57341 29975 57375
rect 29917 57335 29975 57341
rect 31481 57375 31539 57381
rect 31481 57341 31493 57375
rect 31527 57372 31539 57375
rect 32122 57372 32128 57384
rect 31527 57344 32128 57372
rect 31527 57341 31539 57344
rect 31481 57335 31539 57341
rect 32122 57332 32128 57344
rect 32180 57332 32186 57384
rect 32306 57372 32312 57384
rect 32267 57344 32312 57372
rect 32306 57332 32312 57344
rect 32364 57332 32370 57384
rect 32674 57332 32680 57384
rect 32732 57372 32738 57384
rect 32732 57344 33732 57372
rect 32732 57332 32738 57344
rect 11848 57276 12848 57304
rect 11848 57264 11854 57276
rect 20162 57264 20168 57316
rect 20220 57304 20226 57316
rect 20220 57276 22094 57304
rect 20220 57264 20226 57276
rect 5534 57236 5540 57248
rect 5495 57208 5540 57236
rect 5534 57196 5540 57208
rect 5592 57196 5598 57248
rect 9769 57239 9827 57245
rect 9769 57205 9781 57239
rect 9815 57236 9827 57239
rect 11054 57236 11060 57248
rect 9815 57208 11060 57236
rect 9815 57205 9827 57208
rect 9769 57199 9827 57205
rect 11054 57196 11060 57208
rect 11112 57196 11118 57248
rect 11238 57236 11244 57248
rect 11199 57208 11244 57236
rect 11238 57196 11244 57208
rect 11296 57196 11302 57248
rect 12434 57236 12440 57248
rect 12395 57208 12440 57236
rect 12434 57196 12440 57208
rect 12492 57196 12498 57248
rect 13630 57236 13636 57248
rect 13591 57208 13636 57236
rect 13630 57196 13636 57208
rect 13688 57196 13694 57248
rect 14921 57239 14979 57245
rect 14921 57205 14933 57239
rect 14967 57236 14979 57239
rect 15102 57236 15108 57248
rect 14967 57208 15108 57236
rect 14967 57205 14979 57208
rect 14921 57199 14979 57205
rect 15102 57196 15108 57208
rect 15160 57196 15166 57248
rect 15562 57236 15568 57248
rect 15523 57208 15568 57236
rect 15562 57196 15568 57208
rect 15620 57196 15626 57248
rect 15654 57196 15660 57248
rect 15712 57236 15718 57248
rect 16209 57239 16267 57245
rect 16209 57236 16221 57239
rect 15712 57208 16221 57236
rect 15712 57196 15718 57208
rect 16209 57205 16221 57208
rect 16255 57205 16267 57239
rect 16209 57199 16267 57205
rect 17589 57239 17647 57245
rect 17589 57205 17601 57239
rect 17635 57236 17647 57239
rect 17954 57236 17960 57248
rect 17635 57208 17960 57236
rect 17635 57205 17647 57208
rect 17589 57199 17647 57205
rect 17954 57196 17960 57208
rect 18012 57196 18018 57248
rect 18230 57236 18236 57248
rect 18191 57208 18236 57236
rect 18230 57196 18236 57208
rect 18288 57196 18294 57248
rect 18874 57236 18880 57248
rect 18835 57208 18880 57236
rect 18874 57196 18880 57208
rect 18932 57196 18938 57248
rect 20254 57236 20260 57248
rect 20215 57208 20260 57236
rect 20254 57196 20260 57208
rect 20312 57196 20318 57248
rect 20346 57196 20352 57248
rect 20404 57236 20410 57248
rect 20901 57239 20959 57245
rect 20901 57236 20913 57239
rect 20404 57208 20913 57236
rect 20404 57196 20410 57208
rect 20901 57205 20913 57208
rect 20947 57205 20959 57239
rect 21542 57236 21548 57248
rect 21503 57208 21548 57236
rect 20901 57199 20959 57205
rect 21542 57196 21548 57208
rect 21600 57196 21606 57248
rect 22066 57236 22094 57276
rect 23014 57264 23020 57316
rect 23072 57304 23078 57316
rect 26605 57307 26663 57313
rect 26605 57304 26617 57307
rect 23072 57276 26617 57304
rect 23072 57264 23078 57276
rect 26605 57273 26617 57276
rect 26651 57273 26663 57307
rect 26605 57267 26663 57273
rect 26694 57264 26700 57316
rect 26752 57304 26758 57316
rect 28994 57304 29000 57316
rect 26752 57276 29000 57304
rect 26752 57264 26758 57276
rect 28994 57264 29000 57276
rect 29052 57264 29058 57316
rect 29178 57264 29184 57316
rect 29236 57304 29242 57316
rect 33704 57304 33732 57344
rect 33778 57332 33784 57384
rect 33836 57372 33842 57384
rect 34440 57381 34468 57412
rect 36630 57400 36636 57452
rect 36688 57440 36694 57452
rect 36688 57412 38700 57440
rect 36688 57400 36694 57412
rect 34425 57375 34483 57381
rect 33836 57344 33881 57372
rect 33836 57332 33842 57344
rect 34425 57341 34437 57375
rect 34471 57341 34483 57375
rect 34425 57335 34483 57341
rect 35069 57375 35127 57381
rect 35069 57341 35081 57375
rect 35115 57372 35127 57375
rect 35250 57372 35256 57384
rect 35115 57344 35256 57372
rect 35115 57341 35127 57344
rect 35069 57335 35127 57341
rect 35250 57332 35256 57344
rect 35308 57332 35314 57384
rect 36446 57372 36452 57384
rect 36407 57344 36452 57372
rect 36446 57332 36452 57344
rect 36504 57332 36510 57384
rect 37090 57372 37096 57384
rect 37051 57344 37096 57372
rect 37090 57332 37096 57344
rect 37148 57332 37154 57384
rect 37737 57375 37795 57381
rect 37737 57341 37749 57375
rect 37783 57341 37795 57375
rect 38672 57372 38700 57412
rect 39022 57400 39028 57452
rect 39080 57440 39086 57452
rect 39080 57412 40264 57440
rect 39080 57400 39086 57412
rect 40236 57381 40264 57412
rect 41414 57400 41420 57452
rect 41472 57440 41478 57452
rect 41472 57412 42288 57440
rect 41472 57400 41478 57412
rect 39117 57375 39175 57381
rect 39117 57372 39129 57375
rect 38672 57344 39129 57372
rect 37737 57335 37795 57341
rect 39117 57341 39129 57344
rect 39163 57341 39175 57375
rect 39117 57335 39175 57341
rect 39761 57375 39819 57381
rect 39761 57341 39773 57375
rect 39807 57341 39819 57375
rect 39761 57335 39819 57341
rect 40221 57375 40279 57381
rect 40221 57341 40233 57375
rect 40267 57341 40279 57375
rect 40221 57335 40279 57341
rect 37752 57304 37780 57335
rect 29236 57276 33640 57304
rect 33704 57276 37780 57304
rect 29236 57264 29242 57276
rect 22925 57239 22983 57245
rect 22925 57236 22937 57239
rect 22066 57208 22937 57236
rect 22925 57205 22937 57208
rect 22971 57205 22983 57239
rect 24118 57236 24124 57248
rect 24079 57208 24124 57236
rect 22925 57199 22983 57205
rect 24118 57196 24124 57208
rect 24176 57196 24182 57248
rect 25866 57196 25872 57248
rect 25924 57236 25930 57248
rect 26053 57239 26111 57245
rect 26053 57236 26065 57239
rect 25924 57208 26065 57236
rect 25924 57196 25930 57208
rect 26053 57205 26065 57208
rect 26099 57205 26111 57239
rect 26053 57199 26111 57205
rect 26142 57196 26148 57248
rect 26200 57236 26206 57248
rect 27249 57239 27307 57245
rect 27249 57236 27261 57239
rect 26200 57208 27261 57236
rect 26200 57196 26206 57208
rect 27249 57205 27261 57208
rect 27295 57205 27307 57239
rect 28258 57236 28264 57248
rect 28219 57208 28264 57236
rect 27249 57199 27307 57205
rect 28258 57196 28264 57208
rect 28316 57196 28322 57248
rect 31573 57239 31631 57245
rect 31573 57205 31585 57239
rect 31619 57236 31631 57239
rect 31662 57236 31668 57248
rect 31619 57208 31668 57236
rect 31619 57205 31631 57208
rect 31573 57199 31631 57205
rect 31662 57196 31668 57208
rect 31720 57196 31726 57248
rect 33612 57245 33640 57276
rect 38194 57264 38200 57316
rect 38252 57304 38258 57316
rect 39776 57304 39804 57335
rect 40586 57332 40592 57384
rect 40644 57372 40650 57384
rect 42260 57381 42288 57412
rect 45370 57400 45376 57452
rect 45428 57440 45434 57452
rect 46952 57440 46980 57468
rect 45428 57412 45600 57440
rect 46952 57412 47624 57440
rect 45428 57400 45434 57412
rect 41601 57375 41659 57381
rect 41601 57372 41613 57375
rect 40644 57344 41613 57372
rect 40644 57332 40650 57344
rect 41601 57341 41613 57344
rect 41647 57341 41659 57375
rect 41601 57335 41659 57341
rect 42245 57375 42303 57381
rect 42245 57341 42257 57375
rect 42291 57341 42303 57375
rect 42978 57372 42984 57384
rect 42939 57344 42984 57372
rect 42245 57335 42303 57341
rect 42978 57332 42984 57344
rect 43036 57332 43042 57384
rect 43714 57332 43720 57384
rect 43772 57372 43778 57384
rect 44269 57375 44327 57381
rect 44269 57372 44281 57375
rect 43772 57344 44281 57372
rect 43772 57332 43778 57344
rect 44269 57341 44281 57344
rect 44315 57341 44327 57375
rect 44269 57335 44327 57341
rect 44542 57332 44548 57384
rect 44600 57372 44606 57384
rect 45572 57381 45600 57412
rect 44913 57375 44971 57381
rect 44913 57372 44925 57375
rect 44600 57344 44925 57372
rect 44600 57332 44606 57344
rect 44913 57341 44925 57344
rect 44959 57341 44971 57375
rect 44913 57335 44971 57341
rect 45557 57375 45615 57381
rect 45557 57341 45569 57375
rect 45603 57341 45615 57375
rect 45557 57335 45615 57341
rect 46106 57332 46112 57384
rect 46164 57372 46170 57384
rect 47596 57381 47624 57412
rect 49234 57400 49240 57452
rect 49292 57440 49298 57452
rect 49292 57412 49832 57440
rect 49292 57400 49298 57412
rect 46937 57375 46995 57381
rect 46937 57372 46949 57375
rect 46164 57344 46949 57372
rect 46164 57332 46170 57344
rect 46937 57341 46949 57344
rect 46983 57341 46995 57375
rect 46937 57335 46995 57341
rect 47581 57375 47639 57381
rect 47581 57341 47593 57375
rect 47627 57341 47639 57375
rect 47581 57335 47639 57341
rect 47670 57332 47676 57384
rect 47728 57372 47734 57384
rect 48225 57375 48283 57381
rect 48225 57372 48237 57375
rect 47728 57344 48237 57372
rect 47728 57332 47734 57344
rect 48225 57341 48237 57344
rect 48271 57341 48283 57375
rect 48225 57335 48283 57341
rect 48498 57332 48504 57384
rect 48556 57372 48562 57384
rect 49605 57375 49663 57381
rect 49605 57372 49617 57375
rect 48556 57344 49617 57372
rect 48556 57332 48562 57344
rect 49605 57341 49617 57344
rect 49651 57341 49663 57375
rect 49804 57372 49832 57412
rect 50062 57400 50068 57452
rect 50120 57440 50126 57452
rect 54021 57443 54079 57449
rect 50120 57412 50936 57440
rect 50120 57400 50126 57412
rect 50908 57381 50936 57412
rect 54021 57409 54033 57443
rect 54067 57440 54079 57443
rect 56410 57440 56416 57452
rect 54067 57412 56416 57440
rect 54067 57409 54079 57412
rect 54021 57403 54079 57409
rect 56410 57400 56416 57412
rect 56468 57400 56474 57452
rect 58158 57440 58164 57452
rect 58119 57412 58164 57440
rect 58158 57400 58164 57412
rect 58216 57400 58222 57452
rect 50249 57375 50307 57381
rect 50249 57372 50261 57375
rect 49804 57344 50261 57372
rect 49605 57335 49663 57341
rect 50249 57341 50261 57344
rect 50295 57341 50307 57375
rect 50249 57335 50307 57341
rect 50893 57375 50951 57381
rect 50893 57341 50905 57375
rect 50939 57341 50951 57375
rect 50893 57335 50951 57341
rect 52365 57375 52423 57381
rect 52365 57341 52377 57375
rect 52411 57372 52423 57375
rect 53742 57372 53748 57384
rect 52411 57344 53748 57372
rect 52411 57341 52423 57344
rect 52365 57335 52423 57341
rect 53742 57332 53748 57344
rect 53800 57332 53806 57384
rect 54110 57332 54116 57384
rect 54168 57372 54174 57384
rect 56045 57375 56103 57381
rect 56045 57372 56057 57375
rect 54168 57344 56057 57372
rect 54168 57332 54174 57344
rect 56045 57341 56057 57344
rect 56091 57341 56103 57375
rect 56045 57335 56103 57341
rect 56229 57375 56287 57381
rect 56229 57341 56241 57375
rect 56275 57372 56287 57375
rect 56778 57372 56784 57384
rect 56275 57344 56784 57372
rect 56275 57341 56287 57344
rect 56229 57335 56287 57341
rect 56778 57332 56784 57344
rect 56836 57332 56842 57384
rect 53098 57304 53104 57316
rect 38252 57276 39804 57304
rect 53059 57276 53104 57304
rect 38252 57264 38258 57276
rect 53098 57264 53104 57276
rect 53156 57264 53162 57316
rect 53837 57307 53895 57313
rect 53837 57273 53849 57307
rect 53883 57304 53895 57307
rect 55401 57307 55459 57313
rect 53883 57276 55214 57304
rect 53883 57273 53895 57276
rect 53837 57267 53895 57273
rect 33597 57239 33655 57245
rect 33597 57205 33609 57239
rect 33643 57205 33655 57239
rect 34238 57236 34244 57248
rect 34199 57208 34244 57236
rect 33597 57199 33655 57205
rect 34238 57196 34244 57208
rect 34296 57196 34302 57248
rect 34606 57196 34612 57248
rect 34664 57236 34670 57248
rect 35253 57239 35311 57245
rect 35253 57236 35265 57239
rect 34664 57208 35265 57236
rect 34664 57196 34670 57208
rect 35253 57205 35265 57208
rect 35299 57205 35311 57239
rect 36906 57236 36912 57248
rect 36867 57208 36912 57236
rect 35253 57199 35311 57205
rect 36906 57196 36912 57208
rect 36964 57196 36970 57248
rect 38930 57236 38936 57248
rect 38891 57208 38936 57236
rect 38930 57196 38936 57208
rect 38988 57196 38994 57248
rect 39574 57236 39580 57248
rect 39535 57208 39580 57236
rect 39574 57196 39580 57208
rect 39632 57196 39638 57248
rect 40402 57236 40408 57248
rect 40363 57208 40408 57236
rect 40402 57196 40408 57208
rect 40460 57196 40466 57248
rect 55186 57236 55214 57276
rect 55401 57273 55413 57307
rect 55447 57304 55459 57307
rect 56689 57307 56747 57313
rect 56689 57304 56701 57307
rect 55447 57276 56701 57304
rect 55447 57273 55459 57276
rect 55401 57267 55459 57273
rect 56689 57273 56701 57276
rect 56735 57273 56747 57307
rect 57974 57304 57980 57316
rect 57935 57276 57980 57304
rect 56689 57267 56747 57273
rect 57974 57264 57980 57276
rect 58032 57264 58038 57316
rect 58342 57236 58348 57248
rect 55186 57208 58348 57236
rect 58342 57196 58348 57208
rect 58400 57196 58406 57248
rect 1104 57146 58880 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 50326 57146
rect 50378 57094 50390 57146
rect 50442 57094 50454 57146
rect 50506 57094 50518 57146
rect 50570 57094 58880 57146
rect 1104 57072 58880 57094
rect 4246 56992 4252 57044
rect 4304 57032 4310 57044
rect 4893 57035 4951 57041
rect 4893 57032 4905 57035
rect 4304 57004 4905 57032
rect 4304 56992 4310 57004
rect 4893 57001 4905 57004
rect 4939 57001 4951 57035
rect 4893 56995 4951 57001
rect 10597 57035 10655 57041
rect 10597 57001 10609 57035
rect 10643 57001 10655 57035
rect 10597 56995 10655 57001
rect 16117 57035 16175 57041
rect 16117 57001 16129 57035
rect 16163 57032 16175 57035
rect 23661 57035 23719 57041
rect 23661 57032 23673 57035
rect 16163 57004 16574 57032
rect 16163 57001 16175 57004
rect 16117 56995 16175 57001
rect 4525 56967 4583 56973
rect 4525 56964 4537 56967
rect 3160 56936 4537 56964
rect 3160 56908 3188 56936
rect 4525 56933 4537 56936
rect 4571 56933 4583 56967
rect 4525 56927 4583 56933
rect 4617 56967 4675 56973
rect 4617 56933 4629 56967
rect 4663 56964 4675 56967
rect 8294 56964 8300 56976
rect 4663 56936 8300 56964
rect 4663 56933 4675 56936
rect 4617 56927 4675 56933
rect 8294 56924 8300 56936
rect 8352 56924 8358 56976
rect 10612 56964 10640 56995
rect 12250 56964 12256 56976
rect 10612 56936 12256 56964
rect 1394 56896 1400 56908
rect 1355 56868 1400 56896
rect 1394 56856 1400 56868
rect 1452 56856 1458 56908
rect 2130 56896 2136 56908
rect 2091 56868 2136 56896
rect 2130 56856 2136 56868
rect 2188 56856 2194 56908
rect 3142 56896 3148 56908
rect 3103 56868 3148 56896
rect 3142 56856 3148 56868
rect 3200 56856 3206 56908
rect 3326 56856 3332 56908
rect 3384 56896 3390 56908
rect 4734 56899 4792 56905
rect 4734 56896 4746 56899
rect 3384 56868 4746 56896
rect 3384 56856 3390 56868
rect 4734 56865 4746 56868
rect 4780 56865 4792 56899
rect 8202 56896 8208 56908
rect 8163 56868 8208 56896
rect 4734 56859 4792 56865
rect 8202 56856 8208 56868
rect 8260 56856 8266 56908
rect 10594 56856 10600 56908
rect 10652 56896 10658 56908
rect 11716 56905 11744 56936
rect 12250 56924 12256 56936
rect 12308 56924 12314 56976
rect 12986 56924 12992 56976
rect 13044 56964 13050 56976
rect 13081 56967 13139 56973
rect 13081 56964 13093 56967
rect 13044 56936 13093 56964
rect 13044 56924 13050 56936
rect 13081 56933 13093 56936
rect 13127 56933 13139 56967
rect 13081 56927 13139 56933
rect 14737 56967 14795 56973
rect 14737 56933 14749 56967
rect 14783 56964 14795 56967
rect 15562 56964 15568 56976
rect 14783 56936 15568 56964
rect 14783 56933 14795 56936
rect 14737 56927 14795 56933
rect 15562 56924 15568 56936
rect 15620 56924 15626 56976
rect 10781 56899 10839 56905
rect 10781 56896 10793 56899
rect 10652 56868 10793 56896
rect 10652 56856 10658 56868
rect 10781 56865 10793 56868
rect 10827 56865 10839 56899
rect 10781 56859 10839 56865
rect 11701 56899 11759 56905
rect 11701 56865 11713 56899
rect 11747 56865 11759 56899
rect 11974 56896 11980 56908
rect 11935 56868 11980 56896
rect 11701 56859 11759 56865
rect 11974 56856 11980 56868
rect 12032 56856 12038 56908
rect 14884 56899 14942 56905
rect 14884 56865 14896 56899
rect 14930 56896 14942 56899
rect 15654 56896 15660 56908
rect 14930 56868 15660 56896
rect 14930 56865 14942 56868
rect 14884 56859 14942 56865
rect 15654 56856 15660 56868
rect 15712 56856 15718 56908
rect 16114 56856 16120 56908
rect 16172 56896 16178 56908
rect 16301 56899 16359 56905
rect 16301 56896 16313 56899
rect 16172 56868 16313 56896
rect 16172 56856 16178 56868
rect 16301 56865 16313 56868
rect 16347 56865 16359 56899
rect 16301 56859 16359 56865
rect 4249 56831 4307 56837
rect 4249 56797 4261 56831
rect 4295 56828 4307 56831
rect 4614 56828 4620 56840
rect 4295 56800 4620 56828
rect 4295 56797 4307 56800
rect 4249 56791 4307 56797
rect 4614 56788 4620 56800
rect 4672 56788 4678 56840
rect 11054 56788 11060 56840
rect 11112 56828 11118 56840
rect 11790 56828 11796 56840
rect 11112 56800 11796 56828
rect 11112 56788 11118 56800
rect 11790 56788 11796 56800
rect 11848 56788 11854 56840
rect 12158 56828 12164 56840
rect 12119 56800 12164 56828
rect 12158 56788 12164 56800
rect 12216 56788 12222 56840
rect 15102 56828 15108 56840
rect 15063 56800 15108 56828
rect 15102 56788 15108 56800
rect 15160 56788 15166 56840
rect 13170 56720 13176 56772
rect 13228 56760 13234 56772
rect 13265 56763 13323 56769
rect 13265 56760 13277 56763
rect 13228 56732 13277 56760
rect 13228 56720 13234 56732
rect 13265 56729 13277 56732
rect 13311 56760 13323 56763
rect 15013 56763 15071 56769
rect 15013 56760 15025 56763
rect 13311 56732 15025 56760
rect 13311 56729 13323 56732
rect 13265 56723 13323 56729
rect 15013 56729 15025 56732
rect 15059 56729 15071 56763
rect 15013 56723 15071 56729
rect 15381 56763 15439 56769
rect 15381 56729 15393 56763
rect 15427 56760 15439 56763
rect 16546 56760 16574 57004
rect 22066 57004 23673 57032
rect 17589 56967 17647 56973
rect 17589 56933 17601 56967
rect 17635 56964 17647 56967
rect 18230 56964 18236 56976
rect 17635 56936 18236 56964
rect 17635 56933 17647 56936
rect 17589 56927 17647 56933
rect 18230 56924 18236 56936
rect 18288 56924 18294 56976
rect 19981 56967 20039 56973
rect 19981 56933 19993 56967
rect 20027 56964 20039 56967
rect 21542 56964 21548 56976
rect 20027 56936 21548 56964
rect 20027 56933 20039 56936
rect 19981 56927 20039 56933
rect 21542 56924 21548 56936
rect 21600 56924 21606 56976
rect 17736 56899 17794 56905
rect 17736 56865 17748 56899
rect 17782 56896 17794 56899
rect 18874 56896 18880 56908
rect 17782 56868 18880 56896
rect 17782 56865 17794 56868
rect 17736 56859 17794 56865
rect 18874 56856 18880 56868
rect 18932 56856 18938 56908
rect 20717 56899 20775 56905
rect 19812 56868 20484 56896
rect 17954 56828 17960 56840
rect 17915 56800 17960 56828
rect 17954 56788 17960 56800
rect 18012 56788 18018 56840
rect 18325 56831 18383 56837
rect 18325 56797 18337 56831
rect 18371 56828 18383 56831
rect 19812 56828 19840 56868
rect 20162 56837 20168 56840
rect 18371 56800 19840 56828
rect 20128 56831 20168 56837
rect 18371 56797 18383 56800
rect 18325 56791 18383 56797
rect 20128 56797 20140 56831
rect 20128 56791 20168 56797
rect 20162 56788 20168 56791
rect 20220 56788 20226 56840
rect 20346 56828 20352 56840
rect 20307 56800 20352 56828
rect 20346 56788 20352 56800
rect 20404 56788 20410 56840
rect 20456 56828 20484 56868
rect 20717 56865 20729 56899
rect 20763 56896 20775 56899
rect 21177 56899 21235 56905
rect 21177 56896 21189 56899
rect 20763 56868 21189 56896
rect 20763 56865 20775 56868
rect 20717 56859 20775 56865
rect 21177 56865 21189 56868
rect 21223 56865 21235 56899
rect 21177 56859 21235 56865
rect 21324 56899 21382 56905
rect 21324 56865 21336 56899
rect 21370 56896 21382 56899
rect 22066 56896 22094 57004
rect 23661 57001 23673 57004
rect 23707 57001 23719 57035
rect 23661 56995 23719 57001
rect 26878 56992 26884 57044
rect 26936 57032 26942 57044
rect 27341 57035 27399 57041
rect 27341 57032 27353 57035
rect 26936 57004 27353 57032
rect 26936 56992 26942 57004
rect 27341 57001 27353 57004
rect 27387 57001 27399 57035
rect 35713 57035 35771 57041
rect 35713 57032 35725 57035
rect 27341 56995 27399 57001
rect 28644 57004 35725 57032
rect 23017 56967 23075 56973
rect 23017 56933 23029 56967
rect 23063 56964 23075 56967
rect 28258 56964 28264 56976
rect 23063 56936 28264 56964
rect 23063 56933 23075 56936
rect 23017 56927 23075 56933
rect 28258 56924 28264 56936
rect 28316 56924 28322 56976
rect 21370 56868 22094 56896
rect 21370 56865 21382 56868
rect 21324 56859 21382 56865
rect 22462 56856 22468 56908
rect 22520 56896 22526 56908
rect 22557 56899 22615 56905
rect 22557 56896 22569 56899
rect 22520 56868 22569 56896
rect 22520 56856 22526 56868
rect 22557 56865 22569 56868
rect 22603 56865 22615 56899
rect 22557 56859 22615 56865
rect 25777 56899 25835 56905
rect 25777 56865 25789 56899
rect 25823 56896 25835 56899
rect 25866 56896 25872 56908
rect 25823 56868 25872 56896
rect 25823 56865 25835 56868
rect 25777 56859 25835 56865
rect 25866 56856 25872 56868
rect 25924 56856 25930 56908
rect 26694 56896 26700 56908
rect 26655 56868 26700 56896
rect 26694 56856 26700 56868
rect 26752 56856 26758 56908
rect 26844 56899 26902 56905
rect 26844 56865 26856 56899
rect 26890 56896 26902 56899
rect 27246 56896 27252 56908
rect 26890 56868 27252 56896
rect 26890 56865 26902 56868
rect 26844 56859 26902 56865
rect 27246 56856 27252 56868
rect 27304 56856 27310 56908
rect 27982 56896 27988 56908
rect 27943 56868 27988 56896
rect 27982 56856 27988 56868
rect 28040 56856 28046 56908
rect 28644 56905 28672 57004
rect 35713 57001 35725 57004
rect 35759 57001 35771 57035
rect 35713 56995 35771 57001
rect 35894 56992 35900 57044
rect 35952 57032 35958 57044
rect 35952 57004 37044 57032
rect 35952 56992 35958 57004
rect 29178 56924 29184 56976
rect 29236 56964 29242 56976
rect 36906 56964 36912 56976
rect 29236 56936 36912 56964
rect 29236 56924 29242 56936
rect 36906 56924 36912 56936
rect 36964 56924 36970 56976
rect 28629 56899 28687 56905
rect 28629 56865 28641 56899
rect 28675 56865 28687 56899
rect 29914 56896 29920 56908
rect 28629 56859 28687 56865
rect 29012 56868 29920 56896
rect 21545 56831 21603 56837
rect 21545 56828 21557 56831
rect 20456 56800 21557 56828
rect 21545 56797 21557 56800
rect 21591 56797 21603 56831
rect 21545 56791 21603 56797
rect 21913 56831 21971 56837
rect 21913 56797 21925 56831
rect 21959 56828 21971 56831
rect 23014 56828 23020 56840
rect 21959 56800 23020 56828
rect 21959 56797 21971 56800
rect 21913 56791 21971 56797
rect 23014 56788 23020 56800
rect 23072 56788 23078 56840
rect 23382 56828 23388 56840
rect 23343 56800 23388 56828
rect 23382 56788 23388 56800
rect 23440 56788 23446 56840
rect 26053 56831 26111 56837
rect 26053 56797 26065 56831
rect 26099 56828 26111 56831
rect 26326 56828 26332 56840
rect 26099 56800 26332 56828
rect 26099 56797 26111 56800
rect 26053 56791 26111 56797
rect 26326 56788 26332 56800
rect 26384 56788 26390 56840
rect 27065 56831 27123 56837
rect 27065 56797 27077 56831
rect 27111 56828 27123 56831
rect 29012 56828 29040 56868
rect 29914 56856 29920 56868
rect 29972 56856 29978 56908
rect 31294 56905 31300 56908
rect 31288 56859 31300 56905
rect 31352 56896 31358 56908
rect 33588 56899 33646 56905
rect 31352 56868 31388 56896
rect 31294 56856 31300 56859
rect 31352 56856 31358 56868
rect 33588 56865 33600 56899
rect 33634 56896 33646 56899
rect 35434 56896 35440 56908
rect 33634 56868 35440 56896
rect 33634 56865 33646 56868
rect 33588 56859 33646 56865
rect 35434 56856 35440 56868
rect 35492 56856 35498 56908
rect 35894 56896 35900 56908
rect 35855 56868 35900 56896
rect 35894 56856 35900 56868
rect 35952 56856 35958 56908
rect 36541 56899 36599 56905
rect 36541 56865 36553 56899
rect 36587 56865 36599 56899
rect 37016 56896 37044 57004
rect 53098 56992 53104 57044
rect 53156 57032 53162 57044
rect 55217 57035 55275 57041
rect 55217 57032 55229 57035
rect 53156 57004 55229 57032
rect 53156 56992 53162 57004
rect 55217 57001 55229 57004
rect 55263 57001 55275 57035
rect 55217 56995 55275 57001
rect 57974 56992 57980 57044
rect 58032 57032 58038 57044
rect 58161 57035 58219 57041
rect 58161 57032 58173 57035
rect 58032 57004 58173 57032
rect 58032 56992 58038 57004
rect 58161 57001 58173 57004
rect 58207 57001 58219 57035
rect 58161 56995 58219 57001
rect 57054 56964 57060 56976
rect 57015 56936 57060 56964
rect 57054 56924 57060 56936
rect 57112 56924 57118 56976
rect 37185 56899 37243 56905
rect 37185 56896 37197 56899
rect 37016 56868 37197 56896
rect 36541 56859 36599 56865
rect 37185 56865 37197 56868
rect 37231 56865 37243 56899
rect 37185 56859 37243 56865
rect 29178 56828 29184 56840
rect 27111 56800 29040 56828
rect 29139 56800 29184 56828
rect 27111 56797 27123 56800
rect 27065 56791 27123 56797
rect 29178 56788 29184 56800
rect 29236 56788 29242 56840
rect 29270 56788 29276 56840
rect 29328 56828 29334 56840
rect 29328 56800 29373 56828
rect 29328 56788 29334 56800
rect 30742 56788 30748 56840
rect 30800 56828 30806 56840
rect 31021 56831 31079 56837
rect 31021 56828 31033 56831
rect 30800 56800 31033 56828
rect 30800 56788 30806 56800
rect 31021 56797 31033 56800
rect 31067 56797 31079 56831
rect 33318 56828 33324 56840
rect 33279 56800 33324 56828
rect 31021 56791 31079 56797
rect 33318 56788 33324 56800
rect 33376 56788 33382 56840
rect 34422 56788 34428 56840
rect 34480 56828 34486 56840
rect 36556 56828 36584 56859
rect 37458 56856 37464 56908
rect 37516 56896 37522 56908
rect 37829 56899 37887 56905
rect 37829 56896 37841 56899
rect 37516 56868 37841 56896
rect 37516 56856 37522 56868
rect 37829 56865 37841 56868
rect 37875 56865 37887 56899
rect 39758 56896 39764 56908
rect 39719 56868 39764 56896
rect 37829 56859 37887 56865
rect 39758 56856 39764 56868
rect 39816 56856 39822 56908
rect 42150 56896 42156 56908
rect 42111 56868 42156 56896
rect 42150 56856 42156 56868
rect 42208 56856 42214 56908
rect 51074 56856 51080 56908
rect 51132 56896 51138 56908
rect 51445 56899 51503 56905
rect 51445 56896 51457 56899
rect 51132 56868 51457 56896
rect 51132 56856 51138 56868
rect 51445 56865 51457 56868
rect 51491 56865 51503 56899
rect 51445 56859 51503 56865
rect 51626 56856 51632 56908
rect 51684 56896 51690 56908
rect 52089 56899 52147 56905
rect 52089 56896 52101 56899
rect 51684 56868 52101 56896
rect 51684 56856 51690 56868
rect 52089 56865 52101 56868
rect 52135 56865 52147 56899
rect 54110 56896 54116 56908
rect 54071 56868 54116 56896
rect 52089 56859 52147 56865
rect 54110 56856 54116 56868
rect 54168 56856 54174 56908
rect 56873 56899 56931 56905
rect 56873 56865 56885 56899
rect 56919 56896 56931 56899
rect 57146 56896 57152 56908
rect 56919 56868 57152 56896
rect 56919 56865 56931 56868
rect 56873 56859 56931 56865
rect 57146 56856 57152 56868
rect 57204 56856 57210 56908
rect 54570 56828 54576 56840
rect 34480 56800 36584 56828
rect 54531 56800 54576 56828
rect 34480 56788 34486 56800
rect 54570 56788 54576 56800
rect 54628 56788 54634 56840
rect 54754 56828 54760 56840
rect 54715 56800 54760 56828
rect 54754 56788 54760 56800
rect 54812 56788 54818 56840
rect 56594 56788 56600 56840
rect 56652 56828 56658 56840
rect 57517 56831 57575 56837
rect 57517 56828 57529 56831
rect 56652 56800 57529 56828
rect 56652 56788 56658 56800
rect 57517 56797 57529 56800
rect 57563 56797 57575 56831
rect 57517 56791 57575 56797
rect 57701 56831 57759 56837
rect 57701 56797 57713 56831
rect 57747 56797 57759 56831
rect 57701 56791 57759 56797
rect 17865 56763 17923 56769
rect 17865 56760 17877 56763
rect 15427 56732 16252 56760
rect 16546 56732 17877 56760
rect 15427 56729 15439 56732
rect 15381 56723 15439 56729
rect 3234 56692 3240 56704
rect 3195 56664 3240 56692
rect 3234 56652 3240 56664
rect 3292 56652 3298 56704
rect 16224 56692 16252 56732
rect 17865 56729 17877 56732
rect 17911 56729 17923 56763
rect 20254 56760 20260 56772
rect 20215 56732 20260 56760
rect 17865 56723 17923 56729
rect 20254 56720 20260 56732
rect 20312 56720 20318 56772
rect 22373 56763 22431 56769
rect 22373 56729 22385 56763
rect 22419 56760 22431 56763
rect 23293 56763 23351 56769
rect 23293 56760 23305 56763
rect 22419 56732 23305 56760
rect 22419 56729 22431 56732
rect 22373 56723 22431 56729
rect 23293 56729 23305 56732
rect 23339 56729 23351 56763
rect 29086 56760 29092 56772
rect 29047 56732 29092 56760
rect 23293 56723 23351 56729
rect 29086 56720 29092 56732
rect 29144 56720 29150 56772
rect 29196 56732 30420 56760
rect 21453 56695 21511 56701
rect 21453 56692 21465 56695
rect 16224 56664 21465 56692
rect 21453 56661 21465 56664
rect 21499 56661 21511 56695
rect 21453 56655 21511 56661
rect 23106 56652 23112 56704
rect 23164 56701 23170 56704
rect 23164 56695 23213 56701
rect 23164 56661 23167 56695
rect 23201 56661 23213 56695
rect 25590 56692 25596 56704
rect 25551 56664 25596 56692
rect 23164 56655 23213 56661
rect 23164 56652 23170 56655
rect 25590 56652 25596 56664
rect 25648 56652 25654 56704
rect 25958 56692 25964 56704
rect 25919 56664 25964 56692
rect 25958 56652 25964 56664
rect 26016 56652 26022 56704
rect 26973 56695 27031 56701
rect 26973 56661 26985 56695
rect 27019 56692 27031 56695
rect 27062 56692 27068 56704
rect 27019 56664 27068 56692
rect 27019 56661 27031 56664
rect 26973 56655 27031 56661
rect 27062 56652 27068 56664
rect 27120 56652 27126 56704
rect 28077 56695 28135 56701
rect 28077 56661 28089 56695
rect 28123 56692 28135 56695
rect 28902 56692 28908 56704
rect 28123 56664 28908 56692
rect 28123 56661 28135 56664
rect 28077 56655 28135 56661
rect 28902 56652 28908 56664
rect 28960 56652 28966 56704
rect 28997 56695 29055 56701
rect 28997 56661 29009 56695
rect 29043 56692 29055 56695
rect 29196 56692 29224 56732
rect 29043 56664 29224 56692
rect 29043 56661 29055 56664
rect 28997 56655 29055 56661
rect 29270 56652 29276 56704
rect 29328 56692 29334 56704
rect 30282 56692 30288 56704
rect 29328 56664 30288 56692
rect 29328 56652 29334 56664
rect 30282 56652 30288 56664
rect 30340 56652 30346 56704
rect 30392 56692 30420 56732
rect 32122 56720 32128 56772
rect 32180 56760 32186 56772
rect 32401 56763 32459 56769
rect 32401 56760 32413 56763
rect 32180 56732 32413 56760
rect 32180 56720 32186 56732
rect 32401 56729 32413 56732
rect 32447 56729 32459 56763
rect 32401 56723 32459 56729
rect 34330 56720 34336 56772
rect 34388 56760 34394 56772
rect 37001 56763 37059 56769
rect 37001 56760 37013 56763
rect 34388 56732 37013 56760
rect 34388 56720 34394 56732
rect 37001 56729 37013 56732
rect 37047 56729 37059 56763
rect 37001 56723 37059 56729
rect 53469 56763 53527 56769
rect 53469 56729 53481 56763
rect 53515 56760 53527 56763
rect 55766 56760 55772 56772
rect 53515 56732 55772 56760
rect 53515 56729 53527 56732
rect 53469 56723 53527 56729
rect 55766 56720 55772 56732
rect 55824 56720 55830 56772
rect 56410 56720 56416 56772
rect 56468 56760 56474 56772
rect 57716 56760 57744 56791
rect 56468 56732 57744 56760
rect 56468 56720 56474 56732
rect 32950 56692 32956 56704
rect 30392 56664 32956 56692
rect 32950 56652 32956 56664
rect 33008 56652 33014 56704
rect 33134 56652 33140 56704
rect 33192 56692 33198 56704
rect 34422 56692 34428 56704
rect 33192 56664 34428 56692
rect 33192 56652 33198 56664
rect 34422 56652 34428 56664
rect 34480 56652 34486 56704
rect 34701 56695 34759 56701
rect 34701 56661 34713 56695
rect 34747 56692 34759 56695
rect 34790 56692 34796 56704
rect 34747 56664 34796 56692
rect 34747 56661 34759 56664
rect 34701 56655 34759 56661
rect 34790 56652 34796 56664
rect 34848 56652 34854 56704
rect 35250 56652 35256 56704
rect 35308 56692 35314 56704
rect 36357 56695 36415 56701
rect 36357 56692 36369 56695
rect 35308 56664 36369 56692
rect 35308 56652 35314 56664
rect 36357 56661 36369 56664
rect 36403 56661 36415 56695
rect 37642 56692 37648 56704
rect 37603 56664 37648 56692
rect 36357 56655 36415 56661
rect 37642 56652 37648 56664
rect 37700 56652 37706 56704
rect 1104 56602 58880 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 58880 56602
rect 1104 56528 58880 56550
rect 382 56448 388 56500
rect 440 56488 446 56500
rect 1302 56488 1308 56500
rect 440 56460 1308 56488
rect 440 56448 446 56460
rect 1302 56448 1308 56460
rect 1360 56448 1366 56500
rect 3234 56448 3240 56500
rect 3292 56488 3298 56500
rect 3789 56491 3847 56497
rect 3789 56488 3801 56491
rect 3292 56460 3801 56488
rect 3292 56448 3298 56460
rect 3789 56457 3801 56460
rect 3835 56457 3847 56491
rect 4798 56488 4804 56500
rect 4759 56460 4804 56488
rect 3789 56451 3847 56457
rect 4798 56448 4804 56460
rect 4856 56448 4862 56500
rect 22833 56491 22891 56497
rect 22833 56457 22845 56491
rect 22879 56488 22891 56491
rect 23382 56488 23388 56500
rect 22879 56460 23388 56488
rect 22879 56457 22891 56460
rect 22833 56451 22891 56457
rect 23382 56448 23388 56460
rect 23440 56448 23446 56500
rect 24578 56448 24584 56500
rect 24636 56488 24642 56500
rect 24857 56491 24915 56497
rect 24857 56488 24869 56491
rect 24636 56460 24869 56488
rect 24636 56448 24642 56460
rect 24857 56457 24869 56460
rect 24903 56457 24915 56491
rect 24857 56451 24915 56457
rect 26326 56448 26332 56500
rect 26384 56488 26390 56500
rect 26697 56491 26755 56497
rect 26697 56488 26709 56491
rect 26384 56460 26709 56488
rect 26384 56448 26390 56460
rect 26697 56457 26709 56460
rect 26743 56457 26755 56491
rect 26697 56451 26755 56457
rect 26786 56448 26792 56500
rect 26844 56488 26850 56500
rect 26844 56460 31248 56488
rect 26844 56448 26850 56460
rect 2685 56423 2743 56429
rect 2685 56389 2697 56423
rect 2731 56420 2743 56423
rect 3326 56420 3332 56432
rect 2731 56392 3332 56420
rect 2731 56389 2743 56392
rect 2685 56383 2743 56389
rect 3326 56380 3332 56392
rect 3384 56380 3390 56432
rect 3697 56423 3755 56429
rect 3697 56389 3709 56423
rect 3743 56420 3755 56423
rect 4246 56420 4252 56432
rect 3743 56392 4252 56420
rect 3743 56389 3755 56392
rect 3697 56383 3755 56389
rect 4246 56380 4252 56392
rect 4304 56380 4310 56432
rect 11790 56380 11796 56432
rect 11848 56420 11854 56432
rect 12161 56423 12219 56429
rect 12161 56420 12173 56423
rect 11848 56392 12173 56420
rect 11848 56380 11854 56392
rect 12161 56389 12173 56392
rect 12207 56389 12219 56423
rect 31220 56420 31248 56460
rect 31294 56448 31300 56500
rect 31352 56488 31358 56500
rect 31481 56491 31539 56497
rect 31481 56488 31493 56491
rect 31352 56460 31493 56488
rect 31352 56448 31358 56460
rect 31481 56457 31493 56460
rect 31527 56457 31539 56491
rect 31481 56451 31539 56457
rect 31938 56448 31944 56500
rect 31996 56488 32002 56500
rect 33042 56488 33048 56500
rect 31996 56460 33048 56488
rect 31996 56448 32002 56460
rect 33042 56448 33048 56460
rect 33100 56448 33106 56500
rect 33226 56497 33232 56500
rect 33210 56491 33232 56497
rect 33210 56457 33222 56491
rect 33210 56451 33232 56457
rect 33226 56448 33232 56451
rect 33284 56448 33290 56500
rect 33321 56491 33379 56497
rect 33321 56457 33333 56491
rect 33367 56488 33379 56491
rect 34698 56488 34704 56500
rect 33367 56460 34704 56488
rect 33367 56457 33379 56460
rect 33321 56451 33379 56457
rect 34698 56448 34704 56460
rect 34756 56448 34762 56500
rect 34977 56491 35035 56497
rect 34977 56457 34989 56491
rect 35023 56488 35035 56491
rect 35250 56488 35256 56500
rect 35023 56460 35256 56488
rect 35023 56457 35035 56460
rect 34977 56451 35035 56457
rect 35250 56448 35256 56460
rect 35308 56448 35314 56500
rect 38930 56488 38936 56500
rect 35544 56460 38936 56488
rect 33505 56423 33563 56429
rect 33505 56420 33517 56423
rect 31220 56392 33517 56420
rect 12161 56383 12219 56389
rect 33505 56389 33517 56392
rect 33551 56389 33563 56423
rect 33505 56383 33563 56389
rect 34422 56380 34428 56432
rect 34480 56420 34486 56432
rect 35544 56420 35572 56460
rect 38930 56448 38936 56460
rect 38988 56448 38994 56500
rect 54205 56491 54263 56497
rect 54205 56457 54217 56491
rect 54251 56488 54263 56491
rect 54754 56488 54760 56500
rect 54251 56460 54760 56488
rect 54251 56457 54263 56460
rect 54205 56451 54263 56457
rect 54754 56448 54760 56460
rect 54812 56448 54818 56500
rect 55125 56491 55183 56497
rect 55125 56457 55137 56491
rect 55171 56488 55183 56491
rect 56410 56488 56416 56500
rect 55171 56460 56416 56488
rect 55171 56457 55183 56460
rect 55125 56451 55183 56457
rect 56410 56448 56416 56460
rect 56468 56448 56474 56500
rect 56502 56448 56508 56500
rect 56560 56488 56566 56500
rect 59538 56488 59544 56500
rect 56560 56460 59544 56488
rect 56560 56448 56566 56460
rect 59538 56448 59544 56460
rect 59596 56448 59602 56500
rect 34480 56392 35572 56420
rect 34480 56380 34486 56392
rect 35618 56380 35624 56432
rect 35676 56380 35682 56432
rect 53926 56380 53932 56432
rect 53984 56420 53990 56432
rect 54662 56420 54668 56432
rect 53984 56392 54668 56420
rect 53984 56380 53990 56392
rect 54662 56380 54668 56392
rect 54720 56380 54726 56432
rect 56134 56380 56140 56432
rect 56192 56420 56198 56432
rect 58066 56420 58072 56432
rect 56192 56392 58072 56420
rect 56192 56380 56198 56392
rect 58066 56380 58072 56392
rect 58124 56380 58130 56432
rect 1118 56312 1124 56364
rect 1176 56352 1182 56364
rect 3881 56355 3939 56361
rect 1176 56324 2084 56352
rect 1176 56312 1182 56324
rect 1210 56244 1216 56296
rect 1268 56284 1274 56296
rect 2056 56293 2084 56324
rect 3881 56321 3893 56355
rect 3927 56352 3939 56355
rect 4614 56352 4620 56364
rect 3927 56324 4620 56352
rect 3927 56321 3939 56324
rect 3881 56315 3939 56321
rect 4614 56312 4620 56324
rect 4672 56312 4678 56364
rect 11974 56312 11980 56364
rect 12032 56352 12038 56364
rect 33410 56352 33416 56364
rect 12032 56324 12388 56352
rect 33371 56324 33416 56352
rect 12032 56312 12038 56324
rect 1397 56287 1455 56293
rect 1397 56284 1409 56287
rect 1268 56256 1409 56284
rect 1268 56244 1274 56256
rect 1397 56253 1409 56256
rect 1443 56253 1455 56287
rect 1397 56247 1455 56253
rect 2041 56287 2099 56293
rect 2041 56253 2053 56287
rect 2087 56253 2099 56287
rect 2041 56247 2099 56253
rect 2682 56244 2688 56296
rect 2740 56284 2746 56296
rect 2869 56287 2927 56293
rect 2869 56284 2881 56287
rect 2740 56256 2881 56284
rect 2740 56244 2746 56256
rect 2869 56253 2881 56256
rect 2915 56253 2927 56287
rect 2869 56247 2927 56253
rect 4985 56287 5043 56293
rect 4985 56253 4997 56287
rect 5031 56284 5043 56287
rect 5258 56284 5264 56296
rect 5031 56256 5264 56284
rect 5031 56253 5043 56256
rect 4985 56247 5043 56253
rect 5258 56244 5264 56256
rect 5316 56244 5322 56296
rect 11238 56244 11244 56296
rect 11296 56284 11302 56296
rect 12066 56284 12072 56296
rect 11296 56256 12072 56284
rect 11296 56244 11302 56256
rect 12066 56244 12072 56256
rect 12124 56244 12130 56296
rect 12360 56293 12388 56324
rect 33410 56312 33416 56324
rect 33468 56312 33474 56364
rect 34526 56355 34584 56361
rect 34526 56352 34538 56355
rect 34348 56324 34538 56352
rect 12345 56287 12403 56293
rect 12345 56253 12357 56287
rect 12391 56253 12403 56287
rect 12345 56247 12403 56253
rect 23017 56287 23075 56293
rect 23017 56253 23029 56287
rect 23063 56284 23075 56287
rect 23198 56284 23204 56296
rect 23063 56256 23204 56284
rect 23063 56253 23075 56256
rect 23017 56247 23075 56253
rect 23198 56244 23204 56256
rect 23256 56244 23262 56296
rect 23382 56244 23388 56296
rect 23440 56284 23446 56296
rect 23477 56287 23535 56293
rect 23477 56284 23489 56287
rect 23440 56256 23489 56284
rect 23440 56244 23446 56256
rect 23477 56253 23489 56256
rect 23523 56253 23535 56287
rect 23477 56247 23535 56253
rect 23744 56287 23802 56293
rect 23744 56253 23756 56287
rect 23790 56284 23802 56287
rect 24118 56284 24124 56296
rect 23790 56256 24124 56284
rect 23790 56253 23802 56256
rect 23744 56247 23802 56253
rect 24118 56244 24124 56256
rect 24176 56244 24182 56296
rect 25314 56284 25320 56296
rect 25275 56256 25320 56284
rect 25314 56244 25320 56256
rect 25372 56244 25378 56296
rect 25590 56293 25596 56296
rect 25584 56284 25596 56293
rect 25551 56256 25596 56284
rect 25584 56247 25596 56256
rect 25590 56244 25596 56247
rect 25648 56244 25654 56296
rect 27801 56287 27859 56293
rect 27801 56253 27813 56287
rect 27847 56284 27859 56287
rect 29086 56284 29092 56296
rect 27847 56256 29092 56284
rect 27847 56253 27859 56256
rect 27801 56247 27859 56253
rect 29086 56244 29092 56256
rect 29144 56284 29150 56296
rect 29641 56287 29699 56293
rect 29641 56284 29653 56287
rect 29144 56256 29653 56284
rect 29144 56244 29150 56256
rect 29641 56253 29653 56256
rect 29687 56253 29699 56287
rect 31662 56284 31668 56296
rect 31623 56256 31668 56284
rect 29641 56247 29699 56253
rect 31662 56244 31668 56256
rect 31720 56244 31726 56296
rect 32122 56284 32128 56296
rect 32083 56256 32128 56284
rect 32122 56244 32128 56256
rect 32180 56244 32186 56296
rect 32582 56244 32588 56296
rect 32640 56284 32646 56296
rect 34241 56287 34299 56293
rect 34241 56284 34253 56287
rect 32640 56256 34253 56284
rect 32640 56244 32646 56256
rect 34241 56253 34253 56256
rect 34287 56253 34299 56287
rect 34241 56247 34299 56253
rect 12710 56176 12716 56228
rect 12768 56216 12774 56228
rect 12805 56219 12863 56225
rect 12805 56216 12817 56219
rect 12768 56188 12817 56216
rect 12768 56176 12774 56188
rect 12805 56185 12817 56188
rect 12851 56185 12863 56219
rect 12805 56179 12863 56185
rect 27890 56176 27896 56228
rect 27948 56216 27954 56228
rect 28046 56219 28104 56225
rect 28046 56216 28058 56219
rect 27948 56188 28058 56216
rect 27948 56176 27954 56188
rect 28046 56185 28058 56188
rect 28092 56185 28104 56219
rect 29908 56219 29966 56225
rect 28046 56179 28104 56185
rect 28920 56188 29868 56216
rect 4154 56148 4160 56160
rect 4115 56120 4160 56148
rect 4154 56108 4160 56120
rect 4212 56108 4218 56160
rect 27338 56108 27344 56160
rect 27396 56148 27402 56160
rect 28920 56148 28948 56188
rect 27396 56120 28948 56148
rect 27396 56108 27402 56120
rect 28994 56108 29000 56160
rect 29052 56148 29058 56160
rect 29181 56151 29239 56157
rect 29181 56148 29193 56151
rect 29052 56120 29193 56148
rect 29052 56108 29058 56120
rect 29181 56117 29193 56120
rect 29227 56117 29239 56151
rect 29840 56148 29868 56188
rect 29908 56185 29920 56219
rect 29954 56216 29966 56219
rect 30466 56216 30472 56228
rect 29954 56188 30472 56216
rect 29954 56185 29966 56188
rect 29908 56179 29966 56185
rect 30466 56176 30472 56188
rect 30524 56176 30530 56228
rect 31386 56176 31392 56228
rect 31444 56216 31450 56228
rect 32030 56225 32036 56228
rect 31757 56219 31815 56225
rect 31757 56216 31769 56219
rect 31444 56188 31769 56216
rect 31444 56176 31450 56188
rect 31757 56185 31769 56188
rect 31803 56185 31815 56219
rect 31757 56179 31815 56185
rect 31849 56219 31907 56225
rect 31849 56185 31861 56219
rect 31895 56185 31907 56219
rect 31849 56179 31907 56185
rect 31987 56219 32036 56225
rect 31987 56185 31999 56219
rect 32033 56185 32036 56219
rect 31987 56179 32036 56185
rect 30834 56148 30840 56160
rect 29840 56120 30840 56148
rect 29181 56111 29239 56117
rect 30834 56108 30840 56120
rect 30892 56108 30898 56160
rect 31021 56151 31079 56157
rect 31021 56117 31033 56151
rect 31067 56148 31079 56151
rect 31570 56148 31576 56160
rect 31067 56120 31576 56148
rect 31067 56117 31079 56120
rect 31021 56111 31079 56117
rect 31570 56108 31576 56120
rect 31628 56148 31634 56160
rect 31864 56148 31892 56179
rect 32030 56176 32036 56179
rect 32088 56176 32094 56228
rect 33042 56216 33048 56228
rect 33003 56188 33048 56216
rect 33042 56176 33048 56188
rect 33100 56176 33106 56228
rect 33410 56176 33416 56228
rect 33468 56216 33474 56228
rect 34348 56216 34376 56324
rect 34526 56321 34538 56324
rect 34572 56321 34584 56355
rect 34526 56315 34584 56321
rect 34422 56244 34428 56296
rect 34480 56284 34486 56296
rect 34609 56287 34667 56293
rect 34480 56256 34525 56284
rect 34480 56244 34486 56256
rect 34609 56253 34621 56287
rect 34655 56284 34667 56287
rect 34790 56284 34796 56296
rect 34655 56253 34684 56284
rect 34751 56256 34796 56284
rect 34609 56247 34684 56253
rect 33468 56188 34376 56216
rect 33468 56176 33474 56188
rect 34514 56176 34520 56228
rect 34572 56216 34578 56228
rect 34656 56216 34684 56247
rect 34790 56244 34796 56256
rect 34848 56244 34854 56296
rect 35636 56293 35664 56380
rect 55766 56352 55772 56364
rect 55727 56324 55772 56352
rect 55766 56312 55772 56324
rect 55824 56312 55830 56364
rect 56226 56352 56232 56364
rect 56187 56324 56232 56352
rect 56226 56312 56232 56324
rect 56284 56312 56290 56364
rect 35621 56287 35679 56293
rect 35621 56253 35633 56287
rect 35667 56253 35679 56287
rect 36262 56284 36268 56296
rect 36223 56256 36268 56284
rect 35621 56247 35679 56253
rect 36262 56244 36268 56256
rect 36320 56244 36326 56296
rect 51813 56287 51871 56293
rect 51813 56253 51825 56287
rect 51859 56253 51871 56287
rect 52454 56284 52460 56296
rect 52415 56256 52460 56284
rect 51813 56247 51871 56253
rect 34572 56188 34684 56216
rect 34572 56176 34578 56188
rect 31628 56120 31892 56148
rect 31628 56108 31634 56120
rect 34974 56108 34980 56160
rect 35032 56148 35038 56160
rect 35437 56151 35495 56157
rect 35437 56148 35449 56151
rect 35032 56120 35449 56148
rect 35032 56108 35038 56120
rect 35437 56117 35449 56120
rect 35483 56117 35495 56151
rect 36078 56148 36084 56160
rect 36039 56120 36084 56148
rect 35437 56111 35495 56117
rect 36078 56108 36084 56120
rect 36136 56108 36142 56160
rect 51828 56148 51856 56247
rect 52454 56244 52460 56256
rect 52512 56244 52518 56296
rect 54294 56244 54300 56296
rect 54352 56284 54358 56296
rect 54389 56287 54447 56293
rect 54389 56284 54401 56287
rect 54352 56256 54401 56284
rect 54352 56244 54358 56256
rect 54389 56253 54401 56256
rect 54435 56253 54447 56287
rect 54389 56247 54447 56253
rect 55309 56287 55367 56293
rect 55309 56253 55321 56287
rect 55355 56253 55367 56287
rect 55309 56247 55367 56253
rect 55324 56216 55352 56247
rect 55953 56219 56011 56225
rect 55953 56216 55965 56219
rect 55324 56188 55965 56216
rect 55953 56185 55965 56188
rect 55999 56216 56011 56219
rect 56686 56216 56692 56228
rect 55999 56188 56692 56216
rect 55999 56185 56011 56188
rect 55953 56179 56011 56185
rect 56686 56176 56692 56188
rect 56744 56176 56750 56228
rect 58710 56148 58716 56160
rect 51828 56120 58716 56148
rect 58710 56108 58716 56120
rect 58768 56108 58774 56160
rect 1104 56058 58880 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 50326 56058
rect 50378 56006 50390 56058
rect 50442 56006 50454 56058
rect 50506 56006 50518 56058
rect 50570 56006 58880 56058
rect 1104 55984 58880 56006
rect 2225 55947 2283 55953
rect 2225 55913 2237 55947
rect 2271 55944 2283 55947
rect 3142 55944 3148 55956
rect 2271 55916 3148 55944
rect 2271 55913 2283 55916
rect 2225 55907 2283 55913
rect 3142 55904 3148 55916
rect 3200 55904 3206 55956
rect 4154 55904 4160 55956
rect 4212 55944 4218 55956
rect 13354 55944 13360 55956
rect 4212 55916 13360 55944
rect 4212 55904 4218 55916
rect 13354 55904 13360 55916
rect 13412 55904 13418 55956
rect 24302 55944 24308 55956
rect 24263 55916 24308 55944
rect 24302 55904 24308 55916
rect 24360 55944 24366 55956
rect 25958 55944 25964 55956
rect 24360 55916 25452 55944
rect 25919 55916 25964 55944
rect 24360 55904 24366 55916
rect 25317 55879 25375 55885
rect 25317 55876 25329 55879
rect 24228 55848 25329 55876
rect 24228 55820 24256 55848
rect 25317 55845 25329 55848
rect 25363 55845 25375 55879
rect 25317 55839 25375 55845
rect 1394 55808 1400 55820
rect 1355 55780 1400 55808
rect 1394 55768 1400 55780
rect 1452 55768 1458 55820
rect 1946 55768 1952 55820
rect 2004 55808 2010 55820
rect 2041 55811 2099 55817
rect 2041 55808 2053 55811
rect 2004 55780 2053 55808
rect 2004 55768 2010 55780
rect 2041 55777 2053 55780
rect 2087 55777 2099 55811
rect 2041 55771 2099 55777
rect 3510 55768 3516 55820
rect 3568 55808 3574 55820
rect 4433 55811 4491 55817
rect 4433 55808 4445 55811
rect 3568 55780 4445 55808
rect 3568 55768 3574 55780
rect 4433 55777 4445 55780
rect 4479 55777 4491 55811
rect 4433 55771 4491 55777
rect 24121 55811 24179 55817
rect 24121 55777 24133 55811
rect 24167 55808 24179 55811
rect 24210 55808 24216 55820
rect 24167 55780 24216 55808
rect 24167 55777 24179 55780
rect 24121 55771 24179 55777
rect 24210 55768 24216 55780
rect 24268 55768 24274 55820
rect 24305 55811 24363 55817
rect 24305 55777 24317 55811
rect 24351 55808 24363 55811
rect 24578 55808 24584 55820
rect 24351 55780 24584 55808
rect 24351 55777 24363 55780
rect 24305 55771 24363 55777
rect 24578 55768 24584 55780
rect 24636 55768 24642 55820
rect 25222 55808 25228 55820
rect 25183 55780 25228 55808
rect 25222 55768 25228 55780
rect 25280 55768 25286 55820
rect 25424 55808 25452 55916
rect 25958 55904 25964 55916
rect 26016 55904 26022 55956
rect 27890 55944 27896 55956
rect 27851 55916 27896 55944
rect 27890 55904 27896 55916
rect 27948 55904 27954 55956
rect 30466 55944 30472 55956
rect 30427 55916 30472 55944
rect 30466 55904 30472 55916
rect 30524 55904 30530 55956
rect 31573 55947 31631 55953
rect 31573 55913 31585 55947
rect 31619 55944 31631 55947
rect 32122 55944 32128 55956
rect 31619 55916 32128 55944
rect 31619 55913 31631 55916
rect 31573 55907 31631 55913
rect 28905 55879 28963 55885
rect 28905 55876 28917 55879
rect 28092 55848 28917 55876
rect 25869 55811 25927 55817
rect 25869 55808 25881 55811
rect 25424 55780 25881 55808
rect 25869 55777 25881 55780
rect 25915 55777 25927 55811
rect 25869 55771 25927 55777
rect 26697 55811 26755 55817
rect 26697 55777 26709 55811
rect 26743 55808 26755 55811
rect 27890 55808 27896 55820
rect 26743 55780 27896 55808
rect 26743 55777 26755 55780
rect 26697 55771 26755 55777
rect 27890 55768 27896 55780
rect 27948 55768 27954 55820
rect 27982 55768 27988 55820
rect 28040 55808 28046 55820
rect 28092 55817 28120 55848
rect 28905 55845 28917 55848
rect 28951 55845 28963 55879
rect 31588 55876 31616 55907
rect 32122 55904 32128 55916
rect 32180 55904 32186 55956
rect 32585 55947 32643 55953
rect 32585 55913 32597 55947
rect 32631 55944 32643 55947
rect 33134 55944 33140 55956
rect 32631 55916 33140 55944
rect 32631 55913 32643 55916
rect 32585 55907 32643 55913
rect 33134 55904 33140 55916
rect 33192 55904 33198 55956
rect 33226 55904 33232 55956
rect 33284 55944 33290 55956
rect 35713 55947 35771 55953
rect 35713 55944 35725 55947
rect 33284 55916 35725 55944
rect 33284 55904 33290 55916
rect 35713 55913 35725 55916
rect 35759 55913 35771 55947
rect 56778 55944 56784 55956
rect 56739 55916 56784 55944
rect 35713 55907 35771 55913
rect 56778 55904 56784 55916
rect 56836 55904 56842 55956
rect 28905 55839 28963 55845
rect 30760 55848 31616 55876
rect 28077 55811 28135 55817
rect 28077 55808 28089 55811
rect 28040 55780 28089 55808
rect 28040 55768 28046 55780
rect 28077 55777 28089 55780
rect 28123 55777 28135 55811
rect 28077 55771 28135 55777
rect 28258 55768 28264 55820
rect 28316 55808 28322 55820
rect 28813 55811 28871 55817
rect 28813 55808 28825 55811
rect 28316 55780 28825 55808
rect 28316 55768 28322 55780
rect 28813 55777 28825 55780
rect 28859 55777 28871 55811
rect 28994 55808 29000 55820
rect 28955 55780 29000 55808
rect 28813 55771 28871 55777
rect 28994 55768 29000 55780
rect 29052 55768 29058 55820
rect 30653 55811 30711 55817
rect 30653 55777 30665 55811
rect 30699 55808 30711 55811
rect 30760 55808 30788 55848
rect 32030 55836 32036 55888
rect 32088 55876 32094 55888
rect 32677 55879 32735 55885
rect 32677 55876 32689 55879
rect 32088 55848 32689 55876
rect 32088 55836 32094 55848
rect 32677 55845 32689 55848
rect 32723 55845 32735 55879
rect 34790 55876 34796 55888
rect 32677 55839 32735 55845
rect 32876 55848 34796 55876
rect 31386 55808 31392 55820
rect 30699 55780 30788 55808
rect 30852 55780 31392 55808
rect 30699 55777 30711 55780
rect 30653 55771 30711 55777
rect 1854 55700 1860 55752
rect 1912 55740 1918 55752
rect 26973 55743 27031 55749
rect 1912 55712 6914 55740
rect 1912 55700 1918 55712
rect 4246 55672 4252 55684
rect 4207 55644 4252 55672
rect 4246 55632 4252 55644
rect 4304 55632 4310 55684
rect 6886 55672 6914 55712
rect 26973 55709 26985 55743
rect 27019 55740 27031 55743
rect 27430 55740 27436 55752
rect 27019 55712 27436 55740
rect 27019 55709 27031 55712
rect 26973 55703 27031 55709
rect 27430 55700 27436 55712
rect 27488 55700 27494 55752
rect 28353 55743 28411 55749
rect 28353 55709 28365 55743
rect 28399 55740 28411 55743
rect 29012 55740 29040 55768
rect 28399 55712 29040 55740
rect 28399 55709 28411 55712
rect 28353 55703 28411 55709
rect 30374 55700 30380 55752
rect 30432 55740 30438 55752
rect 30852 55749 30880 55780
rect 31386 55768 31392 55780
rect 31444 55768 31450 55820
rect 31570 55808 31576 55820
rect 31531 55780 31576 55808
rect 31570 55768 31576 55780
rect 31628 55768 31634 55820
rect 30837 55743 30895 55749
rect 30837 55740 30849 55743
rect 30432 55712 30849 55740
rect 30432 55700 30438 55712
rect 30837 55709 30849 55712
rect 30883 55709 30895 55743
rect 30837 55703 30895 55709
rect 30929 55743 30987 55749
rect 30929 55709 30941 55743
rect 30975 55740 30987 55743
rect 31588 55740 31616 55768
rect 32876 55749 32904 55848
rect 34790 55836 34796 55848
rect 34848 55836 34854 55888
rect 57238 55876 57244 55888
rect 52564 55848 57244 55876
rect 33686 55817 33692 55820
rect 33680 55771 33692 55817
rect 33744 55808 33750 55820
rect 33744 55780 33780 55808
rect 33686 55768 33692 55771
rect 33744 55768 33750 55780
rect 34146 55768 34152 55820
rect 34204 55808 34210 55820
rect 52564 55817 52592 55848
rect 57238 55836 57244 55848
rect 57296 55836 57302 55888
rect 35897 55811 35955 55817
rect 35897 55808 35909 55811
rect 34204 55780 35909 55808
rect 34204 55768 34210 55780
rect 35897 55777 35909 55780
rect 35943 55777 35955 55811
rect 35897 55771 35955 55777
rect 52549 55811 52607 55817
rect 52549 55777 52561 55811
rect 52595 55777 52607 55811
rect 53190 55808 53196 55820
rect 53151 55780 53196 55808
rect 52549 55771 52607 55777
rect 53190 55768 53196 55780
rect 53248 55768 53254 55820
rect 53837 55811 53895 55817
rect 53837 55777 53849 55811
rect 53883 55808 53895 55811
rect 54018 55808 54024 55820
rect 53883 55780 54024 55808
rect 53883 55777 53895 55780
rect 53837 55771 53895 55777
rect 54018 55768 54024 55780
rect 54076 55768 54082 55820
rect 54570 55768 54576 55820
rect 54628 55808 54634 55820
rect 54665 55811 54723 55817
rect 54665 55808 54677 55811
rect 54628 55780 54677 55808
rect 54628 55768 54634 55780
rect 54665 55777 54677 55780
rect 54711 55777 54723 55811
rect 54665 55771 54723 55777
rect 55769 55811 55827 55817
rect 55769 55777 55781 55811
rect 55815 55808 55827 55811
rect 56594 55808 56600 55820
rect 55815 55780 56600 55808
rect 55815 55777 55827 55780
rect 55769 55771 55827 55777
rect 56594 55768 56600 55780
rect 56652 55768 56658 55820
rect 56686 55768 56692 55820
rect 56744 55808 56750 55820
rect 56965 55811 57023 55817
rect 56965 55808 56977 55811
rect 56744 55780 56977 55808
rect 56744 55768 56750 55780
rect 56965 55777 56977 55780
rect 57011 55777 57023 55811
rect 56965 55771 57023 55777
rect 30975 55712 31616 55740
rect 32861 55743 32919 55749
rect 30975 55709 30987 55712
rect 30929 55703 30987 55709
rect 32861 55709 32873 55743
rect 32907 55709 32919 55743
rect 32861 55703 32919 55709
rect 33226 55700 33232 55752
rect 33284 55740 33290 55752
rect 33413 55743 33471 55749
rect 33413 55740 33425 55743
rect 33284 55712 33425 55740
rect 33284 55700 33290 55712
rect 33413 55709 33425 55712
rect 33459 55709 33471 55743
rect 33413 55703 33471 55709
rect 56042 55700 56048 55752
rect 56100 55740 56106 55752
rect 57517 55743 57575 55749
rect 57517 55740 57529 55743
rect 56100 55712 57529 55740
rect 56100 55700 56106 55712
rect 57517 55709 57529 55712
rect 57563 55709 57575 55743
rect 57698 55740 57704 55752
rect 57659 55712 57704 55740
rect 57517 55703 57575 55709
rect 57698 55700 57704 55712
rect 57756 55700 57762 55752
rect 56226 55672 56232 55684
rect 6886 55644 33456 55672
rect 26510 55604 26516 55616
rect 26471 55576 26516 55604
rect 26510 55564 26516 55576
rect 26568 55564 26574 55616
rect 26878 55604 26884 55616
rect 26839 55576 26884 55604
rect 26878 55564 26884 55576
rect 26936 55564 26942 55616
rect 28258 55604 28264 55616
rect 28219 55576 28264 55604
rect 28258 55564 28264 55576
rect 28316 55564 28322 55616
rect 28718 55564 28724 55616
rect 28776 55604 28782 55616
rect 31938 55604 31944 55616
rect 28776 55576 31944 55604
rect 28776 55564 28782 55576
rect 31938 55564 31944 55576
rect 31996 55564 32002 55616
rect 32214 55604 32220 55616
rect 32175 55576 32220 55604
rect 32214 55564 32220 55576
rect 32272 55564 32278 55616
rect 33428 55604 33456 55644
rect 34348 55644 56232 55672
rect 34348 55604 34376 55644
rect 56226 55632 56232 55644
rect 56284 55632 56290 55684
rect 34790 55604 34796 55616
rect 33428 55576 34376 55604
rect 34751 55576 34796 55604
rect 34790 55564 34796 55576
rect 34848 55564 34854 55616
rect 57974 55604 57980 55616
rect 57935 55576 57980 55604
rect 57974 55564 57980 55576
rect 58032 55564 58038 55616
rect 1104 55514 58880 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 58880 55514
rect 1104 55440 58880 55462
rect 30834 55360 30840 55412
rect 30892 55400 30898 55412
rect 56042 55400 56048 55412
rect 30892 55372 32812 55400
rect 56003 55372 56048 55400
rect 30892 55360 30898 55372
rect 22830 55292 22836 55344
rect 22888 55332 22894 55344
rect 23382 55332 23388 55344
rect 22888 55304 23388 55332
rect 22888 55292 22894 55304
rect 23382 55292 23388 55304
rect 23440 55332 23446 55344
rect 32784 55332 32812 55372
rect 56042 55360 56048 55372
rect 56100 55360 56106 55412
rect 57330 55400 57336 55412
rect 57291 55372 57336 55400
rect 57330 55360 57336 55372
rect 57388 55360 57394 55412
rect 33502 55332 33508 55344
rect 23440 55304 23796 55332
rect 32784 55304 33508 55332
rect 23440 55292 23446 55304
rect 23768 55273 23796 55304
rect 33502 55292 33508 55304
rect 33560 55292 33566 55344
rect 34514 55332 34520 55344
rect 33796 55304 34520 55332
rect 23753 55267 23811 55273
rect 23753 55233 23765 55267
rect 23799 55233 23811 55267
rect 23753 55227 23811 55233
rect 24762 55224 24768 55276
rect 24820 55264 24826 55276
rect 32030 55264 32036 55276
rect 24820 55236 25820 55264
rect 31991 55236 32036 55264
rect 24820 55224 24826 55236
rect 22741 55199 22799 55205
rect 22741 55165 22753 55199
rect 22787 55165 22799 55199
rect 22922 55196 22928 55208
rect 22883 55168 22928 55196
rect 22741 55159 22799 55165
rect 22756 55128 22784 55159
rect 22922 55156 22928 55168
rect 22980 55156 22986 55208
rect 23017 55199 23075 55205
rect 23017 55165 23029 55199
rect 23063 55196 23075 55199
rect 23382 55196 23388 55208
rect 23063 55168 23388 55196
rect 23063 55165 23075 55168
rect 23017 55159 23075 55165
rect 23382 55156 23388 55168
rect 23440 55156 23446 55208
rect 25792 55205 25820 55236
rect 32030 55224 32036 55236
rect 32088 55224 32094 55276
rect 32858 55224 32864 55276
rect 32916 55264 32922 55276
rect 33410 55264 33416 55276
rect 32916 55236 33416 55264
rect 32916 55224 32922 55236
rect 33410 55224 33416 55236
rect 33468 55224 33474 55276
rect 33796 55264 33824 55304
rect 34514 55292 34520 55304
rect 34572 55292 34578 55344
rect 56505 55335 56563 55341
rect 56505 55301 56517 55335
rect 56551 55332 56563 55335
rect 57698 55332 57704 55344
rect 56551 55304 57704 55332
rect 56551 55301 56563 55304
rect 56505 55295 56563 55301
rect 57698 55292 57704 55304
rect 57756 55292 57762 55344
rect 58158 55332 58164 55344
rect 58119 55304 58164 55332
rect 58158 55292 58164 55304
rect 58216 55292 58222 55344
rect 33520 55236 33824 55264
rect 33520 55208 33548 55236
rect 33870 55224 33876 55276
rect 33928 55264 33934 55276
rect 33928 55236 33973 55264
rect 33928 55224 33934 55236
rect 34054 55224 34060 55276
rect 34112 55264 34118 55276
rect 34793 55267 34851 55273
rect 34793 55264 34805 55267
rect 34112 55236 34805 55264
rect 34112 55224 34118 55236
rect 34793 55233 34805 55236
rect 34839 55233 34851 55267
rect 34793 55227 34851 55233
rect 25777 55199 25835 55205
rect 25777 55165 25789 55199
rect 25823 55165 25835 55199
rect 25777 55159 25835 55165
rect 25866 55156 25872 55208
rect 25924 55196 25930 55208
rect 26421 55199 26479 55205
rect 26421 55196 26433 55199
rect 25924 55168 26433 55196
rect 25924 55156 25930 55168
rect 26421 55165 26433 55168
rect 26467 55165 26479 55199
rect 26421 55159 26479 55165
rect 26513 55199 26571 55205
rect 26513 55165 26525 55199
rect 26559 55196 26571 55199
rect 26878 55196 26884 55208
rect 26559 55168 26884 55196
rect 26559 55165 26571 55168
rect 26513 55159 26571 55165
rect 26878 55156 26884 55168
rect 26936 55196 26942 55208
rect 27801 55199 27859 55205
rect 27801 55196 27813 55199
rect 26936 55168 27813 55196
rect 26936 55156 26942 55168
rect 27801 55165 27813 55168
rect 27847 55165 27859 55199
rect 27801 55159 27859 55165
rect 27985 55199 28043 55205
rect 27985 55165 27997 55199
rect 28031 55165 28043 55199
rect 27985 55159 28043 55165
rect 23290 55128 23296 55140
rect 22756 55100 23296 55128
rect 23290 55088 23296 55100
rect 23348 55088 23354 55140
rect 23842 55088 23848 55140
rect 23900 55128 23906 55140
rect 23998 55131 24056 55137
rect 23998 55128 24010 55131
rect 23900 55100 24010 55128
rect 23900 55088 23906 55100
rect 23998 55097 24010 55100
rect 24044 55097 24056 55131
rect 27890 55128 27896 55140
rect 23998 55091 24056 55097
rect 24228 55100 25636 55128
rect 27851 55100 27896 55128
rect 22554 55060 22560 55072
rect 22515 55032 22560 55060
rect 22554 55020 22560 55032
rect 22612 55020 22618 55072
rect 23106 55020 23112 55072
rect 23164 55060 23170 55072
rect 24228 55060 24256 55100
rect 23164 55032 24256 55060
rect 23164 55020 23170 55032
rect 24302 55020 24308 55072
rect 24360 55060 24366 55072
rect 25608 55069 25636 55100
rect 27890 55088 27896 55100
rect 27948 55088 27954 55140
rect 25133 55063 25191 55069
rect 25133 55060 25145 55063
rect 24360 55032 25145 55060
rect 24360 55020 24366 55032
rect 25133 55029 25145 55032
rect 25179 55029 25191 55063
rect 25133 55023 25191 55029
rect 25593 55063 25651 55069
rect 25593 55029 25605 55063
rect 25639 55029 25651 55063
rect 25593 55023 25651 55029
rect 27430 55020 27436 55072
rect 27488 55060 27494 55072
rect 28000 55060 28028 55159
rect 28994 55156 29000 55208
rect 29052 55196 29058 55208
rect 31757 55199 31815 55205
rect 29052 55168 29097 55196
rect 29052 55156 29058 55168
rect 31757 55165 31769 55199
rect 31803 55196 31815 55199
rect 32214 55196 32220 55208
rect 31803 55168 32220 55196
rect 31803 55165 31815 55168
rect 31757 55159 31815 55165
rect 32214 55156 32220 55168
rect 32272 55156 32278 55208
rect 33157 55199 33215 55205
rect 33157 55165 33169 55199
rect 33203 55165 33215 55199
rect 33157 55159 33215 55165
rect 33321 55199 33379 55205
rect 33321 55165 33333 55199
rect 33367 55165 33379 55199
rect 33502 55196 33508 55208
rect 33463 55168 33508 55196
rect 33321 55159 33379 55165
rect 29086 55088 29092 55140
rect 29144 55128 29150 55140
rect 29242 55131 29300 55137
rect 29242 55128 29254 55131
rect 29144 55100 29254 55128
rect 29144 55088 29150 55100
rect 29242 55097 29254 55100
rect 29288 55097 29300 55131
rect 31849 55131 31907 55137
rect 31849 55128 31861 55131
rect 29242 55091 29300 55097
rect 30392 55100 31861 55128
rect 27488 55032 28028 55060
rect 27488 55020 27494 55032
rect 29546 55020 29552 55072
rect 29604 55060 29610 55072
rect 30392 55069 30420 55100
rect 31849 55097 31861 55100
rect 31895 55097 31907 55131
rect 31849 55091 31907 55097
rect 32582 55088 32588 55140
rect 32640 55128 32646 55140
rect 33172 55128 33200 55159
rect 32640 55100 33200 55128
rect 33336 55128 33364 55159
rect 33502 55156 33508 55168
rect 33560 55156 33566 55208
rect 33689 55199 33747 55205
rect 33689 55165 33701 55199
rect 33735 55196 33747 55199
rect 34698 55196 34704 55208
rect 33735 55168 34704 55196
rect 33735 55165 33747 55168
rect 33689 55159 33747 55165
rect 34698 55156 34704 55168
rect 34756 55156 34762 55208
rect 53926 55156 53932 55208
rect 53984 55196 53990 55208
rect 54573 55199 54631 55205
rect 54573 55196 54585 55199
rect 53984 55168 54585 55196
rect 53984 55156 53990 55168
rect 54573 55165 54585 55168
rect 54619 55165 54631 55199
rect 54573 55159 54631 55165
rect 55214 55156 55220 55208
rect 55272 55196 55278 55208
rect 56686 55196 56692 55208
rect 55272 55168 55317 55196
rect 56647 55168 56692 55196
rect 55272 55156 55278 55168
rect 56686 55156 56692 55168
rect 56744 55156 56750 55208
rect 57974 55196 57980 55208
rect 57935 55168 57980 55196
rect 57974 55156 57980 55168
rect 58032 55156 58038 55208
rect 34238 55128 34244 55140
rect 33336 55100 34244 55128
rect 32640 55088 32646 55100
rect 34238 55088 34244 55100
rect 34296 55088 34302 55140
rect 35060 55131 35118 55137
rect 35060 55097 35072 55131
rect 35106 55128 35118 55131
rect 35250 55128 35256 55140
rect 35106 55100 35256 55128
rect 35106 55097 35118 55100
rect 35060 55091 35118 55097
rect 35250 55088 35256 55100
rect 35308 55088 35314 55140
rect 57241 55131 57299 55137
rect 57241 55097 57253 55131
rect 57287 55128 57299 55131
rect 58526 55128 58532 55140
rect 57287 55100 58532 55128
rect 57287 55097 57299 55100
rect 57241 55091 57299 55097
rect 58526 55088 58532 55100
rect 58584 55088 58590 55140
rect 30377 55063 30435 55069
rect 30377 55060 30389 55063
rect 29604 55032 30389 55060
rect 29604 55020 29610 55032
rect 30377 55029 30389 55032
rect 30423 55029 30435 55063
rect 30377 55023 30435 55029
rect 31389 55063 31447 55069
rect 31389 55029 31401 55063
rect 31435 55060 31447 55063
rect 33410 55060 33416 55072
rect 31435 55032 33416 55060
rect 31435 55029 31447 55032
rect 31389 55023 31447 55029
rect 33410 55020 33416 55032
rect 33468 55020 33474 55072
rect 36170 55060 36176 55072
rect 36131 55032 36176 55060
rect 36170 55020 36176 55032
rect 36228 55020 36234 55072
rect 1104 54970 58880 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 50326 54970
rect 50378 54918 50390 54970
rect 50442 54918 50454 54970
rect 50506 54918 50518 54970
rect 50570 54918 58880 54970
rect 1104 54896 58880 54918
rect 23382 54856 23388 54868
rect 22066 54828 22692 54856
rect 23343 54828 23388 54856
rect 8294 54748 8300 54800
rect 8352 54788 8358 54800
rect 22066 54788 22094 54828
rect 8352 54760 22094 54788
rect 22272 54791 22330 54797
rect 8352 54748 8358 54760
rect 22272 54757 22284 54791
rect 22318 54788 22330 54791
rect 22554 54788 22560 54800
rect 22318 54760 22560 54788
rect 22318 54757 22330 54760
rect 22272 54751 22330 54757
rect 22554 54748 22560 54760
rect 22612 54748 22618 54800
rect 22664 54788 22692 54828
rect 23382 54816 23388 54828
rect 23440 54816 23446 54868
rect 23842 54856 23848 54868
rect 23803 54828 23848 54856
rect 23842 54816 23848 54828
rect 23900 54816 23906 54868
rect 27430 54856 27436 54868
rect 27391 54828 27436 54856
rect 27430 54816 27436 54828
rect 27488 54816 27494 54868
rect 27985 54859 28043 54865
rect 27985 54825 27997 54859
rect 28031 54856 28043 54859
rect 28258 54856 28264 54868
rect 28031 54828 28264 54856
rect 28031 54825 28043 54828
rect 27985 54819 28043 54825
rect 28258 54816 28264 54828
rect 28316 54816 28322 54868
rect 32030 54816 32036 54868
rect 32088 54856 32094 54868
rect 32125 54859 32183 54865
rect 32125 54856 32137 54859
rect 32088 54828 32137 54856
rect 32088 54816 32094 54828
rect 32125 54825 32137 54828
rect 32171 54825 32183 54859
rect 32125 54819 32183 54825
rect 26320 54791 26378 54797
rect 22664 54760 26280 54788
rect 1394 54720 1400 54732
rect 1355 54692 1400 54720
rect 1394 54680 1400 54692
rect 1452 54680 1458 54732
rect 22005 54723 22063 54729
rect 22005 54689 22017 54723
rect 22051 54720 22063 54723
rect 22094 54720 22100 54732
rect 22051 54692 22100 54720
rect 22051 54689 22063 54692
rect 22005 54683 22063 54689
rect 22094 54680 22100 54692
rect 22152 54720 22158 54732
rect 22830 54720 22836 54732
rect 22152 54692 22836 54720
rect 22152 54680 22158 54692
rect 22830 54680 22836 54692
rect 22888 54680 22894 54732
rect 24029 54723 24087 54729
rect 24029 54689 24041 54723
rect 24075 54689 24087 54723
rect 24302 54720 24308 54732
rect 24263 54692 24308 54720
rect 24029 54683 24087 54689
rect 24044 54652 24072 54683
rect 24302 54680 24308 54692
rect 24360 54680 24366 54732
rect 25314 54680 25320 54732
rect 25372 54720 25378 54732
rect 26053 54723 26111 54729
rect 26053 54720 26065 54723
rect 25372 54692 26065 54720
rect 25372 54680 25378 54692
rect 26053 54689 26065 54692
rect 26099 54720 26111 54723
rect 26142 54720 26148 54732
rect 26099 54692 26148 54720
rect 26099 54689 26111 54692
rect 26053 54683 26111 54689
rect 26142 54680 26148 54692
rect 26200 54680 26206 54732
rect 26252 54720 26280 54760
rect 26320 54757 26332 54791
rect 26366 54788 26378 54791
rect 26510 54788 26516 54800
rect 26366 54760 26516 54788
rect 26366 54757 26378 54760
rect 26320 54751 26378 54757
rect 26510 54748 26516 54760
rect 26568 54748 26574 54800
rect 31012 54791 31070 54797
rect 26620 54760 28856 54788
rect 26620 54720 26648 54760
rect 27890 54720 27896 54732
rect 26252 54692 26648 54720
rect 27851 54692 27896 54720
rect 27890 54680 27896 54692
rect 27948 54680 27954 54732
rect 28721 54723 28779 54729
rect 28721 54689 28733 54723
rect 28767 54689 28779 54723
rect 28828 54720 28856 54760
rect 31012 54757 31024 54791
rect 31058 54788 31070 54791
rect 31754 54788 31760 54800
rect 31058 54760 31760 54788
rect 31058 54757 31070 54760
rect 31012 54751 31070 54757
rect 31754 54748 31760 54760
rect 31812 54748 31818 54800
rect 32140 54788 32168 54819
rect 33134 54816 33140 54868
rect 33192 54856 33198 54868
rect 33781 54859 33839 54865
rect 33781 54856 33793 54859
rect 33192 54828 33793 54856
rect 33192 54816 33198 54828
rect 33781 54825 33793 54828
rect 33827 54825 33839 54859
rect 33781 54819 33839 54825
rect 58161 54859 58219 54865
rect 58161 54825 58173 54859
rect 58207 54856 58219 54859
rect 58342 54856 58348 54868
rect 58207 54828 58348 54856
rect 58207 54825 58219 54828
rect 58161 54819 58219 54825
rect 58342 54816 58348 54828
rect 58400 54816 58406 54868
rect 37642 54788 37648 54800
rect 32140 54760 33180 54788
rect 32582 54720 32588 54732
rect 28828 54692 32588 54720
rect 28721 54683 28779 54689
rect 25222 54652 25228 54664
rect 24044 54624 25228 54652
rect 25222 54612 25228 54624
rect 25280 54612 25286 54664
rect 28736 54584 28764 54683
rect 32582 54680 32588 54692
rect 32640 54680 32646 54732
rect 32769 54723 32827 54729
rect 32769 54689 32781 54723
rect 32815 54689 32827 54723
rect 32769 54683 32827 54689
rect 28997 54655 29055 54661
rect 28997 54621 29009 54655
rect 29043 54652 29055 54655
rect 29362 54652 29368 54664
rect 29043 54624 29368 54652
rect 29043 54621 29055 54624
rect 28997 54615 29055 54621
rect 29362 54612 29368 54624
rect 29420 54612 29426 54664
rect 30742 54652 30748 54664
rect 30703 54624 30748 54652
rect 30742 54612 30748 54624
rect 30800 54612 30806 54664
rect 32784 54652 32812 54683
rect 32858 54680 32864 54732
rect 32916 54720 32922 54732
rect 33042 54729 33048 54732
rect 32999 54723 33048 54729
rect 32916 54692 32961 54720
rect 32916 54680 32922 54692
rect 32999 54689 33011 54723
rect 33045 54689 33048 54723
rect 32999 54683 33048 54689
rect 33042 54680 33048 54683
rect 33100 54680 33106 54732
rect 33152 54729 33180 54760
rect 33980 54760 37648 54788
rect 33137 54723 33195 54729
rect 33137 54689 33149 54723
rect 33183 54689 33195 54723
rect 33137 54683 33195 54689
rect 33980 54652 34008 54760
rect 37642 54748 37648 54760
rect 37700 54748 37706 54800
rect 56134 54788 56140 54800
rect 54312 54760 56140 54788
rect 34146 54720 34152 54732
rect 34107 54692 34152 54720
rect 34146 54680 34152 54692
rect 34204 54680 34210 54732
rect 34241 54723 34299 54729
rect 34241 54689 34253 54723
rect 34287 54720 34299 54723
rect 36170 54720 36176 54732
rect 34287 54692 36176 54720
rect 34287 54689 34299 54692
rect 34241 54683 34299 54689
rect 36170 54680 36176 54692
rect 36228 54720 36234 54732
rect 54312 54729 54340 54760
rect 56134 54748 56140 54760
rect 56192 54748 56198 54800
rect 36817 54723 36875 54729
rect 36817 54720 36829 54723
rect 36228 54692 36829 54720
rect 36228 54680 36234 54692
rect 36817 54689 36829 54692
rect 36863 54689 36875 54723
rect 36817 54683 36875 54689
rect 54297 54723 54355 54729
rect 54297 54689 54309 54723
rect 54343 54689 54355 54723
rect 54297 54683 54355 54689
rect 54941 54723 54999 54729
rect 54941 54689 54953 54723
rect 54987 54720 54999 54723
rect 55306 54720 55312 54732
rect 54987 54692 55312 54720
rect 54987 54689 54999 54692
rect 54941 54683 54999 54689
rect 55306 54680 55312 54692
rect 55364 54680 55370 54732
rect 55582 54720 55588 54732
rect 55543 54692 55588 54720
rect 55582 54680 55588 54692
rect 55640 54680 55646 54732
rect 32784 54624 34008 54652
rect 34425 54655 34483 54661
rect 34425 54621 34437 54655
rect 34471 54652 34483 54655
rect 34790 54652 34796 54664
rect 34471 54624 34796 54652
rect 34471 54621 34483 54624
rect 34425 54615 34483 54621
rect 34790 54612 34796 54624
rect 34848 54612 34854 54664
rect 35713 54655 35771 54661
rect 35713 54652 35725 54655
rect 34900 54624 35725 54652
rect 29914 54584 29920 54596
rect 28736 54556 29920 54584
rect 29914 54544 29920 54556
rect 29972 54544 29978 54596
rect 23934 54476 23940 54528
rect 23992 54516 23998 54528
rect 24213 54519 24271 54525
rect 24213 54516 24225 54519
rect 23992 54488 24225 54516
rect 23992 54476 23998 54488
rect 24213 54485 24225 54488
rect 24259 54485 24271 54519
rect 28534 54516 28540 54528
rect 28495 54488 28540 54516
rect 24213 54479 24271 54485
rect 28534 54476 28540 54488
rect 28592 54476 28598 54528
rect 28902 54516 28908 54528
rect 28863 54488 28908 54516
rect 28902 54476 28908 54488
rect 28960 54476 28966 54528
rect 30760 54516 30788 54612
rect 31754 54544 31760 54596
rect 31812 54584 31818 54596
rect 33321 54587 33379 54593
rect 33321 54584 33333 54587
rect 31812 54556 33333 54584
rect 31812 54544 31818 54556
rect 33321 54553 33333 54556
rect 33367 54553 33379 54587
rect 33321 54547 33379 54553
rect 33686 54544 33692 54596
rect 33744 54584 33750 54596
rect 34900 54584 34928 54624
rect 35713 54621 35725 54624
rect 35759 54621 35771 54655
rect 35713 54615 35771 54621
rect 57057 54655 57115 54661
rect 57057 54621 57069 54655
rect 57103 54652 57115 54655
rect 57517 54655 57575 54661
rect 57517 54652 57529 54655
rect 57103 54624 57529 54652
rect 57103 54621 57115 54624
rect 57057 54615 57115 54621
rect 57517 54621 57529 54624
rect 57563 54621 57575 54655
rect 57698 54652 57704 54664
rect 57659 54624 57704 54652
rect 57517 54615 57575 54621
rect 57698 54612 57704 54624
rect 57756 54612 57762 54664
rect 33744 54556 34928 54584
rect 33744 54544 33750 54556
rect 35434 54544 35440 54596
rect 35492 54584 35498 54596
rect 36909 54587 36967 54593
rect 36909 54584 36921 54587
rect 35492 54556 36921 54584
rect 35492 54544 35498 54556
rect 36909 54553 36921 54556
rect 36955 54553 36967 54587
rect 36909 54547 36967 54553
rect 33226 54516 33232 54528
rect 30760 54488 33232 54516
rect 33226 54476 33232 54488
rect 33284 54476 33290 54528
rect 33870 54476 33876 54528
rect 33928 54516 33934 54528
rect 36357 54519 36415 54525
rect 36357 54516 36369 54519
rect 33928 54488 36369 54516
rect 33928 54476 33934 54488
rect 36357 54485 36369 54488
rect 36403 54485 36415 54519
rect 36357 54479 36415 54485
rect 1104 54426 58880 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 58880 54426
rect 1104 54352 58880 54374
rect 22649 54315 22707 54321
rect 22649 54281 22661 54315
rect 22695 54312 22707 54315
rect 22922 54312 22928 54324
rect 22695 54284 22928 54312
rect 22695 54281 22707 54284
rect 22649 54275 22707 54281
rect 22922 54272 22928 54284
rect 22980 54272 22986 54324
rect 23290 54312 23296 54324
rect 23251 54284 23296 54312
rect 23290 54272 23296 54284
rect 23348 54272 23354 54324
rect 23934 54312 23940 54324
rect 23895 54284 23940 54312
rect 23934 54272 23940 54284
rect 23992 54272 23998 54324
rect 24581 54315 24639 54321
rect 24581 54281 24593 54315
rect 24627 54312 24639 54315
rect 25222 54312 25228 54324
rect 24627 54284 25228 54312
rect 24627 54281 24639 54284
rect 24581 54275 24639 54281
rect 25222 54272 25228 54284
rect 25280 54272 25286 54324
rect 28997 54315 29055 54321
rect 28997 54281 29009 54315
rect 29043 54312 29055 54315
rect 29086 54312 29092 54324
rect 29043 54284 29092 54312
rect 29043 54281 29055 54284
rect 28997 54275 29055 54281
rect 29086 54272 29092 54284
rect 29144 54272 29150 54324
rect 31021 54315 31079 54321
rect 31021 54281 31033 54315
rect 31067 54312 31079 54315
rect 33686 54312 33692 54324
rect 31067 54284 33692 54312
rect 31067 54281 31079 54284
rect 31021 54275 31079 54281
rect 33686 54272 33692 54284
rect 33744 54272 33750 54324
rect 35250 54312 35256 54324
rect 35211 54284 35256 54312
rect 35250 54272 35256 54284
rect 35308 54272 35314 54324
rect 57241 54315 57299 54321
rect 57241 54281 57253 54315
rect 57287 54312 57299 54315
rect 57698 54312 57704 54324
rect 57287 54284 57704 54312
rect 57287 54281 57299 54284
rect 57241 54275 57299 54281
rect 57698 54272 57704 54284
rect 57756 54272 57762 54324
rect 1394 54108 1400 54120
rect 1355 54080 1400 54108
rect 1394 54068 1400 54080
rect 1452 54068 1458 54120
rect 22186 54068 22192 54120
rect 22244 54108 22250 54120
rect 22557 54111 22615 54117
rect 22557 54108 22569 54111
rect 22244 54080 22569 54108
rect 22244 54068 22250 54080
rect 22557 54077 22569 54080
rect 22603 54077 22615 54111
rect 22940 54108 22968 54272
rect 23308 54176 23336 54272
rect 23308 54148 23888 54176
rect 23201 54111 23259 54117
rect 23201 54108 23213 54111
rect 22940 54080 23213 54108
rect 22557 54071 22615 54077
rect 23201 54077 23213 54080
rect 23247 54077 23259 54111
rect 23382 54108 23388 54120
rect 23343 54080 23388 54108
rect 23201 54071 23259 54077
rect 23382 54068 23388 54080
rect 23440 54068 23446 54120
rect 23860 54117 23888 54148
rect 23845 54111 23903 54117
rect 23845 54077 23857 54111
rect 23891 54077 23903 54111
rect 23952 54108 23980 54272
rect 39574 54244 39580 54256
rect 33244 54216 39580 54244
rect 24302 54136 24308 54188
rect 24360 54176 24366 54188
rect 25869 54179 25927 54185
rect 24360 54148 24716 54176
rect 24360 54136 24366 54148
rect 24688 54117 24716 54148
rect 25869 54145 25881 54179
rect 25915 54176 25927 54179
rect 26789 54179 26847 54185
rect 26789 54176 26801 54179
rect 25915 54148 26801 54176
rect 25915 54145 25927 54148
rect 25869 54139 25927 54145
rect 26789 54145 26801 54148
rect 26835 54145 26847 54179
rect 26789 54139 26847 54145
rect 26881 54179 26939 54185
rect 26881 54145 26893 54179
rect 26927 54176 26939 54179
rect 27706 54176 27712 54188
rect 26927 54148 27712 54176
rect 26927 54145 26939 54148
rect 26881 54139 26939 54145
rect 24489 54111 24547 54117
rect 24489 54108 24501 54111
rect 23952 54080 24501 54108
rect 23845 54071 23903 54077
rect 24489 54077 24501 54080
rect 24535 54077 24547 54111
rect 24489 54071 24547 54077
rect 24673 54111 24731 54117
rect 24673 54077 24685 54111
rect 24719 54077 24731 54111
rect 24673 54071 24731 54077
rect 24762 54068 24768 54120
rect 24820 54108 24826 54120
rect 25133 54111 25191 54117
rect 25133 54108 25145 54111
rect 24820 54080 25145 54108
rect 24820 54068 24826 54080
rect 25133 54077 25145 54080
rect 25179 54077 25191 54111
rect 25133 54071 25191 54077
rect 25406 54068 25412 54120
rect 25464 54108 25470 54120
rect 25777 54111 25835 54117
rect 25777 54108 25789 54111
rect 25464 54080 25789 54108
rect 25464 54068 25470 54080
rect 25777 54077 25789 54080
rect 25823 54077 25835 54111
rect 25777 54071 25835 54077
rect 26605 54111 26663 54117
rect 26605 54077 26617 54111
rect 26651 54077 26663 54111
rect 26804 54108 26832 54139
rect 27706 54136 27712 54148
rect 27764 54176 27770 54188
rect 30469 54179 30527 54185
rect 27764 54148 28028 54176
rect 27764 54136 27770 54148
rect 28000 54117 28028 54148
rect 30469 54145 30481 54179
rect 30515 54176 30527 54179
rect 32125 54179 32183 54185
rect 32125 54176 32137 54179
rect 30515 54148 32137 54176
rect 30515 54145 30527 54148
rect 30469 54139 30527 54145
rect 32125 54145 32137 54148
rect 32171 54145 32183 54179
rect 32125 54139 32183 54145
rect 27801 54111 27859 54117
rect 27801 54108 27813 54111
rect 26804 54080 27813 54108
rect 26605 54071 26663 54077
rect 27801 54077 27813 54080
rect 27847 54077 27859 54111
rect 27801 54071 27859 54077
rect 27985 54111 28043 54117
rect 27985 54077 27997 54111
rect 28031 54077 28043 54111
rect 29178 54108 29184 54120
rect 29139 54080 29184 54108
rect 27985 54071 28043 54077
rect 26620 54040 26648 54071
rect 29178 54068 29184 54080
rect 29236 54068 29242 54120
rect 29362 54108 29368 54120
rect 29323 54080 29368 54108
rect 29362 54068 29368 54080
rect 29420 54068 29426 54120
rect 29546 54117 29552 54120
rect 29503 54111 29552 54117
rect 29503 54077 29515 54111
rect 29549 54077 29552 54111
rect 29503 54071 29552 54077
rect 29546 54068 29552 54071
rect 29604 54068 29610 54120
rect 29641 54111 29699 54117
rect 29641 54077 29653 54111
rect 29687 54108 29699 54111
rect 29914 54108 29920 54120
rect 29687 54080 29920 54108
rect 29687 54077 29699 54080
rect 29641 54071 29699 54077
rect 29914 54068 29920 54080
rect 29972 54068 29978 54120
rect 31478 54108 31484 54120
rect 31439 54080 31484 54108
rect 31478 54068 31484 54080
rect 31536 54068 31542 54120
rect 33042 54108 33048 54120
rect 33003 54080 33048 54108
rect 33042 54068 33048 54080
rect 33100 54068 33106 54120
rect 33244 54117 33272 54216
rect 39574 54204 39580 54216
rect 39632 54204 39638 54256
rect 58158 54244 58164 54256
rect 58119 54216 58164 54244
rect 58158 54204 58164 54216
rect 58216 54204 58222 54256
rect 35894 54176 35900 54188
rect 35807 54148 35900 54176
rect 35894 54136 35900 54148
rect 35952 54176 35958 54188
rect 36449 54179 36507 54185
rect 36449 54176 36461 54179
rect 35952 54148 36461 54176
rect 35952 54136 35958 54148
rect 36449 54145 36461 54148
rect 36495 54145 36507 54179
rect 36449 54139 36507 54145
rect 33229 54111 33287 54117
rect 33229 54077 33241 54111
rect 33275 54077 33287 54111
rect 33229 54071 33287 54077
rect 33321 54111 33379 54117
rect 33321 54077 33333 54111
rect 33367 54077 33379 54111
rect 33321 54071 33379 54077
rect 33413 54111 33471 54117
rect 33413 54077 33425 54111
rect 33459 54077 33471 54111
rect 33594 54108 33600 54120
rect 33555 54080 33600 54108
rect 33413 54071 33471 54077
rect 27890 54040 27896 54052
rect 26620 54012 27896 54040
rect 27890 54000 27896 54012
rect 27948 54000 27954 54052
rect 28902 54000 28908 54052
rect 28960 54040 28966 54052
rect 29273 54043 29331 54049
rect 29273 54040 29285 54043
rect 28960 54012 29285 54040
rect 28960 54000 28966 54012
rect 29273 54009 29285 54012
rect 29319 54009 29331 54043
rect 29273 54003 29331 54009
rect 32858 54000 32864 54052
rect 32916 54040 32922 54052
rect 33134 54040 33140 54052
rect 32916 54012 33140 54040
rect 32916 54000 32922 54012
rect 33134 54000 33140 54012
rect 33192 54040 33198 54052
rect 33336 54040 33364 54071
rect 33192 54012 33364 54040
rect 33428 54040 33456 54071
rect 33594 54068 33600 54080
rect 33652 54068 33658 54120
rect 35434 54108 35440 54120
rect 35395 54080 35440 54108
rect 35434 54068 35440 54080
rect 35492 54068 35498 54120
rect 35621 54111 35679 54117
rect 35621 54077 35633 54111
rect 35667 54108 35679 54111
rect 36170 54108 36176 54120
rect 35667 54080 36176 54108
rect 35667 54077 35679 54080
rect 35621 54071 35679 54077
rect 36170 54068 36176 54080
rect 36228 54108 36234 54120
rect 36228 54080 36308 54108
rect 36228 54068 36234 54080
rect 33502 54040 33508 54052
rect 33428 54012 33508 54040
rect 33192 54000 33198 54012
rect 8294 53932 8300 53984
rect 8352 53972 8358 53984
rect 8846 53972 8852 53984
rect 8352 53944 8852 53972
rect 8352 53932 8358 53944
rect 8846 53932 8852 53944
rect 8904 53932 8910 53984
rect 25225 53975 25283 53981
rect 25225 53941 25237 53975
rect 25271 53972 25283 53975
rect 25590 53972 25596 53984
rect 25271 53944 25596 53972
rect 25271 53941 25283 53944
rect 25225 53935 25283 53941
rect 25590 53932 25596 53944
rect 25648 53932 25654 53984
rect 26418 53972 26424 53984
rect 26379 53944 26424 53972
rect 26418 53932 26424 53944
rect 26476 53932 26482 53984
rect 32950 53932 32956 53984
rect 33008 53972 33014 53984
rect 33318 53972 33324 53984
rect 33008 53944 33324 53972
rect 33008 53932 33014 53944
rect 33318 53932 33324 53944
rect 33376 53972 33382 53984
rect 33428 53972 33456 54012
rect 33502 54000 33508 54012
rect 33560 54000 33566 54052
rect 35529 54043 35587 54049
rect 35529 54009 35541 54043
rect 35575 54009 35587 54043
rect 35529 54003 35587 54009
rect 35759 54043 35817 54049
rect 35759 54009 35771 54043
rect 35805 54040 35817 54043
rect 36078 54040 36084 54052
rect 35805 54012 36084 54040
rect 35805 54009 35817 54012
rect 35759 54003 35817 54009
rect 33778 53972 33784 53984
rect 33376 53944 33456 53972
rect 33739 53944 33784 53972
rect 33376 53932 33382 53944
rect 33778 53932 33784 53944
rect 33836 53932 33842 53984
rect 35544 53972 35572 54003
rect 36078 54000 36084 54012
rect 36136 54000 36142 54052
rect 36280 54040 36308 54080
rect 36354 54068 36360 54120
rect 36412 54108 36418 54120
rect 36541 54111 36599 54117
rect 36412 54080 36457 54108
rect 36412 54068 36418 54080
rect 36541 54077 36553 54111
rect 36587 54077 36599 54111
rect 36541 54071 36599 54077
rect 55585 54111 55643 54117
rect 55585 54077 55597 54111
rect 55631 54108 55643 54111
rect 55674 54108 55680 54120
rect 55631 54080 55680 54108
rect 55631 54077 55643 54080
rect 55585 54071 55643 54077
rect 36556 54040 36584 54071
rect 55674 54068 55680 54080
rect 55732 54068 55738 54120
rect 56781 54111 56839 54117
rect 56781 54077 56793 54111
rect 56827 54108 56839 54111
rect 57330 54108 57336 54120
rect 56827 54080 57336 54108
rect 56827 54077 56839 54080
rect 56781 54071 56839 54077
rect 57330 54068 57336 54080
rect 57388 54068 57394 54120
rect 57422 54068 57428 54120
rect 57480 54108 57486 54120
rect 57480 54080 57525 54108
rect 57480 54068 57486 54080
rect 57974 54040 57980 54052
rect 36280 54012 36584 54040
rect 57935 54012 57980 54040
rect 57974 54000 57980 54012
rect 58032 54000 58038 54052
rect 36354 53972 36360 53984
rect 35544 53944 36360 53972
rect 36354 53932 36360 53944
rect 36412 53932 36418 53984
rect 1104 53882 58880 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 50326 53882
rect 50378 53830 50390 53882
rect 50442 53830 50454 53882
rect 50506 53830 50518 53882
rect 50570 53830 58880 53882
rect 1104 53808 58880 53830
rect 27706 53768 27712 53780
rect 27667 53740 27712 53768
rect 27706 53728 27712 53740
rect 27764 53728 27770 53780
rect 29362 53728 29368 53780
rect 29420 53768 29426 53780
rect 29549 53771 29607 53777
rect 29549 53768 29561 53771
rect 29420 53740 29561 53768
rect 29420 53728 29426 53740
rect 29549 53737 29561 53740
rect 29595 53737 29607 53771
rect 29549 53731 29607 53737
rect 33594 53728 33600 53780
rect 33652 53768 33658 53780
rect 34517 53771 34575 53777
rect 34517 53768 34529 53771
rect 33652 53740 34529 53768
rect 33652 53728 33658 53740
rect 34517 53737 34529 53740
rect 34563 53737 34575 53771
rect 56962 53768 56968 53780
rect 56923 53740 56968 53768
rect 34517 53731 34575 53737
rect 56962 53728 56968 53740
rect 57020 53728 57026 53780
rect 57974 53728 57980 53780
rect 58032 53768 58038 53780
rect 58161 53771 58219 53777
rect 58161 53768 58173 53771
rect 58032 53740 58173 53768
rect 58032 53728 58038 53740
rect 58161 53737 58173 53740
rect 58207 53737 58219 53771
rect 58161 53731 58219 53737
rect 22094 53700 22100 53712
rect 21192 53672 22100 53700
rect 21192 53641 21220 53672
rect 22094 53660 22100 53672
rect 22152 53660 22158 53712
rect 26418 53660 26424 53712
rect 26476 53700 26482 53712
rect 26574 53703 26632 53709
rect 26574 53700 26586 53703
rect 26476 53672 26586 53700
rect 26476 53660 26482 53672
rect 26574 53669 26586 53672
rect 26620 53669 26632 53703
rect 26574 53663 26632 53669
rect 28436 53703 28494 53709
rect 28436 53669 28448 53703
rect 28482 53700 28494 53703
rect 28534 53700 28540 53712
rect 28482 53672 28540 53700
rect 28482 53669 28494 53672
rect 28436 53663 28494 53669
rect 28534 53660 28540 53672
rect 28592 53660 28598 53712
rect 30650 53660 30656 53712
rect 30708 53700 30714 53712
rect 30708 53672 31156 53700
rect 30708 53660 30714 53672
rect 21177 53635 21235 53641
rect 21177 53601 21189 53635
rect 21223 53601 21235 53635
rect 21177 53595 21235 53601
rect 21444 53635 21502 53641
rect 21444 53601 21456 53635
rect 21490 53632 21502 53635
rect 21726 53632 21732 53644
rect 21490 53604 21732 53632
rect 21490 53601 21502 53604
rect 21444 53595 21502 53601
rect 21726 53592 21732 53604
rect 21784 53592 21790 53644
rect 23566 53592 23572 53644
rect 23624 53632 23630 53644
rect 23661 53635 23719 53641
rect 23661 53632 23673 53635
rect 23624 53604 23673 53632
rect 23624 53592 23630 53604
rect 23661 53601 23673 53604
rect 23707 53632 23719 53635
rect 24762 53632 24768 53644
rect 23707 53604 24768 53632
rect 23707 53601 23719 53604
rect 23661 53595 23719 53601
rect 24762 53592 24768 53604
rect 24820 53592 24826 53644
rect 25406 53632 25412 53644
rect 25367 53604 25412 53632
rect 25406 53592 25412 53604
rect 25464 53592 25470 53644
rect 25590 53632 25596 53644
rect 25551 53604 25596 53632
rect 25590 53592 25596 53604
rect 25648 53592 25654 53644
rect 26142 53592 26148 53644
rect 26200 53632 26206 53644
rect 26326 53632 26332 53644
rect 26200 53604 26332 53632
rect 26200 53592 26206 53604
rect 26326 53592 26332 53604
rect 26384 53592 26390 53644
rect 28169 53635 28227 53641
rect 28169 53601 28181 53635
rect 28215 53632 28227 53635
rect 28994 53632 29000 53644
rect 28215 53604 29000 53632
rect 28215 53601 28227 53604
rect 28169 53595 28227 53601
rect 28994 53592 29000 53604
rect 29052 53632 29058 53644
rect 30926 53641 30932 53644
rect 29052 53604 30052 53632
rect 29052 53592 29058 53604
rect 30024 53576 30052 53604
rect 30920 53595 30932 53641
rect 30984 53632 30990 53644
rect 31128 53632 31156 53672
rect 31294 53660 31300 53712
rect 31352 53700 31358 53712
rect 33404 53703 33462 53709
rect 31352 53672 33364 53700
rect 31352 53660 31358 53672
rect 32493 53635 32551 53641
rect 32493 53632 32505 53635
rect 30984 53604 31020 53632
rect 31128 53604 32505 53632
rect 30926 53592 30932 53595
rect 30984 53592 30990 53604
rect 32493 53601 32505 53604
rect 32539 53601 32551 53635
rect 32493 53595 32551 53601
rect 33137 53635 33195 53641
rect 33137 53601 33149 53635
rect 33183 53632 33195 53635
rect 33226 53632 33232 53644
rect 33183 53604 33232 53632
rect 33183 53601 33195 53604
rect 33137 53595 33195 53601
rect 33226 53592 33232 53604
rect 33284 53592 33290 53644
rect 33336 53632 33364 53672
rect 33404 53669 33416 53703
rect 33450 53700 33462 53703
rect 33778 53700 33784 53712
rect 33450 53672 33784 53700
rect 33450 53669 33462 53672
rect 33404 53663 33462 53669
rect 33778 53660 33784 53672
rect 33836 53660 33842 53712
rect 56873 53703 56931 53709
rect 56873 53669 56885 53703
rect 56919 53700 56931 53703
rect 57790 53700 57796 53712
rect 56919 53672 57796 53700
rect 56919 53669 56931 53672
rect 56873 53663 56931 53669
rect 57790 53660 57796 53672
rect 57848 53660 57854 53712
rect 34606 53632 34612 53644
rect 33336 53604 34612 53632
rect 34606 53592 34612 53604
rect 34664 53592 34670 53644
rect 35894 53632 35900 53644
rect 35855 53604 35900 53632
rect 35894 53592 35900 53604
rect 35952 53592 35958 53644
rect 36170 53632 36176 53644
rect 36131 53604 36176 53632
rect 36170 53592 36176 53604
rect 36228 53592 36234 53644
rect 55585 53635 55643 53641
rect 55585 53601 55597 53635
rect 55631 53632 55643 53635
rect 56502 53632 56508 53644
rect 55631 53604 56508 53632
rect 55631 53601 55643 53604
rect 55585 53595 55643 53601
rect 56502 53592 56508 53604
rect 56560 53592 56566 53644
rect 57330 53592 57336 53644
rect 57388 53632 57394 53644
rect 57517 53635 57575 53641
rect 57517 53632 57529 53635
rect 57388 53604 57529 53632
rect 57388 53592 57394 53604
rect 57517 53601 57529 53604
rect 57563 53601 57575 53635
rect 57517 53595 57575 53601
rect 23934 53564 23940 53576
rect 23895 53536 23940 53564
rect 23934 53524 23940 53536
rect 23992 53524 23998 53576
rect 25685 53567 25743 53573
rect 25685 53533 25697 53567
rect 25731 53564 25743 53567
rect 26050 53564 26056 53576
rect 25731 53536 26056 53564
rect 25731 53533 25743 53536
rect 25685 53527 25743 53533
rect 26050 53524 26056 53536
rect 26108 53524 26114 53576
rect 30006 53524 30012 53576
rect 30064 53564 30070 53576
rect 30653 53567 30711 53573
rect 30653 53564 30665 53567
rect 30064 53536 30665 53564
rect 30064 53524 30070 53536
rect 30653 53533 30665 53536
rect 30699 53533 30711 53567
rect 57698 53564 57704 53576
rect 57659 53536 57704 53564
rect 30653 53527 30711 53533
rect 57698 53524 57704 53536
rect 57756 53524 57762 53576
rect 31754 53456 31760 53508
rect 31812 53496 31818 53508
rect 32585 53499 32643 53505
rect 32585 53496 32597 53499
rect 31812 53468 32597 53496
rect 31812 53456 31818 53468
rect 32585 53465 32597 53468
rect 32631 53465 32643 53499
rect 32585 53459 32643 53465
rect 22554 53428 22560 53440
rect 22515 53400 22560 53428
rect 22554 53388 22560 53400
rect 22612 53388 22618 53440
rect 23474 53428 23480 53440
rect 23435 53400 23480 53428
rect 23474 53388 23480 53400
rect 23532 53388 23538 53440
rect 23658 53388 23664 53440
rect 23716 53428 23722 53440
rect 23845 53431 23903 53437
rect 23845 53428 23857 53431
rect 23716 53400 23857 53428
rect 23716 53388 23722 53400
rect 23845 53397 23857 53400
rect 23891 53397 23903 53431
rect 25222 53428 25228 53440
rect 25183 53400 25228 53428
rect 23845 53391 23903 53397
rect 25222 53388 25228 53400
rect 25280 53388 25286 53440
rect 32030 53428 32036 53440
rect 31991 53400 32036 53428
rect 32030 53388 32036 53400
rect 32088 53388 32094 53440
rect 32214 53388 32220 53440
rect 32272 53428 32278 53440
rect 33870 53428 33876 53440
rect 32272 53400 33876 53428
rect 32272 53388 32278 53400
rect 33870 53388 33876 53400
rect 33928 53388 33934 53440
rect 35710 53428 35716 53440
rect 35671 53400 35716 53428
rect 35710 53388 35716 53400
rect 35768 53388 35774 53440
rect 36081 53431 36139 53437
rect 36081 53397 36093 53431
rect 36127 53428 36139 53431
rect 36354 53428 36360 53440
rect 36127 53400 36360 53428
rect 36127 53397 36139 53400
rect 36081 53391 36139 53397
rect 36354 53388 36360 53400
rect 36412 53428 36418 53440
rect 36722 53428 36728 53440
rect 36412 53400 36728 53428
rect 36412 53388 36418 53400
rect 36722 53388 36728 53400
rect 36780 53388 36786 53440
rect 1104 53338 58880 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 58880 53338
rect 1104 53264 58880 53286
rect 11882 53184 11888 53236
rect 11940 53224 11946 53236
rect 11940 53196 26924 53224
rect 11940 53184 11946 53196
rect 21545 53159 21603 53165
rect 21545 53125 21557 53159
rect 21591 53156 21603 53159
rect 22186 53156 22192 53168
rect 21591 53128 22192 53156
rect 21591 53125 21603 53128
rect 21545 53119 21603 53125
rect 22186 53116 22192 53128
rect 22244 53116 22250 53168
rect 26050 53156 26056 53168
rect 26011 53128 26056 53156
rect 26050 53116 26056 53128
rect 26108 53116 26114 53168
rect 26896 53156 26924 53196
rect 29178 53184 29184 53236
rect 29236 53224 29242 53236
rect 29273 53227 29331 53233
rect 29273 53224 29285 53227
rect 29236 53196 29285 53224
rect 29236 53184 29242 53196
rect 29273 53193 29285 53196
rect 29319 53193 29331 53227
rect 29914 53224 29920 53236
rect 29875 53196 29920 53224
rect 29273 53187 29331 53193
rect 29914 53184 29920 53196
rect 29972 53184 29978 53236
rect 30926 53184 30932 53236
rect 30984 53224 30990 53236
rect 31113 53227 31171 53233
rect 31113 53224 31125 53227
rect 30984 53196 31125 53224
rect 30984 53184 30990 53196
rect 31113 53193 31125 53196
rect 31159 53193 31171 53227
rect 31113 53187 31171 53193
rect 32033 53227 32091 53233
rect 32033 53193 32045 53227
rect 32079 53224 32091 53227
rect 34146 53224 34152 53236
rect 32079 53196 34152 53224
rect 32079 53193 32091 53196
rect 32033 53187 32091 53193
rect 34146 53184 34152 53196
rect 34204 53184 34210 53236
rect 36081 53227 36139 53233
rect 34716 53196 35940 53224
rect 33042 53156 33048 53168
rect 26896 53128 33048 53156
rect 33042 53116 33048 53128
rect 33100 53116 33106 53168
rect 34716 53156 34744 53196
rect 33172 53128 34744 53156
rect 35912 53156 35940 53196
rect 36081 53193 36093 53227
rect 36127 53224 36139 53227
rect 36170 53224 36176 53236
rect 36127 53196 36176 53224
rect 36127 53193 36139 53196
rect 36081 53187 36139 53193
rect 36170 53184 36176 53196
rect 36228 53184 36234 53236
rect 57241 53227 57299 53233
rect 57241 53193 57253 53227
rect 57287 53224 57299 53227
rect 57698 53224 57704 53236
rect 57287 53196 57704 53224
rect 57287 53193 57299 53196
rect 57241 53187 57299 53193
rect 57698 53184 57704 53196
rect 57756 53184 57762 53236
rect 40402 53156 40408 53168
rect 35912 53128 40408 53156
rect 22094 53048 22100 53100
rect 22152 53088 22158 53100
rect 22830 53088 22836 53100
rect 22152 53060 22836 53088
rect 22152 53048 22158 53060
rect 22830 53048 22836 53060
rect 22888 53048 22894 53100
rect 26068 53088 26096 53116
rect 26068 53060 26740 53088
rect 1394 53020 1400 53032
rect 1355 52992 1400 53020
rect 1394 52980 1400 52992
rect 1452 52980 1458 53032
rect 21450 53020 21456 53032
rect 21411 52992 21456 53020
rect 21450 52980 21456 52992
rect 21508 52980 21514 53032
rect 21637 53023 21695 53029
rect 21637 52989 21649 53023
rect 21683 53020 21695 53023
rect 22554 53020 22560 53032
rect 21683 52992 22560 53020
rect 21683 52989 21695 52992
rect 21637 52983 21695 52989
rect 22554 52980 22560 52992
rect 22612 52980 22618 53032
rect 23100 53023 23158 53029
rect 23100 52989 23112 53023
rect 23146 53020 23158 53023
rect 23474 53020 23480 53032
rect 23146 52992 23480 53020
rect 23146 52989 23158 52992
rect 23100 52983 23158 52989
rect 23474 52980 23480 52992
rect 23532 52980 23538 53032
rect 24673 53023 24731 53029
rect 24673 52989 24685 53023
rect 24719 52989 24731 53023
rect 24673 52983 24731 52989
rect 24940 53023 24998 53029
rect 24940 52989 24952 53023
rect 24986 53020 24998 53023
rect 25222 53020 25228 53032
rect 24986 52992 25228 53020
rect 24986 52989 24998 52992
rect 24940 52983 24998 52989
rect 24688 52952 24716 52983
rect 25222 52980 25228 52992
rect 25280 52980 25286 53032
rect 25682 52980 25688 53032
rect 25740 53020 25746 53032
rect 26712 53029 26740 53060
rect 29362 53048 29368 53100
rect 29420 53088 29426 53100
rect 30742 53088 30748 53100
rect 29420 53060 30052 53088
rect 29420 53048 29426 53060
rect 26513 53023 26571 53029
rect 26513 53020 26525 53023
rect 25740 52992 26525 53020
rect 25740 52980 25746 52992
rect 26513 52989 26525 52992
rect 26559 52989 26571 53023
rect 26513 52983 26571 52989
rect 26697 53023 26755 53029
rect 26697 52989 26709 53023
rect 26743 52989 26755 53023
rect 27890 53020 27896 53032
rect 27851 52992 27896 53020
rect 26697 52983 26755 52989
rect 27890 52980 27896 52992
rect 27948 52980 27954 53032
rect 29181 53023 29239 53029
rect 29181 52989 29193 53023
rect 29227 53020 29239 53023
rect 29546 53020 29552 53032
rect 29227 52992 29552 53020
rect 29227 52989 29239 52992
rect 29181 52983 29239 52989
rect 29546 52980 29552 52992
rect 29604 52980 29610 53032
rect 30024 53029 30052 53060
rect 30484 53060 30748 53088
rect 30484 53029 30512 53060
rect 30742 53048 30748 53060
rect 30800 53048 30806 53100
rect 32030 53088 32036 53100
rect 30852 53060 32036 53088
rect 30650 53029 30656 53032
rect 29825 53023 29883 53029
rect 29825 52989 29837 53023
rect 29871 52989 29883 53023
rect 29825 52983 29883 52989
rect 30009 53023 30067 53029
rect 30009 52989 30021 53023
rect 30055 52989 30067 53023
rect 30009 52983 30067 52989
rect 30469 53023 30527 53029
rect 30469 52989 30481 53023
rect 30515 52989 30527 53023
rect 30469 52983 30527 52989
rect 30617 53023 30656 53029
rect 30617 52989 30629 53023
rect 30617 52983 30656 52989
rect 25314 52952 25320 52964
rect 24688 52924 25320 52952
rect 25314 52912 25320 52924
rect 25372 52912 25378 52964
rect 25406 52912 25412 52964
rect 25464 52952 25470 52964
rect 26605 52955 26663 52961
rect 26605 52952 26617 52955
rect 25464 52924 26617 52952
rect 25464 52912 25470 52924
rect 26605 52921 26617 52924
rect 26651 52921 26663 52955
rect 26605 52915 26663 52921
rect 27985 52955 28043 52961
rect 27985 52921 27997 52955
rect 28031 52952 28043 52955
rect 28902 52952 28908 52964
rect 28031 52924 28908 52952
rect 28031 52921 28043 52924
rect 27985 52915 28043 52921
rect 28902 52912 28908 52924
rect 28960 52952 28966 52964
rect 29840 52952 29868 52983
rect 30650 52980 30656 52983
rect 30708 52980 30714 53032
rect 30852 53020 30880 53060
rect 32030 53048 32036 53060
rect 32088 53048 32094 53100
rect 30760 52992 30880 53020
rect 30975 53023 31033 53029
rect 30760 52961 30788 52992
rect 30975 52989 30987 53023
rect 31021 53020 31033 53023
rect 31662 53020 31668 53032
rect 31021 52992 31668 53020
rect 31021 52989 31033 52992
rect 30975 52983 31033 52989
rect 31662 52980 31668 52992
rect 31720 52980 31726 53032
rect 31757 53023 31815 53029
rect 31757 52989 31769 53023
rect 31803 52989 31815 53023
rect 31757 52983 31815 52989
rect 31849 53023 31907 53029
rect 31849 52989 31861 53023
rect 31895 53020 31907 53023
rect 31938 53020 31944 53032
rect 31895 52992 31944 53020
rect 31895 52989 31907 52992
rect 31849 52983 31907 52989
rect 28960 52924 29868 52952
rect 30745 52955 30803 52961
rect 28960 52912 28966 52924
rect 30745 52921 30757 52955
rect 30791 52921 30803 52955
rect 30745 52915 30803 52921
rect 30837 52955 30895 52961
rect 30837 52921 30849 52955
rect 30883 52952 30895 52955
rect 31294 52952 31300 52964
rect 30883 52924 31300 52952
rect 30883 52921 30895 52924
rect 30837 52915 30895 52921
rect 23106 52844 23112 52896
rect 23164 52884 23170 52896
rect 23934 52884 23940 52896
rect 23164 52856 23940 52884
rect 23164 52844 23170 52856
rect 23934 52844 23940 52856
rect 23992 52884 23998 52896
rect 24213 52887 24271 52893
rect 24213 52884 24225 52887
rect 23992 52856 24225 52884
rect 23992 52844 23998 52856
rect 24213 52853 24225 52856
rect 24259 52853 24271 52887
rect 24213 52847 24271 52853
rect 30650 52844 30656 52896
rect 30708 52884 30714 52896
rect 30760 52884 30788 52915
rect 31294 52912 31300 52924
rect 31352 52912 31358 52964
rect 31772 52952 31800 52983
rect 31938 52980 31944 52992
rect 31996 52980 32002 53032
rect 33042 53020 33048 53032
rect 33003 52992 33048 53020
rect 33042 52980 33048 52992
rect 33100 52980 33106 53032
rect 33172 53020 33200 53128
rect 40402 53116 40408 53128
rect 40460 53116 40466 53168
rect 33233 53023 33291 53029
rect 33233 53020 33245 53023
rect 33172 52992 33245 53020
rect 33233 52989 33245 52992
rect 33279 52989 33291 53023
rect 33233 52983 33291 52989
rect 33321 53023 33379 53029
rect 33321 52989 33333 53023
rect 33367 52989 33379 53023
rect 33321 52983 33379 52989
rect 33413 53023 33471 53029
rect 33413 52989 33425 53023
rect 33459 52989 33471 53023
rect 33413 52983 33471 52989
rect 32214 52952 32220 52964
rect 31772 52924 32220 52952
rect 32214 52912 32220 52924
rect 32272 52912 32278 52964
rect 33134 52912 33140 52964
rect 33192 52952 33198 52964
rect 33336 52952 33364 52983
rect 33192 52924 33364 52952
rect 33192 52912 33198 52924
rect 30708 52856 30788 52884
rect 30708 52844 30714 52856
rect 32122 52844 32128 52896
rect 32180 52884 32186 52896
rect 33318 52884 33324 52896
rect 32180 52856 33324 52884
rect 32180 52844 32186 52856
rect 33318 52844 33324 52856
rect 33376 52884 33382 52896
rect 33419 52884 33447 52983
rect 33502 52980 33508 53032
rect 33560 53020 33566 53032
rect 33597 53023 33655 53029
rect 33597 53020 33609 53023
rect 33560 52992 33609 53020
rect 33560 52980 33566 52992
rect 33597 52989 33609 52992
rect 33643 52989 33655 53023
rect 34698 53020 34704 53032
rect 34659 52992 34704 53020
rect 33597 52983 33655 52989
rect 34698 52980 34704 52992
rect 34756 52980 34762 53032
rect 34968 53023 35026 53029
rect 34968 52989 34980 53023
rect 35014 53020 35026 53023
rect 35710 53020 35716 53032
rect 35014 52992 35716 53020
rect 35014 52989 35026 52992
rect 34968 52983 35026 52989
rect 35710 52980 35716 52992
rect 35768 52980 35774 53032
rect 56502 52980 56508 53032
rect 56560 53020 56566 53032
rect 56597 53023 56655 53029
rect 56597 53020 56609 53023
rect 56560 52992 56609 53020
rect 56560 52980 56566 52992
rect 56597 52989 56609 52992
rect 56643 52989 56655 53023
rect 56597 52983 56655 52989
rect 57425 53023 57483 53029
rect 57425 52989 57437 53023
rect 57471 53020 57483 53023
rect 57514 53020 57520 53032
rect 57471 52992 57520 53020
rect 57471 52989 57483 52992
rect 57425 52983 57483 52989
rect 57514 52980 57520 52992
rect 57572 52980 57578 53032
rect 57974 52952 57980 52964
rect 57935 52924 57980 52952
rect 57974 52912 57980 52924
rect 58032 52912 58038 52964
rect 58158 52952 58164 52964
rect 58119 52924 58164 52952
rect 58158 52912 58164 52924
rect 58216 52912 58222 52964
rect 33778 52884 33784 52896
rect 33376 52856 33447 52884
rect 33739 52856 33784 52884
rect 33376 52844 33382 52856
rect 33778 52844 33784 52856
rect 33836 52844 33842 52896
rect 1104 52794 58880 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 50326 52794
rect 50378 52742 50390 52794
rect 50442 52742 50454 52794
rect 50506 52742 50518 52794
rect 50570 52742 58880 52794
rect 1104 52720 58880 52742
rect 21726 52680 21732 52692
rect 21687 52652 21732 52680
rect 21726 52640 21732 52652
rect 21784 52640 21790 52692
rect 22186 52680 22192 52692
rect 22066 52652 22192 52680
rect 22066 52612 22094 52652
rect 22186 52640 22192 52652
rect 22244 52640 22250 52692
rect 23109 52683 23167 52689
rect 23109 52649 23121 52683
rect 23155 52680 23167 52683
rect 23474 52680 23480 52692
rect 23155 52652 23480 52680
rect 23155 52649 23167 52652
rect 23109 52643 23167 52649
rect 23474 52640 23480 52652
rect 23532 52640 23538 52692
rect 23658 52680 23664 52692
rect 23619 52652 23664 52680
rect 23658 52640 23664 52652
rect 23716 52640 23722 52692
rect 31205 52683 31263 52689
rect 31205 52649 31217 52683
rect 31251 52680 31263 52683
rect 31478 52680 31484 52692
rect 31251 52652 31484 52680
rect 31251 52649 31263 52652
rect 31205 52643 31263 52649
rect 31478 52640 31484 52652
rect 31536 52640 31542 52692
rect 31665 52683 31723 52689
rect 31665 52649 31677 52683
rect 31711 52649 31723 52683
rect 33226 52680 33232 52692
rect 31665 52643 31723 52649
rect 33060 52652 33232 52680
rect 23676 52612 23704 52640
rect 21928 52584 22094 52612
rect 22940 52584 23704 52612
rect 28436 52615 28494 52621
rect 20898 52504 20904 52556
rect 20956 52544 20962 52556
rect 21928 52553 21956 52584
rect 21085 52547 21143 52553
rect 21085 52544 21097 52547
rect 20956 52516 21097 52544
rect 20956 52504 20962 52516
rect 21085 52513 21097 52516
rect 21131 52513 21143 52547
rect 21085 52507 21143 52513
rect 21913 52547 21971 52553
rect 21913 52513 21925 52547
rect 21959 52513 21971 52547
rect 21913 52507 21971 52513
rect 22189 52547 22247 52553
rect 22189 52513 22201 52547
rect 22235 52544 22247 52547
rect 22554 52544 22560 52556
rect 22235 52516 22560 52544
rect 22235 52513 22247 52516
rect 22189 52507 22247 52513
rect 22554 52504 22560 52516
rect 22612 52504 22618 52556
rect 22940 52553 22968 52584
rect 28436 52581 28448 52615
rect 28482 52612 28494 52615
rect 29086 52612 29092 52624
rect 28482 52584 29092 52612
rect 28482 52581 28494 52584
rect 28436 52575 28494 52581
rect 29086 52572 29092 52584
rect 29144 52572 29150 52624
rect 30374 52572 30380 52624
rect 30432 52612 30438 52624
rect 31680 52612 31708 52643
rect 30432 52584 31708 52612
rect 30432 52572 30438 52584
rect 22925 52547 22983 52553
rect 22925 52513 22937 52547
rect 22971 52513 22983 52547
rect 23106 52544 23112 52556
rect 23067 52516 23112 52544
rect 22925 52507 22983 52513
rect 23106 52504 23112 52516
rect 23164 52504 23170 52556
rect 23569 52547 23627 52553
rect 23569 52513 23581 52547
rect 23615 52544 23627 52547
rect 23750 52544 23756 52556
rect 23615 52516 23756 52544
rect 23615 52513 23627 52516
rect 23569 52507 23627 52513
rect 23750 52504 23756 52516
rect 23808 52504 23814 52556
rect 25685 52547 25743 52553
rect 25685 52513 25697 52547
rect 25731 52513 25743 52547
rect 25685 52507 25743 52513
rect 25869 52547 25927 52553
rect 25869 52513 25881 52547
rect 25915 52544 25927 52547
rect 26142 52544 26148 52556
rect 25915 52516 26148 52544
rect 25915 52513 25927 52516
rect 25869 52507 25927 52513
rect 21177 52479 21235 52485
rect 21177 52445 21189 52479
rect 21223 52476 21235 52479
rect 21450 52476 21456 52488
rect 21223 52448 21456 52476
rect 21223 52445 21235 52448
rect 21177 52439 21235 52445
rect 21450 52436 21456 52448
rect 21508 52476 21514 52488
rect 22097 52479 22155 52485
rect 22097 52476 22109 52479
rect 21508 52448 22109 52476
rect 21508 52436 21514 52448
rect 22097 52445 22109 52448
rect 22143 52445 22155 52479
rect 25700 52476 25728 52507
rect 26142 52504 26148 52516
rect 26200 52504 26206 52556
rect 28169 52547 28227 52553
rect 28169 52513 28181 52547
rect 28215 52544 28227 52547
rect 30006 52544 30012 52556
rect 28215 52516 30012 52544
rect 28215 52513 28227 52516
rect 28169 52507 28227 52513
rect 30006 52504 30012 52516
rect 30064 52504 30070 52556
rect 30650 52544 30656 52556
rect 30611 52516 30656 52544
rect 30650 52504 30656 52516
rect 30708 52504 30714 52556
rect 32030 52544 32036 52556
rect 31991 52516 32036 52544
rect 32030 52504 32036 52516
rect 32088 52504 32094 52556
rect 32125 52547 32183 52553
rect 32125 52513 32137 52547
rect 32171 52544 32183 52547
rect 32582 52544 32588 52556
rect 32171 52516 32588 52544
rect 32171 52513 32183 52516
rect 32125 52507 32183 52513
rect 32582 52504 32588 52516
rect 32640 52504 32646 52556
rect 32861 52547 32919 52553
rect 32861 52513 32873 52547
rect 32907 52544 32919 52547
rect 33060 52544 33088 52652
rect 33226 52640 33232 52652
rect 33284 52640 33290 52692
rect 36722 52680 36728 52692
rect 36683 52652 36728 52680
rect 36722 52640 36728 52652
rect 36780 52640 36786 52692
rect 57974 52640 57980 52692
rect 58032 52680 58038 52692
rect 58161 52683 58219 52689
rect 58161 52680 58173 52683
rect 58032 52652 58173 52680
rect 58032 52640 58038 52652
rect 58161 52649 58173 52652
rect 58207 52649 58219 52683
rect 58161 52643 58219 52649
rect 33128 52615 33186 52621
rect 33128 52581 33140 52615
rect 33174 52612 33186 52615
rect 33778 52612 33784 52624
rect 33174 52584 33784 52612
rect 33174 52581 33186 52584
rect 33128 52575 33186 52581
rect 33778 52572 33784 52584
rect 33836 52572 33842 52624
rect 34054 52544 34060 52556
rect 32907 52516 34060 52544
rect 32907 52513 32919 52516
rect 32861 52507 32919 52513
rect 34054 52504 34060 52516
rect 34112 52544 34118 52556
rect 34330 52544 34336 52556
rect 34112 52516 34336 52544
rect 34112 52504 34118 52516
rect 34330 52504 34336 52516
rect 34388 52504 34394 52556
rect 35897 52547 35955 52553
rect 35897 52513 35909 52547
rect 35943 52544 35955 52547
rect 36262 52544 36268 52556
rect 35943 52516 36268 52544
rect 35943 52513 35955 52516
rect 35897 52507 35955 52513
rect 36262 52504 36268 52516
rect 36320 52544 36326 52556
rect 36633 52547 36691 52553
rect 36633 52544 36645 52547
rect 36320 52516 36645 52544
rect 36320 52504 36326 52516
rect 36633 52513 36645 52516
rect 36679 52513 36691 52547
rect 36633 52507 36691 52513
rect 26234 52476 26240 52488
rect 25700 52448 26240 52476
rect 22097 52439 22155 52445
rect 26234 52436 26240 52448
rect 26292 52436 26298 52488
rect 32309 52479 32367 52485
rect 32309 52445 32321 52479
rect 32355 52445 32367 52479
rect 32309 52439 32367 52445
rect 25682 52340 25688 52352
rect 25643 52312 25688 52340
rect 25682 52300 25688 52312
rect 25740 52300 25746 52352
rect 29270 52300 29276 52352
rect 29328 52340 29334 52352
rect 29549 52343 29607 52349
rect 29549 52340 29561 52343
rect 29328 52312 29561 52340
rect 29328 52300 29334 52312
rect 29549 52309 29561 52312
rect 29595 52309 29607 52343
rect 32324 52340 32352 52439
rect 36078 52436 36084 52488
rect 36136 52476 36142 52488
rect 36173 52479 36231 52485
rect 36173 52476 36185 52479
rect 36136 52448 36185 52476
rect 36136 52436 36142 52448
rect 36173 52445 36185 52448
rect 36219 52445 36231 52479
rect 36173 52439 36231 52445
rect 57057 52479 57115 52485
rect 57057 52445 57069 52479
rect 57103 52476 57115 52479
rect 57517 52479 57575 52485
rect 57517 52476 57529 52479
rect 57103 52448 57529 52476
rect 57103 52445 57115 52448
rect 57057 52439 57115 52445
rect 57517 52445 57529 52448
rect 57563 52445 57575 52479
rect 57698 52476 57704 52488
rect 57659 52448 57704 52476
rect 57517 52439 57575 52445
rect 57698 52436 57704 52448
rect 57756 52436 57762 52488
rect 33502 52340 33508 52352
rect 32324 52312 33508 52340
rect 29549 52303 29607 52309
rect 33502 52300 33508 52312
rect 33560 52340 33566 52352
rect 34241 52343 34299 52349
rect 34241 52340 34253 52343
rect 33560 52312 34253 52340
rect 33560 52300 33566 52312
rect 34241 52309 34253 52312
rect 34287 52309 34299 52343
rect 35710 52340 35716 52352
rect 35671 52312 35716 52340
rect 34241 52303 34299 52309
rect 35710 52300 35716 52312
rect 35768 52300 35774 52352
rect 36081 52343 36139 52349
rect 36081 52309 36093 52343
rect 36127 52340 36139 52343
rect 36170 52340 36176 52352
rect 36127 52312 36176 52340
rect 36127 52309 36139 52312
rect 36081 52303 36139 52309
rect 36170 52300 36176 52312
rect 36228 52300 36234 52352
rect 1104 52250 58880 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 58880 52250
rect 1104 52176 58880 52198
rect 25958 52136 25964 52148
rect 25919 52108 25964 52136
rect 25958 52096 25964 52108
rect 26016 52096 26022 52148
rect 26326 52096 26332 52148
rect 26384 52136 26390 52148
rect 26605 52139 26663 52145
rect 26605 52136 26617 52139
rect 26384 52108 26617 52136
rect 26384 52096 26390 52108
rect 26605 52105 26617 52108
rect 26651 52105 26663 52139
rect 26605 52099 26663 52105
rect 32030 52096 32036 52148
rect 32088 52136 32094 52148
rect 33045 52139 33103 52145
rect 33045 52136 33057 52139
rect 32088 52108 33057 52136
rect 32088 52096 32094 52108
rect 33045 52105 33057 52108
rect 33091 52105 33103 52139
rect 36262 52136 36268 52148
rect 36223 52108 36268 52136
rect 33045 52099 33103 52105
rect 36262 52096 36268 52108
rect 36320 52096 36326 52148
rect 57241 52139 57299 52145
rect 57241 52105 57253 52139
rect 57287 52136 57299 52139
rect 57698 52136 57704 52148
rect 57287 52108 57704 52136
rect 57287 52105 57299 52108
rect 57241 52099 57299 52105
rect 57698 52096 57704 52108
rect 57756 52096 57762 52148
rect 32122 52068 32128 52080
rect 32083 52040 32128 52068
rect 32122 52028 32128 52040
rect 32180 52028 32186 52080
rect 58158 52068 58164 52080
rect 58119 52040 58164 52068
rect 58158 52028 58164 52040
rect 58216 52028 58222 52080
rect 21358 51960 21364 52012
rect 21416 52000 21422 52012
rect 21545 52003 21603 52009
rect 21545 52000 21557 52003
rect 21416 51972 21557 52000
rect 21416 51960 21422 51972
rect 21545 51969 21557 51972
rect 21591 51969 21603 52003
rect 21545 51963 21603 51969
rect 22830 51960 22836 52012
rect 22888 52000 22894 52012
rect 23937 52003 23995 52009
rect 23937 52000 23949 52003
rect 22888 51972 23949 52000
rect 22888 51960 22894 51972
rect 23937 51969 23949 51972
rect 23983 51969 23995 52003
rect 23937 51963 23995 51969
rect 28905 52003 28963 52009
rect 28905 51969 28917 52003
rect 28951 52000 28963 52003
rect 33594 52000 33600 52012
rect 28951 51972 30144 52000
rect 33555 51972 33600 52000
rect 28951 51969 28963 51972
rect 28905 51963 28963 51969
rect 1394 51932 1400 51944
rect 1355 51904 1400 51932
rect 1394 51892 1400 51904
rect 1452 51892 1458 51944
rect 20898 51892 20904 51944
rect 20956 51932 20962 51944
rect 21269 51935 21327 51941
rect 21269 51932 21281 51935
rect 20956 51904 21281 51932
rect 20956 51892 20962 51904
rect 21269 51901 21281 51904
rect 21315 51901 21327 51935
rect 21450 51932 21456 51944
rect 21411 51904 21456 51932
rect 21269 51895 21327 51901
rect 21450 51892 21456 51904
rect 21508 51892 21514 51944
rect 23109 51935 23167 51941
rect 23109 51901 23121 51935
rect 23155 51901 23167 51935
rect 23290 51932 23296 51944
rect 23251 51904 23296 51932
rect 23109 51895 23167 51901
rect 23124 51864 23152 51895
rect 23290 51892 23296 51904
rect 23348 51892 23354 51944
rect 23385 51935 23443 51941
rect 23385 51901 23397 51935
rect 23431 51932 23443 51935
rect 23658 51932 23664 51944
rect 23431 51904 23664 51932
rect 23431 51901 23443 51904
rect 23385 51895 23443 51901
rect 23658 51892 23664 51904
rect 23716 51892 23722 51944
rect 24026 51892 24032 51944
rect 24084 51932 24090 51944
rect 26789 51935 26847 51941
rect 26789 51932 26801 51935
rect 24084 51904 26801 51932
rect 24084 51892 24090 51904
rect 26789 51901 26801 51904
rect 26835 51901 26847 51935
rect 26789 51895 26847 51901
rect 27985 51935 28043 51941
rect 27985 51901 27997 51935
rect 28031 51901 28043 51935
rect 28166 51932 28172 51944
rect 28127 51904 28172 51932
rect 27985 51895 28043 51901
rect 23750 51864 23756 51876
rect 23124 51836 23756 51864
rect 23750 51824 23756 51836
rect 23808 51824 23814 51876
rect 24204 51867 24262 51873
rect 24204 51833 24216 51867
rect 24250 51864 24262 51867
rect 25038 51864 25044 51876
rect 24250 51836 25044 51864
rect 24250 51833 24262 51836
rect 24204 51827 24262 51833
rect 25038 51824 25044 51836
rect 25096 51824 25102 51876
rect 25777 51867 25835 51873
rect 25777 51833 25789 51867
rect 25823 51833 25835 51867
rect 28000 51864 28028 51895
rect 28166 51892 28172 51904
rect 28224 51892 28230 51944
rect 28261 51935 28319 51941
rect 28261 51901 28273 51935
rect 28307 51932 28319 51935
rect 28626 51932 28632 51944
rect 28307 51904 28632 51932
rect 28307 51901 28319 51904
rect 28261 51895 28319 51901
rect 28626 51892 28632 51904
rect 28684 51892 28690 51944
rect 29089 51935 29147 51941
rect 29089 51932 29101 51935
rect 29012 51904 29101 51932
rect 28810 51864 28816 51876
rect 28000 51836 28816 51864
rect 25777 51827 25835 51833
rect 21082 51796 21088 51808
rect 21043 51768 21088 51796
rect 21082 51756 21088 51768
rect 21140 51756 21146 51808
rect 22922 51796 22928 51808
rect 22883 51768 22928 51796
rect 22922 51756 22928 51768
rect 22980 51756 22986 51808
rect 25317 51799 25375 51805
rect 25317 51765 25329 51799
rect 25363 51796 25375 51799
rect 25590 51796 25596 51808
rect 25363 51768 25596 51796
rect 25363 51765 25375 51768
rect 25317 51759 25375 51765
rect 25590 51756 25596 51768
rect 25648 51796 25654 51808
rect 25792 51796 25820 51827
rect 28810 51824 28816 51836
rect 28868 51824 28874 51876
rect 25648 51768 25820 51796
rect 25648 51756 25654 51768
rect 25866 51756 25872 51808
rect 25924 51796 25930 51808
rect 25982 51799 26040 51805
rect 25982 51796 25994 51799
rect 25924 51768 25994 51796
rect 25924 51756 25930 51768
rect 25982 51765 25994 51768
rect 26028 51765 26040 51799
rect 26142 51796 26148 51808
rect 26103 51768 26148 51796
rect 25982 51759 26040 51765
rect 26142 51756 26148 51768
rect 26200 51756 26206 51808
rect 27798 51796 27804 51808
rect 27759 51768 27804 51796
rect 27798 51756 27804 51768
rect 27856 51756 27862 51808
rect 29012 51796 29040 51904
rect 29089 51901 29101 51904
rect 29135 51901 29147 51935
rect 29089 51895 29147 51901
rect 29549 51935 29607 51941
rect 29549 51901 29561 51935
rect 29595 51932 29607 51935
rect 29638 51932 29644 51944
rect 29595 51904 29644 51932
rect 29595 51901 29607 51904
rect 29549 51895 29607 51901
rect 29638 51892 29644 51904
rect 29696 51892 29702 51944
rect 30006 51932 30012 51944
rect 29967 51904 30012 51932
rect 30006 51892 30012 51904
rect 30064 51892 30070 51944
rect 30116 51932 30144 51972
rect 33594 51960 33600 51972
rect 33652 51960 33658 52012
rect 30265 51935 30323 51941
rect 30265 51932 30277 51935
rect 30116 51904 30277 51932
rect 30265 51901 30277 51904
rect 30311 51901 30323 51935
rect 30265 51895 30323 51901
rect 31754 51892 31760 51944
rect 31812 51932 31818 51944
rect 31941 51935 31999 51941
rect 31941 51932 31953 51935
rect 31812 51904 31953 51932
rect 31812 51892 31818 51904
rect 31941 51901 31953 51904
rect 31987 51901 31999 51935
rect 33410 51932 33416 51944
rect 33371 51904 33416 51932
rect 31941 51895 31999 51901
rect 33410 51892 33416 51904
rect 33468 51892 33474 51944
rect 34330 51932 34336 51944
rect 34291 51904 34336 51932
rect 34330 51892 34336 51904
rect 34388 51892 34394 51944
rect 34600 51935 34658 51941
rect 34600 51901 34612 51935
rect 34646 51932 34658 51935
rect 35710 51932 35716 51944
rect 34646 51904 35716 51932
rect 34646 51901 34658 51904
rect 34600 51895 34658 51901
rect 35710 51892 35716 51904
rect 35768 51892 35774 51944
rect 36170 51932 36176 51944
rect 36131 51904 36176 51932
rect 36170 51892 36176 51904
rect 36228 51892 36234 51944
rect 36357 51935 36415 51941
rect 36357 51901 36369 51935
rect 36403 51901 36415 51935
rect 36357 51895 36415 51901
rect 29178 51864 29184 51876
rect 29139 51836 29184 51864
rect 29178 51824 29184 51836
rect 29236 51824 29242 51876
rect 29270 51824 29276 51876
rect 29328 51864 29334 51876
rect 29411 51867 29469 51873
rect 29328 51836 29373 51864
rect 29328 51824 29334 51836
rect 29411 51833 29423 51867
rect 29457 51864 29469 51867
rect 32582 51864 32588 51876
rect 29457 51836 30236 51864
rect 29457 51833 29469 51836
rect 29411 51827 29469 51833
rect 29546 51796 29552 51808
rect 29012 51768 29552 51796
rect 29546 51756 29552 51768
rect 29604 51756 29610 51808
rect 30208 51796 30236 51836
rect 31726 51836 32588 51864
rect 31389 51799 31447 51805
rect 31389 51796 31401 51799
rect 30208 51768 31401 51796
rect 31389 51765 31401 51768
rect 31435 51796 31447 51799
rect 31726 51796 31754 51836
rect 32582 51824 32588 51836
rect 32640 51824 32646 51876
rect 36078 51864 36084 51876
rect 35728 51836 36084 51864
rect 31435 51768 31754 51796
rect 31435 51765 31447 51768
rect 31389 51759 31447 51765
rect 33502 51756 33508 51808
rect 33560 51796 33566 51808
rect 35728 51805 35756 51836
rect 36078 51824 36084 51836
rect 36136 51864 36142 51876
rect 36372 51864 36400 51895
rect 56502 51892 56508 51944
rect 56560 51932 56566 51944
rect 56597 51935 56655 51941
rect 56597 51932 56609 51935
rect 56560 51904 56609 51932
rect 56560 51892 56566 51904
rect 56597 51901 56609 51904
rect 56643 51901 56655 51935
rect 56597 51895 56655 51901
rect 57425 51935 57483 51941
rect 57425 51901 57437 51935
rect 57471 51932 57483 51935
rect 57514 51932 57520 51944
rect 57471 51904 57520 51932
rect 57471 51901 57483 51904
rect 57425 51895 57483 51901
rect 57514 51892 57520 51904
rect 57572 51892 57578 51944
rect 36136 51836 36400 51864
rect 57977 51867 58035 51873
rect 36136 51824 36142 51836
rect 57977 51833 57989 51867
rect 58023 51864 58035 51867
rect 58342 51864 58348 51876
rect 58023 51836 58348 51864
rect 58023 51833 58035 51836
rect 57977 51827 58035 51833
rect 58342 51824 58348 51836
rect 58400 51824 58406 51876
rect 35713 51799 35771 51805
rect 33560 51768 33605 51796
rect 33560 51756 33566 51768
rect 35713 51765 35725 51799
rect 35759 51765 35771 51799
rect 35713 51759 35771 51765
rect 1104 51706 58880 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 50326 51706
rect 50378 51654 50390 51706
rect 50442 51654 50454 51706
rect 50506 51654 50518 51706
rect 50570 51654 58880 51706
rect 1104 51632 58880 51654
rect 23658 51592 23664 51604
rect 23619 51564 23664 51592
rect 23658 51552 23664 51564
rect 23716 51552 23722 51604
rect 23750 51552 23756 51604
rect 23808 51592 23814 51604
rect 24213 51595 24271 51601
rect 24213 51592 24225 51595
rect 23808 51564 24225 51592
rect 23808 51552 23814 51564
rect 24213 51561 24225 51564
rect 24259 51561 24271 51595
rect 24213 51555 24271 51561
rect 25958 51552 25964 51604
rect 26016 51592 26022 51604
rect 26789 51595 26847 51601
rect 26789 51592 26801 51595
rect 26016 51564 26801 51592
rect 26016 51552 26022 51564
rect 26789 51561 26801 51564
rect 26835 51561 26847 51595
rect 28626 51592 28632 51604
rect 28587 51564 28632 51592
rect 26789 51555 26847 51561
rect 28626 51552 28632 51564
rect 28684 51592 28690 51604
rect 28994 51592 29000 51604
rect 28684 51564 29000 51592
rect 28684 51552 28690 51564
rect 28994 51552 29000 51564
rect 29052 51552 29058 51604
rect 29086 51552 29092 51604
rect 29144 51592 29150 51604
rect 31113 51595 31171 51601
rect 29144 51564 29189 51592
rect 29144 51552 29150 51564
rect 31113 51561 31125 51595
rect 31159 51592 31171 51595
rect 33134 51592 33140 51604
rect 31159 51564 33140 51592
rect 31159 51561 31171 51564
rect 31113 51555 31171 51561
rect 33134 51552 33140 51564
rect 33192 51552 33198 51604
rect 33413 51595 33471 51601
rect 33413 51561 33425 51595
rect 33459 51592 33471 51595
rect 33502 51592 33508 51604
rect 33459 51564 33508 51592
rect 33459 51561 33471 51564
rect 33413 51555 33471 51561
rect 33502 51552 33508 51564
rect 33560 51552 33566 51604
rect 20708 51527 20766 51533
rect 20708 51493 20720 51527
rect 20754 51524 20766 51527
rect 21082 51524 21088 51536
rect 20754 51496 21088 51524
rect 20754 51493 20766 51496
rect 20708 51487 20766 51493
rect 21082 51484 21088 51496
rect 21140 51484 21146 51536
rect 22548 51527 22606 51533
rect 22548 51493 22560 51527
rect 22594 51524 22606 51527
rect 22922 51524 22928 51536
rect 22594 51496 22928 51524
rect 22594 51493 22606 51496
rect 22548 51487 22606 51493
rect 22922 51484 22928 51496
rect 22980 51484 22986 51536
rect 23676 51524 23704 51552
rect 25682 51533 25688 51536
rect 25676 51524 25688 51533
rect 23676 51496 24348 51524
rect 25643 51496 25688 51524
rect 1394 51456 1400 51468
rect 1355 51428 1400 51456
rect 1394 51416 1400 51428
rect 1452 51416 1458 51468
rect 22278 51456 22284 51468
rect 22191 51428 22284 51456
rect 22278 51416 22284 51428
rect 22336 51456 22342 51468
rect 22830 51456 22836 51468
rect 22336 51428 22836 51456
rect 22336 51416 22342 51428
rect 22830 51416 22836 51428
rect 22888 51416 22894 51468
rect 23290 51416 23296 51468
rect 23348 51456 23354 51468
rect 24320 51465 24348 51496
rect 25676 51487 25688 51496
rect 25682 51484 25688 51487
rect 25740 51484 25746 51536
rect 27516 51527 27574 51533
rect 27516 51493 27528 51527
rect 27562 51524 27574 51527
rect 27798 51524 27804 51536
rect 27562 51496 27804 51524
rect 27562 51493 27574 51496
rect 27516 51487 27574 51493
rect 27798 51484 27804 51496
rect 27856 51484 27862 51536
rect 29546 51484 29552 51536
rect 29604 51524 29610 51536
rect 33965 51527 34023 51533
rect 33965 51524 33977 51527
rect 29604 51496 33977 51524
rect 29604 51484 29610 51496
rect 33965 51493 33977 51496
rect 34011 51493 34023 51527
rect 33965 51487 34023 51493
rect 24121 51459 24179 51465
rect 24121 51456 24133 51459
rect 23348 51428 24133 51456
rect 23348 51416 23354 51428
rect 24121 51425 24133 51428
rect 24167 51425 24179 51459
rect 24121 51419 24179 51425
rect 24305 51459 24363 51465
rect 24305 51425 24317 51459
rect 24351 51425 24363 51459
rect 26142 51456 26148 51468
rect 24305 51419 24363 51425
rect 25332 51428 26148 51456
rect 20438 51388 20444 51400
rect 20399 51360 20444 51388
rect 20438 51348 20444 51360
rect 20496 51348 20502 51400
rect 24136 51388 24164 51419
rect 25332 51388 25360 51428
rect 26142 51416 26148 51428
rect 26200 51416 26206 51468
rect 29273 51459 29331 51465
rect 29273 51425 29285 51459
rect 29319 51456 29331 51459
rect 29638 51456 29644 51468
rect 29319 51428 29644 51456
rect 29319 51425 29331 51428
rect 29273 51419 29331 51425
rect 29638 51416 29644 51428
rect 29696 51456 29702 51468
rect 30558 51456 30564 51468
rect 29696 51428 30564 51456
rect 29696 51416 29702 51428
rect 30558 51416 30564 51428
rect 30616 51416 30622 51468
rect 30834 51416 30840 51468
rect 30892 51456 30898 51468
rect 32306 51465 32312 51468
rect 31021 51459 31079 51465
rect 31021 51456 31033 51459
rect 30892 51428 31033 51456
rect 30892 51416 30898 51428
rect 31021 51425 31033 51428
rect 31067 51425 31079 51459
rect 31021 51419 31079 51425
rect 32300 51419 32312 51465
rect 32364 51456 32370 51468
rect 32364 51428 32400 51456
rect 32306 51416 32312 51419
rect 32364 51416 32370 51428
rect 32582 51416 32588 51468
rect 32640 51456 32646 51468
rect 33873 51459 33931 51465
rect 33873 51456 33885 51459
rect 32640 51428 33885 51456
rect 32640 51416 32646 51428
rect 33873 51425 33885 51428
rect 33919 51425 33931 51459
rect 57974 51456 57980 51468
rect 57935 51428 57980 51456
rect 33873 51419 33931 51425
rect 57974 51416 57980 51428
rect 58032 51416 58038 51468
rect 24136 51360 25360 51388
rect 25409 51391 25467 51397
rect 25409 51357 25421 51391
rect 25455 51357 25467 51391
rect 25409 51351 25467 51357
rect 27249 51391 27307 51397
rect 27249 51357 27261 51391
rect 27295 51357 27307 51391
rect 27249 51351 27307 51357
rect 21358 51212 21364 51264
rect 21416 51252 21422 51264
rect 21821 51255 21879 51261
rect 21821 51252 21833 51255
rect 21416 51224 21833 51252
rect 21416 51212 21422 51224
rect 21821 51221 21833 51224
rect 21867 51221 21879 51255
rect 25424 51252 25452 51351
rect 27264 51320 27292 51351
rect 29362 51348 29368 51400
rect 29420 51388 29426 51400
rect 29549 51391 29607 51397
rect 29549 51388 29561 51391
rect 29420 51360 29561 51388
rect 29420 51348 29426 51360
rect 29549 51357 29561 51360
rect 29595 51388 29607 51391
rect 30650 51388 30656 51400
rect 29595 51360 30656 51388
rect 29595 51357 29607 51360
rect 29549 51351 29607 51357
rect 30650 51348 30656 51360
rect 30708 51348 30714 51400
rect 31938 51348 31944 51400
rect 31996 51388 32002 51400
rect 32033 51391 32091 51397
rect 32033 51388 32045 51391
rect 31996 51360 32045 51388
rect 31996 51348 32002 51360
rect 32033 51357 32045 51360
rect 32079 51357 32091 51391
rect 32033 51351 32091 51357
rect 58158 51320 58164 51332
rect 26344 51292 27292 51320
rect 58119 51292 58164 51320
rect 26344 51264 26372 51292
rect 58158 51280 58164 51292
rect 58216 51280 58222 51332
rect 26326 51252 26332 51264
rect 25424 51224 26332 51252
rect 21821 51215 21879 51221
rect 26326 51212 26332 51224
rect 26384 51212 26390 51264
rect 29178 51212 29184 51264
rect 29236 51252 29242 51264
rect 29457 51255 29515 51261
rect 29457 51252 29469 51255
rect 29236 51224 29469 51252
rect 29236 51212 29242 51224
rect 29457 51221 29469 51224
rect 29503 51221 29515 51255
rect 57422 51252 57428 51264
rect 57383 51224 57428 51252
rect 29457 51215 29515 51221
rect 57422 51212 57428 51224
rect 57480 51212 57486 51264
rect 1104 51162 58880 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 58880 51162
rect 1104 51088 58880 51110
rect 20898 51048 20904 51060
rect 20859 51020 20904 51048
rect 20898 51008 20904 51020
rect 20956 51008 20962 51060
rect 21450 51008 21456 51060
rect 21508 51048 21514 51060
rect 21545 51051 21603 51057
rect 21545 51048 21557 51051
rect 21508 51020 21557 51048
rect 21508 51008 21514 51020
rect 21545 51017 21557 51020
rect 21591 51017 21603 51051
rect 25038 51048 25044 51060
rect 24999 51020 25044 51048
rect 21545 51011 21603 51017
rect 25038 51008 25044 51020
rect 25096 51008 25102 51060
rect 26145 51051 26203 51057
rect 26145 51017 26157 51051
rect 26191 51048 26203 51051
rect 26234 51048 26240 51060
rect 26191 51020 26240 51048
rect 26191 51017 26203 51020
rect 26145 51011 26203 51017
rect 26234 51008 26240 51020
rect 26292 51008 26298 51060
rect 28166 51008 28172 51060
rect 28224 51048 28230 51060
rect 28261 51051 28319 51057
rect 28261 51048 28273 51051
rect 28224 51020 28273 51048
rect 28224 51008 28230 51020
rect 28261 51017 28273 51020
rect 28307 51017 28319 51051
rect 28261 51011 28319 51017
rect 21468 50912 21496 51008
rect 20824 50884 21496 50912
rect 25593 50915 25651 50921
rect 20824 50853 20852 50884
rect 25593 50881 25605 50915
rect 25639 50912 25651 50915
rect 25866 50912 25872 50924
rect 25639 50884 25872 50912
rect 25639 50881 25651 50884
rect 25593 50875 25651 50881
rect 25866 50872 25872 50884
rect 25924 50872 25930 50924
rect 20809 50847 20867 50853
rect 20809 50813 20821 50847
rect 20855 50813 20867 50847
rect 20809 50807 20867 50813
rect 20993 50847 21051 50853
rect 20993 50813 21005 50847
rect 21039 50844 21051 50847
rect 21358 50844 21364 50856
rect 21039 50816 21364 50844
rect 21039 50813 21051 50816
rect 20993 50807 21051 50813
rect 21358 50804 21364 50816
rect 21416 50804 21422 50856
rect 21453 50847 21511 50853
rect 21453 50813 21465 50847
rect 21499 50844 21511 50847
rect 21634 50844 21640 50856
rect 21499 50816 21640 50844
rect 21499 50813 21511 50816
rect 21453 50807 21511 50813
rect 21634 50804 21640 50816
rect 21692 50804 21698 50856
rect 22833 50847 22891 50853
rect 22833 50813 22845 50847
rect 22879 50844 22891 50847
rect 24026 50844 24032 50856
rect 22879 50816 24032 50844
rect 22879 50813 22891 50816
rect 22833 50807 22891 50813
rect 24026 50804 24032 50816
rect 24084 50804 24090 50856
rect 25222 50847 25280 50853
rect 25222 50813 25234 50847
rect 25268 50844 25280 50847
rect 25498 50844 25504 50856
rect 25268 50816 25504 50844
rect 25268 50813 25280 50816
rect 25222 50807 25280 50813
rect 25498 50804 25504 50816
rect 25556 50804 25562 50856
rect 25685 50847 25743 50853
rect 25685 50813 25697 50847
rect 25731 50813 25743 50847
rect 25685 50807 25743 50813
rect 25516 50776 25544 50804
rect 25700 50776 25728 50807
rect 25958 50804 25964 50856
rect 26016 50844 26022 50856
rect 26145 50847 26203 50853
rect 26145 50844 26157 50847
rect 26016 50816 26157 50844
rect 26016 50804 26022 50816
rect 26145 50813 26157 50816
rect 26191 50813 26203 50847
rect 26145 50807 26203 50813
rect 26421 50847 26479 50853
rect 26421 50813 26433 50847
rect 26467 50844 26479 50847
rect 26694 50844 26700 50856
rect 26467 50816 26700 50844
rect 26467 50813 26479 50816
rect 26421 50807 26479 50813
rect 26694 50804 26700 50816
rect 26752 50804 26758 50856
rect 28166 50844 28172 50856
rect 28127 50816 28172 50844
rect 28166 50804 28172 50816
rect 28224 50804 28230 50856
rect 28276 50844 28304 51011
rect 28810 51008 28816 51060
rect 28868 51048 28874 51060
rect 28905 51051 28963 51057
rect 28905 51048 28917 51051
rect 28868 51020 28917 51048
rect 28868 51008 28874 51020
rect 28905 51017 28917 51020
rect 28951 51017 28963 51051
rect 28905 51011 28963 51017
rect 28920 50912 28948 51011
rect 29178 51008 29184 51060
rect 29236 51048 29242 51060
rect 29549 51051 29607 51057
rect 29549 51048 29561 51051
rect 29236 51020 29561 51048
rect 29236 51008 29242 51020
rect 29549 51017 29561 51020
rect 29595 51017 29607 51051
rect 30558 51048 30564 51060
rect 30519 51020 30564 51048
rect 29549 51011 29607 51017
rect 28920 50884 29500 50912
rect 28813 50847 28871 50853
rect 28813 50844 28825 50847
rect 28276 50816 28825 50844
rect 28813 50813 28825 50816
rect 28859 50813 28871 50847
rect 28994 50844 29000 50856
rect 28955 50816 29000 50844
rect 28813 50807 28871 50813
rect 28994 50804 29000 50816
rect 29052 50804 29058 50856
rect 29472 50853 29500 50884
rect 29457 50847 29515 50853
rect 29457 50813 29469 50847
rect 29503 50813 29515 50847
rect 29564 50844 29592 51011
rect 30558 51008 30564 51020
rect 30616 51008 30622 51060
rect 35805 51051 35863 51057
rect 35805 51017 35817 51051
rect 35851 51048 35863 51051
rect 36170 51048 36176 51060
rect 35851 51020 36176 51048
rect 35851 51017 35863 51020
rect 35805 51011 35863 51017
rect 36170 51008 36176 51020
rect 36228 51008 36234 51060
rect 57974 51048 57980 51060
rect 57935 51020 57980 51048
rect 57974 51008 57980 51020
rect 58032 51008 58038 51060
rect 56873 50983 56931 50989
rect 56873 50949 56885 50983
rect 56919 50980 56931 50983
rect 56919 50952 57744 50980
rect 56919 50949 56931 50952
rect 56873 50943 56931 50949
rect 31478 50872 31484 50924
rect 31536 50912 31542 50924
rect 31757 50915 31815 50921
rect 31536 50884 31708 50912
rect 31536 50872 31542 50884
rect 30469 50847 30527 50853
rect 30469 50844 30481 50847
rect 29564 50816 30481 50844
rect 29457 50807 29515 50813
rect 30469 50813 30481 50816
rect 30515 50813 30527 50847
rect 30650 50844 30656 50856
rect 30611 50816 30656 50844
rect 30469 50807 30527 50813
rect 30650 50804 30656 50816
rect 30708 50804 30714 50856
rect 31573 50847 31631 50853
rect 31573 50813 31585 50847
rect 31619 50813 31631 50847
rect 31680 50844 31708 50884
rect 31757 50881 31769 50915
rect 31803 50912 31815 50915
rect 34609 50915 34667 50921
rect 31803 50884 33088 50912
rect 31803 50881 31815 50884
rect 31757 50875 31815 50881
rect 31772 50844 31800 50875
rect 31680 50816 31800 50844
rect 31573 50807 31631 50813
rect 26329 50779 26387 50785
rect 26329 50776 26341 50779
rect 25516 50748 26341 50776
rect 26329 50745 26341 50748
rect 26375 50745 26387 50779
rect 31588 50776 31616 50807
rect 31846 50804 31852 50856
rect 31904 50844 31910 50856
rect 33060 50853 33088 50884
rect 34609 50881 34621 50915
rect 34655 50912 34667 50915
rect 34790 50912 34796 50924
rect 34655 50884 34796 50912
rect 34655 50881 34667 50884
rect 34609 50875 34667 50881
rect 34790 50872 34796 50884
rect 34848 50912 34854 50924
rect 34848 50884 35296 50912
rect 34848 50872 34854 50884
rect 33045 50847 33103 50853
rect 31904 50816 31949 50844
rect 31904 50804 31910 50816
rect 33045 50813 33057 50847
rect 33091 50813 33103 50847
rect 33226 50844 33232 50856
rect 33187 50816 33232 50844
rect 33045 50807 33103 50813
rect 33226 50804 33232 50816
rect 33284 50804 33290 50856
rect 34333 50847 34391 50853
rect 34333 50813 34345 50847
rect 34379 50813 34391 50847
rect 34333 50807 34391 50813
rect 34517 50847 34575 50853
rect 34517 50813 34529 50847
rect 34563 50844 34575 50847
rect 34698 50844 34704 50856
rect 34563 50816 34704 50844
rect 34563 50813 34575 50816
rect 34517 50807 34575 50813
rect 32950 50776 32956 50788
rect 31588 50748 32956 50776
rect 26329 50739 26387 50745
rect 32950 50736 32956 50748
rect 33008 50776 33014 50788
rect 33137 50779 33195 50785
rect 33137 50776 33149 50779
rect 33008 50748 33149 50776
rect 33008 50736 33014 50748
rect 33137 50745 33149 50748
rect 33183 50745 33195 50779
rect 34348 50776 34376 50807
rect 34698 50804 34704 50816
rect 34756 50844 34762 50856
rect 35268 50853 35296 50884
rect 57422 50872 57428 50924
rect 57480 50912 57486 50924
rect 57716 50921 57744 50952
rect 57517 50915 57575 50921
rect 57517 50912 57529 50915
rect 57480 50884 57529 50912
rect 57480 50872 57486 50884
rect 57517 50881 57529 50884
rect 57563 50881 57575 50915
rect 57517 50875 57575 50881
rect 57701 50915 57759 50921
rect 57701 50881 57713 50915
rect 57747 50881 57759 50915
rect 57701 50875 57759 50881
rect 35069 50847 35127 50853
rect 35069 50844 35081 50847
rect 34756 50816 35081 50844
rect 34756 50804 34762 50816
rect 35069 50813 35081 50816
rect 35115 50813 35127 50847
rect 35069 50807 35127 50813
rect 35253 50847 35311 50853
rect 35253 50813 35265 50847
rect 35299 50813 35311 50847
rect 35253 50807 35311 50813
rect 35713 50847 35771 50853
rect 35713 50813 35725 50847
rect 35759 50813 35771 50847
rect 35713 50807 35771 50813
rect 57057 50847 57115 50853
rect 57057 50813 57069 50847
rect 57103 50844 57115 50847
rect 57103 50816 57560 50844
rect 57103 50813 57115 50816
rect 57057 50807 57115 50813
rect 35161 50779 35219 50785
rect 35161 50776 35173 50779
rect 34348 50748 35173 50776
rect 33137 50739 33195 50745
rect 35161 50745 35173 50748
rect 35207 50776 35219 50779
rect 35728 50776 35756 50807
rect 57532 50788 57560 50816
rect 35207 50748 35756 50776
rect 35207 50745 35219 50748
rect 35161 50739 35219 50745
rect 57514 50736 57520 50788
rect 57572 50736 57578 50788
rect 22278 50668 22284 50720
rect 22336 50708 22342 50720
rect 22646 50708 22652 50720
rect 22336 50680 22652 50708
rect 22336 50668 22342 50680
rect 22646 50668 22652 50680
rect 22704 50668 22710 50720
rect 25225 50711 25283 50717
rect 25225 50677 25237 50711
rect 25271 50708 25283 50711
rect 25866 50708 25872 50720
rect 25271 50680 25872 50708
rect 25271 50677 25283 50680
rect 25225 50671 25283 50677
rect 25866 50668 25872 50680
rect 25924 50668 25930 50720
rect 31386 50708 31392 50720
rect 31347 50680 31392 50708
rect 31386 50668 31392 50680
rect 31444 50668 31450 50720
rect 34146 50708 34152 50720
rect 34107 50680 34152 50708
rect 34146 50668 34152 50680
rect 34204 50668 34210 50720
rect 1104 50618 58880 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 50326 50618
rect 50378 50566 50390 50618
rect 50442 50566 50454 50618
rect 50506 50566 50518 50618
rect 50570 50566 58880 50618
rect 1104 50544 58880 50566
rect 23937 50507 23995 50513
rect 23937 50473 23949 50507
rect 23983 50504 23995 50507
rect 24026 50504 24032 50516
rect 23983 50476 24032 50504
rect 23983 50473 23995 50476
rect 23937 50467 23995 50473
rect 24026 50464 24032 50476
rect 24084 50464 24090 50516
rect 31846 50504 31852 50516
rect 31759 50476 31852 50504
rect 31846 50464 31852 50476
rect 31904 50464 31910 50516
rect 32306 50504 32312 50516
rect 32267 50476 32312 50504
rect 32306 50464 32312 50476
rect 32364 50464 32370 50516
rect 33226 50504 33232 50516
rect 32692 50476 33232 50504
rect 28166 50436 28172 50448
rect 28079 50408 28172 50436
rect 1394 50368 1400 50380
rect 1355 50340 1400 50368
rect 1394 50328 1400 50340
rect 1452 50328 1458 50380
rect 20349 50371 20407 50377
rect 20349 50337 20361 50371
rect 20395 50368 20407 50371
rect 21266 50368 21272 50380
rect 20395 50340 21272 50368
rect 20395 50337 20407 50340
rect 20349 50331 20407 50337
rect 21266 50328 21272 50340
rect 21324 50328 21330 50380
rect 21450 50377 21456 50380
rect 21444 50331 21456 50377
rect 21508 50368 21514 50380
rect 21508 50340 21544 50368
rect 21450 50328 21456 50331
rect 21508 50328 21514 50340
rect 23474 50328 23480 50380
rect 23532 50368 23538 50380
rect 24121 50371 24179 50377
rect 24121 50368 24133 50371
rect 23532 50340 24133 50368
rect 23532 50328 23538 50340
rect 24121 50337 24133 50340
rect 24167 50337 24179 50371
rect 24121 50331 24179 50337
rect 25498 50328 25504 50380
rect 25556 50368 25562 50380
rect 25777 50371 25835 50377
rect 25777 50368 25789 50371
rect 25556 50340 25789 50368
rect 25556 50328 25562 50340
rect 25777 50337 25789 50340
rect 25823 50337 25835 50371
rect 25777 50331 25835 50337
rect 25866 50328 25872 50380
rect 25924 50368 25930 50380
rect 25961 50371 26019 50377
rect 25961 50368 25973 50371
rect 25924 50340 25973 50368
rect 25924 50328 25930 50340
rect 25961 50337 25973 50340
rect 26007 50368 26019 50371
rect 26694 50368 26700 50380
rect 26007 50340 26700 50368
rect 26007 50337 26019 50340
rect 25961 50331 26019 50337
rect 26694 50328 26700 50340
rect 26752 50328 26758 50380
rect 28092 50377 28120 50408
rect 28166 50396 28172 50408
rect 28224 50436 28230 50448
rect 28905 50439 28963 50445
rect 28905 50436 28917 50439
rect 28224 50408 28917 50436
rect 28224 50396 28230 50408
rect 28905 50405 28917 50408
rect 28951 50405 28963 50439
rect 28905 50399 28963 50405
rect 30736 50439 30794 50445
rect 30736 50405 30748 50439
rect 30782 50436 30794 50439
rect 31386 50436 31392 50448
rect 30782 50408 31392 50436
rect 30782 50405 30794 50408
rect 30736 50399 30794 50405
rect 31386 50396 31392 50408
rect 31444 50396 31450 50448
rect 31864 50436 31892 50464
rect 32692 50445 32720 50476
rect 33226 50464 33232 50476
rect 33284 50464 33290 50516
rect 34790 50504 34796 50516
rect 34751 50476 34796 50504
rect 34790 50464 34796 50476
rect 34848 50464 34854 50516
rect 32677 50439 32735 50445
rect 32677 50436 32689 50439
rect 31864 50408 32689 50436
rect 32677 50405 32689 50408
rect 32723 50405 32735 50439
rect 32677 50399 32735 50405
rect 32815 50439 32873 50445
rect 32815 50405 32827 50439
rect 32861 50436 32873 50439
rect 33502 50436 33508 50448
rect 32861 50408 33508 50436
rect 32861 50405 32873 50408
rect 32815 50399 32873 50405
rect 33502 50396 33508 50408
rect 33560 50396 33566 50448
rect 33680 50439 33738 50445
rect 33680 50405 33692 50439
rect 33726 50436 33738 50439
rect 34146 50436 34152 50448
rect 33726 50408 34152 50436
rect 33726 50405 33738 50408
rect 33680 50399 33738 50405
rect 34146 50396 34152 50408
rect 34204 50396 34210 50448
rect 58158 50436 58164 50448
rect 58119 50408 58164 50436
rect 58158 50396 58164 50408
rect 58216 50396 58222 50448
rect 28077 50371 28135 50377
rect 28077 50337 28089 50371
rect 28123 50337 28135 50371
rect 28813 50371 28871 50377
rect 28813 50368 28825 50371
rect 28077 50331 28135 50337
rect 28276 50340 28825 50368
rect 20625 50303 20683 50309
rect 20625 50269 20637 50303
rect 20671 50300 20683 50303
rect 20806 50300 20812 50312
rect 20671 50272 20812 50300
rect 20671 50269 20683 50272
rect 20625 50263 20683 50269
rect 20806 50260 20812 50272
rect 20864 50260 20870 50312
rect 21177 50303 21235 50309
rect 21177 50269 21189 50303
rect 21223 50269 21235 50303
rect 21177 50263 21235 50269
rect 19426 50192 19432 50244
rect 19484 50232 19490 50244
rect 20438 50232 20444 50244
rect 19484 50204 20444 50232
rect 19484 50192 19490 50204
rect 20438 50192 20444 50204
rect 20496 50232 20502 50244
rect 21192 50232 21220 50263
rect 22646 50232 22652 50244
rect 20496 50204 21220 50232
rect 20496 50192 20502 50204
rect 20162 50164 20168 50176
rect 20123 50136 20168 50164
rect 20162 50124 20168 50136
rect 20220 50124 20226 50176
rect 20530 50164 20536 50176
rect 20491 50136 20536 50164
rect 20530 50124 20536 50136
rect 20588 50124 20594 50176
rect 21192 50164 21220 50204
rect 22480 50204 22652 50232
rect 22480 50164 22508 50204
rect 22646 50192 22652 50204
rect 22704 50192 22710 50244
rect 21192 50136 22508 50164
rect 22554 50124 22560 50176
rect 22612 50164 22618 50176
rect 25774 50164 25780 50176
rect 22612 50136 22657 50164
rect 25735 50136 25780 50164
rect 22612 50124 22618 50136
rect 25774 50124 25780 50136
rect 25832 50124 25838 50176
rect 27890 50164 27896 50176
rect 27851 50136 27896 50164
rect 27890 50124 27896 50136
rect 27948 50124 27954 50176
rect 28276 50173 28304 50340
rect 28813 50337 28825 50340
rect 28859 50337 28871 50371
rect 28994 50368 29000 50380
rect 28955 50340 29000 50368
rect 28813 50331 28871 50337
rect 28994 50328 29000 50340
rect 29052 50328 29058 50380
rect 30006 50328 30012 50380
rect 30064 50368 30070 50380
rect 30469 50371 30527 50377
rect 30469 50368 30481 50371
rect 30064 50340 30481 50368
rect 30064 50328 30070 50340
rect 30469 50337 30481 50340
rect 30515 50368 30527 50371
rect 31938 50368 31944 50380
rect 30515 50340 31944 50368
rect 30515 50337 30527 50340
rect 30469 50331 30527 50337
rect 31938 50328 31944 50340
rect 31996 50328 32002 50380
rect 32490 50368 32496 50380
rect 32451 50340 32496 50368
rect 32490 50328 32496 50340
rect 32548 50328 32554 50380
rect 32585 50371 32643 50377
rect 32585 50337 32597 50371
rect 32631 50337 32643 50371
rect 32950 50368 32956 50380
rect 32911 50340 32956 50368
rect 32585 50331 32643 50337
rect 28353 50303 28411 50309
rect 28353 50269 28365 50303
rect 28399 50300 28411 50303
rect 29012 50300 29040 50328
rect 28399 50272 29040 50300
rect 28399 50269 28411 50272
rect 28353 50263 28411 50269
rect 31478 50260 31484 50312
rect 31536 50300 31542 50312
rect 32600 50300 32628 50331
rect 32950 50328 32956 50340
rect 33008 50328 33014 50380
rect 57238 50368 57244 50380
rect 57199 50340 57244 50368
rect 57238 50328 57244 50340
rect 57296 50328 57302 50380
rect 57977 50371 58035 50377
rect 57977 50337 57989 50371
rect 58023 50368 58035 50371
rect 58250 50368 58256 50380
rect 58023 50340 58256 50368
rect 58023 50337 58035 50340
rect 57977 50331 58035 50337
rect 58250 50328 58256 50340
rect 58308 50328 58314 50380
rect 31536 50272 32628 50300
rect 33413 50303 33471 50309
rect 31536 50260 31542 50272
rect 33413 50269 33425 50303
rect 33459 50269 33471 50303
rect 33413 50263 33471 50269
rect 31938 50192 31944 50244
rect 31996 50232 32002 50244
rect 33428 50232 33456 50263
rect 31996 50204 33456 50232
rect 31996 50192 32002 50204
rect 28261 50167 28319 50173
rect 28261 50133 28273 50167
rect 28307 50164 28319 50167
rect 28350 50164 28356 50176
rect 28307 50136 28356 50164
rect 28307 50133 28319 50136
rect 28261 50127 28319 50133
rect 28350 50124 28356 50136
rect 28408 50124 28414 50176
rect 1104 50074 58880 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 58880 50074
rect 1104 50000 58880 50022
rect 20806 49960 20812 49972
rect 20767 49932 20812 49960
rect 20806 49920 20812 49932
rect 20864 49920 20870 49972
rect 21266 49920 21272 49972
rect 21324 49960 21330 49972
rect 21361 49963 21419 49969
rect 21361 49960 21373 49963
rect 21324 49932 21373 49960
rect 21324 49920 21330 49932
rect 21361 49929 21373 49932
rect 21407 49929 21419 49963
rect 21361 49923 21419 49929
rect 19426 49824 19432 49836
rect 19387 49796 19432 49824
rect 19426 49784 19432 49796
rect 19484 49784 19490 49836
rect 20824 49824 20852 49920
rect 21376 49892 21404 49923
rect 28994 49920 29000 49972
rect 29052 49960 29058 49972
rect 29181 49963 29239 49969
rect 29181 49960 29193 49963
rect 29052 49932 29193 49960
rect 29052 49920 29058 49932
rect 29181 49929 29193 49932
rect 29227 49929 29239 49963
rect 29181 49923 29239 49929
rect 31113 49963 31171 49969
rect 31113 49929 31125 49963
rect 31159 49960 31171 49963
rect 31478 49960 31484 49972
rect 31159 49932 31484 49960
rect 31159 49929 31171 49932
rect 31113 49923 31171 49929
rect 31478 49920 31484 49932
rect 31536 49920 31542 49972
rect 32490 49920 32496 49972
rect 32548 49960 32554 49972
rect 33137 49963 33195 49969
rect 33137 49960 33149 49963
rect 32548 49932 33149 49960
rect 32548 49920 32554 49932
rect 33137 49929 33149 49932
rect 33183 49929 33195 49963
rect 33137 49923 33195 49929
rect 33689 49963 33747 49969
rect 33689 49929 33701 49963
rect 33735 49960 33747 49963
rect 34330 49960 34336 49972
rect 33735 49932 34336 49960
rect 33735 49929 33747 49932
rect 33689 49923 33747 49929
rect 34330 49920 34336 49932
rect 34388 49920 34394 49972
rect 21376 49864 22094 49892
rect 20824 49796 21496 49824
rect 19696 49759 19754 49765
rect 19696 49725 19708 49759
rect 19742 49756 19754 49759
rect 20162 49756 20168 49768
rect 19742 49728 20168 49756
rect 19742 49725 19754 49728
rect 19696 49719 19754 49725
rect 20162 49716 20168 49728
rect 20220 49716 20226 49768
rect 20530 49716 20536 49768
rect 20588 49756 20594 49768
rect 21468 49765 21496 49796
rect 21269 49759 21327 49765
rect 21269 49756 21281 49759
rect 20588 49728 21281 49756
rect 20588 49716 20594 49728
rect 21269 49725 21281 49728
rect 21315 49725 21327 49759
rect 21269 49719 21327 49725
rect 21453 49759 21511 49765
rect 21453 49725 21465 49759
rect 21499 49725 21511 49759
rect 22066 49756 22094 49864
rect 22646 49784 22652 49836
rect 22704 49824 22710 49836
rect 23569 49827 23627 49833
rect 23569 49824 23581 49827
rect 22704 49796 23581 49824
rect 22704 49784 22710 49796
rect 23569 49793 23581 49796
rect 23615 49793 23627 49827
rect 23569 49787 23627 49793
rect 30101 49827 30159 49833
rect 30101 49793 30113 49827
rect 30147 49824 30159 49827
rect 31110 49824 31116 49836
rect 30147 49796 31116 49824
rect 30147 49793 30159 49796
rect 30101 49787 30159 49793
rect 31110 49784 31116 49796
rect 31168 49784 31174 49836
rect 31757 49827 31815 49833
rect 31757 49824 31769 49827
rect 31496 49796 31769 49824
rect 31496 49768 31524 49796
rect 31757 49793 31769 49796
rect 31803 49793 31815 49827
rect 31757 49787 31815 49793
rect 33134 49784 33140 49836
rect 33192 49824 33198 49836
rect 33192 49796 33916 49824
rect 33192 49784 33198 49796
rect 22557 49759 22615 49765
rect 22557 49756 22569 49759
rect 22066 49728 22569 49756
rect 21453 49719 21511 49725
rect 22557 49725 22569 49728
rect 22603 49725 22615 49759
rect 22557 49719 22615 49725
rect 23836 49759 23894 49765
rect 23836 49725 23848 49759
rect 23882 49756 23894 49759
rect 25222 49756 25228 49768
rect 23882 49728 25228 49756
rect 23882 49725 23894 49728
rect 23836 49719 23894 49725
rect 25222 49716 25228 49728
rect 25280 49716 25286 49768
rect 25774 49765 25780 49768
rect 25501 49759 25559 49765
rect 25501 49725 25513 49759
rect 25547 49756 25559 49759
rect 25768 49756 25780 49765
rect 25547 49728 25636 49756
rect 25735 49728 25780 49756
rect 25547 49725 25559 49728
rect 25501 49719 25559 49725
rect 25608 49688 25636 49728
rect 25768 49719 25780 49728
rect 25774 49716 25780 49719
rect 25832 49716 25838 49768
rect 26326 49756 26332 49768
rect 25884 49728 26332 49756
rect 25884 49688 25912 49728
rect 26326 49716 26332 49728
rect 26384 49756 26390 49768
rect 27522 49756 27528 49768
rect 26384 49728 27528 49756
rect 26384 49716 26390 49728
rect 27522 49716 27528 49728
rect 27580 49756 27586 49768
rect 27801 49759 27859 49765
rect 27801 49756 27813 49759
rect 27580 49728 27813 49756
rect 27580 49716 27586 49728
rect 27801 49725 27813 49728
rect 27847 49725 27859 49759
rect 27801 49719 27859 49725
rect 27890 49716 27896 49768
rect 27948 49756 27954 49768
rect 28057 49759 28115 49765
rect 28057 49756 28069 49759
rect 27948 49728 28069 49756
rect 27948 49716 27954 49728
rect 28057 49725 28069 49728
rect 28103 49725 28115 49759
rect 28057 49719 28115 49725
rect 30009 49759 30067 49765
rect 30009 49725 30021 49759
rect 30055 49756 30067 49759
rect 30193 49759 30251 49765
rect 30055 49728 30144 49756
rect 30055 49725 30067 49728
rect 30009 49719 30067 49725
rect 25608 49660 25912 49688
rect 30116 49688 30144 49728
rect 30193 49725 30205 49759
rect 30239 49756 30251 49759
rect 30466 49756 30472 49768
rect 30239 49728 30472 49756
rect 30239 49725 30251 49728
rect 30193 49719 30251 49725
rect 30466 49716 30472 49728
rect 30524 49716 30530 49768
rect 31021 49759 31079 49765
rect 31021 49725 31033 49759
rect 31067 49756 31079 49759
rect 31478 49756 31484 49768
rect 31067 49728 31484 49756
rect 31067 49725 31079 49728
rect 31021 49719 31079 49725
rect 31478 49716 31484 49728
rect 31536 49716 31542 49768
rect 31662 49756 31668 49768
rect 31623 49728 31668 49756
rect 31662 49716 31668 49728
rect 31720 49716 31726 49768
rect 31849 49759 31907 49765
rect 31849 49725 31861 49759
rect 31895 49725 31907 49759
rect 31849 49719 31907 49725
rect 33045 49759 33103 49765
rect 33045 49725 33057 49759
rect 33091 49756 33103 49759
rect 33502 49756 33508 49768
rect 33091 49728 33508 49756
rect 33091 49725 33103 49728
rect 33045 49719 33103 49725
rect 30926 49688 30932 49700
rect 30116 49660 30932 49688
rect 30926 49648 30932 49660
rect 30984 49648 30990 49700
rect 31754 49648 31760 49700
rect 31812 49688 31818 49700
rect 31864 49688 31892 49719
rect 33502 49716 33508 49728
rect 33560 49716 33566 49768
rect 33888 49765 33916 49796
rect 33873 49759 33931 49765
rect 33873 49725 33885 49759
rect 33919 49725 33931 49759
rect 33873 49719 33931 49725
rect 34238 49716 34244 49768
rect 34296 49756 34302 49768
rect 34517 49759 34575 49765
rect 34517 49756 34529 49759
rect 34296 49728 34529 49756
rect 34296 49716 34302 49728
rect 34517 49725 34529 49728
rect 34563 49725 34575 49759
rect 34698 49756 34704 49768
rect 34659 49728 34704 49756
rect 34517 49719 34575 49725
rect 34698 49716 34704 49728
rect 34756 49716 34762 49768
rect 57425 49759 57483 49765
rect 57425 49725 57437 49759
rect 57471 49756 57483 49759
rect 57514 49756 57520 49768
rect 57471 49728 57520 49756
rect 57471 49725 57483 49728
rect 57425 49719 57483 49725
rect 57514 49716 57520 49728
rect 57572 49716 57578 49768
rect 58158 49756 58164 49768
rect 58119 49728 58164 49756
rect 58158 49716 58164 49728
rect 58216 49716 58222 49768
rect 57974 49688 57980 49700
rect 31812 49660 31892 49688
rect 57935 49660 57980 49688
rect 31812 49648 31818 49660
rect 57974 49648 57980 49660
rect 58032 49648 58038 49700
rect 22370 49580 22376 49632
rect 22428 49620 22434 49632
rect 22649 49623 22707 49629
rect 22649 49620 22661 49623
rect 22428 49592 22661 49620
rect 22428 49580 22434 49592
rect 22649 49589 22661 49592
rect 22695 49589 22707 49623
rect 24946 49620 24952 49632
rect 24907 49592 24952 49620
rect 22649 49583 22707 49589
rect 24946 49580 24952 49592
rect 25004 49580 25010 49632
rect 26510 49580 26516 49632
rect 26568 49620 26574 49632
rect 26881 49623 26939 49629
rect 26881 49620 26893 49623
rect 26568 49592 26893 49620
rect 26568 49580 26574 49592
rect 26881 49589 26893 49592
rect 26927 49589 26939 49623
rect 34606 49620 34612 49632
rect 34567 49592 34612 49620
rect 26881 49583 26939 49589
rect 34606 49580 34612 49592
rect 34664 49580 34670 49632
rect 57238 49620 57244 49632
rect 57199 49592 57244 49620
rect 57238 49580 57244 49592
rect 57296 49580 57302 49632
rect 1104 49530 58880 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 50326 49530
rect 50378 49478 50390 49530
rect 50442 49478 50454 49530
rect 50506 49478 50518 49530
rect 50570 49478 58880 49530
rect 1104 49456 58880 49478
rect 21450 49416 21456 49428
rect 21411 49388 21456 49416
rect 21450 49376 21456 49388
rect 21508 49376 21514 49428
rect 25222 49416 25228 49428
rect 25183 49388 25228 49416
rect 25222 49376 25228 49388
rect 25280 49376 25286 49428
rect 25409 49419 25467 49425
rect 25409 49385 25421 49419
rect 25455 49416 25467 49419
rect 26694 49416 26700 49428
rect 25455 49388 26464 49416
rect 26655 49388 26700 49416
rect 25455 49385 25467 49388
rect 25409 49379 25467 49385
rect 22465 49351 22523 49357
rect 22465 49348 22477 49351
rect 21652 49320 22477 49348
rect 21652 49292 21680 49320
rect 22465 49317 22477 49320
rect 22511 49317 22523 49351
rect 22465 49311 22523 49317
rect 26329 49351 26387 49357
rect 26329 49317 26341 49351
rect 26375 49317 26387 49351
rect 26329 49311 26387 49317
rect 26436 49348 26464 49388
rect 26694 49376 26700 49388
rect 26752 49376 26758 49428
rect 28350 49376 28356 49428
rect 28408 49416 28414 49428
rect 33505 49419 33563 49425
rect 28408 49388 29500 49416
rect 28408 49376 28414 49388
rect 26534 49351 26592 49357
rect 26534 49348 26546 49351
rect 26436 49320 26546 49348
rect 1394 49280 1400 49292
rect 1355 49252 1400 49280
rect 1394 49240 1400 49252
rect 1452 49240 1458 49292
rect 21634 49280 21640 49292
rect 21595 49252 21640 49280
rect 21634 49240 21640 49252
rect 21692 49240 21698 49292
rect 21821 49283 21879 49289
rect 21821 49249 21833 49283
rect 21867 49280 21879 49283
rect 22370 49280 22376 49292
rect 21867 49252 22376 49280
rect 21867 49249 21879 49252
rect 21821 49243 21879 49249
rect 22370 49240 22376 49252
rect 22428 49240 22434 49292
rect 22554 49280 22560 49292
rect 22515 49252 22560 49280
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 24946 49240 24952 49292
rect 25004 49280 25010 49292
rect 25350 49283 25408 49289
rect 25350 49280 25362 49283
rect 25004 49252 25362 49280
rect 25004 49240 25010 49252
rect 25350 49249 25362 49252
rect 25396 49280 25408 49283
rect 25682 49280 25688 49292
rect 25396 49252 25688 49280
rect 25396 49249 25408 49252
rect 25350 49243 25408 49249
rect 25682 49240 25688 49252
rect 25740 49280 25746 49292
rect 25869 49283 25927 49289
rect 25869 49280 25881 49283
rect 25740 49252 25881 49280
rect 25740 49240 25746 49252
rect 25869 49249 25881 49252
rect 25915 49280 25927 49283
rect 26344 49280 26372 49311
rect 25915 49252 26372 49280
rect 25915 49249 25927 49252
rect 25869 49243 25927 49249
rect 21913 49215 21971 49221
rect 21913 49181 21925 49215
rect 21959 49212 21971 49215
rect 22572 49212 22600 49240
rect 25774 49212 25780 49224
rect 21959 49184 22600 49212
rect 25687 49184 25780 49212
rect 21959 49181 21971 49184
rect 21913 49175 21971 49181
rect 25774 49172 25780 49184
rect 25832 49212 25838 49224
rect 26436 49212 26464 49320
rect 26534 49317 26546 49320
rect 26580 49317 26592 49351
rect 26534 49311 26592 49317
rect 27700 49351 27758 49357
rect 27700 49317 27712 49351
rect 27746 49348 27758 49351
rect 29365 49351 29423 49357
rect 29365 49348 29377 49351
rect 27746 49320 29377 49348
rect 27746 49317 27758 49320
rect 27700 49311 27758 49317
rect 29365 49317 29377 49320
rect 29411 49317 29423 49351
rect 29365 49311 29423 49317
rect 29270 49280 29276 49292
rect 29231 49252 29276 49280
rect 29270 49240 29276 49252
rect 29328 49240 29334 49292
rect 29472 49289 29500 49388
rect 33505 49385 33517 49419
rect 33551 49385 33563 49419
rect 34790 49416 34796 49428
rect 34751 49388 34796 49416
rect 33505 49379 33563 49385
rect 33520 49348 33548 49379
rect 34790 49376 34796 49388
rect 34848 49376 34854 49428
rect 57974 49376 57980 49428
rect 58032 49416 58038 49428
rect 58161 49419 58219 49425
rect 58161 49416 58173 49419
rect 58032 49388 58173 49416
rect 58032 49376 58038 49388
rect 58161 49385 58173 49388
rect 58207 49385 58219 49419
rect 58161 49379 58219 49385
rect 34422 49348 34428 49360
rect 34480 49357 34486 49360
rect 34480 49351 34509 49357
rect 33428 49320 33548 49348
rect 33980 49320 34428 49348
rect 31294 49289 31300 49292
rect 29457 49283 29515 49289
rect 29457 49249 29469 49283
rect 29503 49249 29515 49283
rect 29457 49243 29515 49249
rect 31288 49243 31300 49289
rect 31352 49280 31358 49292
rect 31352 49252 31388 49280
rect 31294 49240 31300 49243
rect 31352 49240 31358 49252
rect 27430 49212 27436 49224
rect 25832 49184 26464 49212
rect 27391 49184 27436 49212
rect 25832 49172 25838 49184
rect 27430 49172 27436 49184
rect 27488 49172 27494 49224
rect 30650 49172 30656 49224
rect 30708 49212 30714 49224
rect 31021 49215 31079 49221
rect 31021 49212 31033 49215
rect 30708 49184 31033 49212
rect 30708 49172 30714 49184
rect 31021 49181 31033 49184
rect 31067 49181 31079 49215
rect 33428 49212 33456 49320
rect 33980 49289 34008 49320
rect 34422 49308 34428 49320
rect 34497 49317 34509 49351
rect 34480 49311 34509 49317
rect 34641 49351 34699 49357
rect 34641 49317 34653 49351
rect 34687 49348 34699 49351
rect 35250 49348 35256 49360
rect 34687 49320 35256 49348
rect 34687 49317 34699 49320
rect 34641 49311 34699 49317
rect 34480 49308 34486 49311
rect 35250 49308 35256 49320
rect 35308 49308 35314 49360
rect 33502 49283 33560 49289
rect 33502 49249 33514 49283
rect 33548 49280 33560 49283
rect 33965 49283 34023 49289
rect 33965 49280 33977 49283
rect 33548 49252 33977 49280
rect 33548 49249 33560 49252
rect 33502 49243 33560 49249
rect 33965 49249 33977 49252
rect 34011 49249 34023 49283
rect 33965 49243 34023 49249
rect 55030 49240 55036 49292
rect 55088 49280 55094 49292
rect 56873 49283 56931 49289
rect 56873 49280 56885 49283
rect 55088 49252 56885 49280
rect 55088 49240 55094 49252
rect 56873 49249 56885 49252
rect 56919 49249 56931 49283
rect 56873 49243 56931 49249
rect 57238 49240 57244 49292
rect 57296 49280 57302 49292
rect 57701 49283 57759 49289
rect 57701 49280 57713 49283
rect 57296 49252 57713 49280
rect 57296 49240 57302 49252
rect 57701 49249 57713 49252
rect 57747 49249 57759 49283
rect 57701 49243 57759 49249
rect 33686 49212 33692 49224
rect 33428 49184 33692 49212
rect 31021 49175 31079 49181
rect 33686 49172 33692 49184
rect 33744 49212 33750 49224
rect 33873 49215 33931 49221
rect 33873 49212 33885 49215
rect 33744 49184 33885 49212
rect 33744 49172 33750 49184
rect 33873 49181 33885 49184
rect 33919 49181 33931 49215
rect 33873 49175 33931 49181
rect 26510 49076 26516 49088
rect 26471 49048 26516 49076
rect 26510 49036 26516 49048
rect 26568 49036 26574 49088
rect 28442 49036 28448 49088
rect 28500 49076 28506 49088
rect 28813 49079 28871 49085
rect 28813 49076 28825 49079
rect 28500 49048 28825 49076
rect 28500 49036 28506 49048
rect 28813 49045 28825 49048
rect 28859 49045 28871 49079
rect 28813 49039 28871 49045
rect 31754 49036 31760 49088
rect 31812 49076 31818 49088
rect 32401 49079 32459 49085
rect 32401 49076 32413 49079
rect 31812 49048 32413 49076
rect 31812 49036 31818 49048
rect 32401 49045 32413 49048
rect 32447 49045 32459 49079
rect 33318 49076 33324 49088
rect 33279 49048 33324 49076
rect 32401 49039 32459 49045
rect 33318 49036 33324 49048
rect 33376 49036 33382 49088
rect 33888 49076 33916 49175
rect 57422 49172 57428 49224
rect 57480 49212 57486 49224
rect 57517 49215 57575 49221
rect 57517 49212 57529 49215
rect 57480 49184 57529 49212
rect 57480 49172 57486 49184
rect 57517 49181 57529 49184
rect 57563 49181 57575 49215
rect 57517 49175 57575 49181
rect 57054 49144 57060 49156
rect 57015 49116 57060 49144
rect 57054 49104 57060 49116
rect 57112 49104 57118 49156
rect 34609 49079 34667 49085
rect 34609 49076 34621 49079
rect 33888 49048 34621 49076
rect 34609 49045 34621 49048
rect 34655 49045 34667 49079
rect 34609 49039 34667 49045
rect 1104 48986 58880 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 58880 48986
rect 1104 48912 58880 48934
rect 20438 48872 20444 48884
rect 20399 48844 20444 48872
rect 20438 48832 20444 48844
rect 20496 48832 20502 48884
rect 20530 48832 20536 48884
rect 20588 48872 20594 48884
rect 20625 48875 20683 48881
rect 20625 48872 20637 48875
rect 20588 48844 20637 48872
rect 20588 48832 20594 48844
rect 20625 48841 20637 48844
rect 20671 48841 20683 48875
rect 25498 48872 25504 48884
rect 25459 48844 25504 48872
rect 20625 48835 20683 48841
rect 20640 48736 20668 48835
rect 25498 48832 25504 48844
rect 25556 48832 25562 48884
rect 30466 48872 30472 48884
rect 30427 48844 30472 48872
rect 30466 48832 30472 48844
rect 30524 48832 30530 48884
rect 30926 48832 30932 48884
rect 30984 48872 30990 48884
rect 31297 48875 31355 48881
rect 31297 48872 31309 48875
rect 30984 48844 31309 48872
rect 30984 48832 30990 48844
rect 31297 48841 31309 48844
rect 31343 48841 31355 48875
rect 31297 48835 31355 48841
rect 31662 48832 31668 48884
rect 31720 48872 31726 48884
rect 31941 48875 31999 48881
rect 31941 48872 31953 48875
rect 31720 48844 31953 48872
rect 31720 48832 31726 48844
rect 31941 48841 31953 48844
rect 31987 48841 31999 48875
rect 34422 48872 34428 48884
rect 34383 48844 34428 48872
rect 31941 48835 31999 48841
rect 34422 48832 34428 48844
rect 34480 48832 34486 48884
rect 35250 48832 35256 48884
rect 35308 48872 35314 48884
rect 36265 48875 36323 48881
rect 36265 48872 36277 48875
rect 35308 48844 36277 48872
rect 35308 48832 35314 48844
rect 36265 48841 36277 48844
rect 36311 48841 36323 48875
rect 57422 48872 57428 48884
rect 57383 48844 57428 48872
rect 36265 48835 36323 48841
rect 57422 48832 57428 48844
rect 57480 48832 57486 48884
rect 24949 48739 25007 48745
rect 20640 48708 21312 48736
rect 18138 48668 18144 48680
rect 18099 48640 18144 48668
rect 18138 48628 18144 48640
rect 18196 48628 18202 48680
rect 21082 48668 21088 48680
rect 21043 48640 21088 48668
rect 21082 48628 21088 48640
rect 21140 48628 21146 48680
rect 21284 48677 21312 48708
rect 24949 48705 24961 48739
rect 24995 48736 25007 48739
rect 24995 48708 25820 48736
rect 24995 48705 25007 48708
rect 24949 48699 25007 48705
rect 25792 48680 25820 48708
rect 27522 48696 27528 48748
rect 27580 48736 27586 48748
rect 29089 48739 29147 48745
rect 29089 48736 29101 48739
rect 27580 48708 29101 48736
rect 27580 48696 27586 48708
rect 29089 48705 29101 48708
rect 29135 48705 29147 48739
rect 30484 48736 30512 48832
rect 30650 48764 30656 48816
rect 30708 48804 30714 48816
rect 30708 48776 31754 48804
rect 30708 48764 30714 48776
rect 31389 48739 31447 48745
rect 31389 48736 31401 48739
rect 30484 48708 31401 48736
rect 29089 48699 29147 48705
rect 31389 48705 31401 48708
rect 31435 48705 31447 48739
rect 31726 48736 31754 48776
rect 31726 48708 33088 48736
rect 31389 48699 31447 48705
rect 21269 48671 21327 48677
rect 21269 48637 21281 48671
rect 21315 48637 21327 48671
rect 24854 48668 24860 48680
rect 24815 48640 24860 48668
rect 21269 48631 21327 48637
rect 24854 48628 24860 48640
rect 24912 48628 24918 48680
rect 25682 48668 25688 48680
rect 25643 48640 25688 48668
rect 25682 48628 25688 48640
rect 25740 48628 25746 48680
rect 25774 48628 25780 48680
rect 25832 48668 25838 48680
rect 26694 48668 26700 48680
rect 25832 48640 25877 48668
rect 26655 48640 26700 48668
rect 25832 48628 25838 48640
rect 26694 48628 26700 48640
rect 26752 48628 26758 48680
rect 27798 48668 27804 48680
rect 27759 48640 27804 48668
rect 27798 48628 27804 48640
rect 27856 48628 27862 48680
rect 28442 48668 28448 48680
rect 28403 48640 28448 48668
rect 28442 48628 28448 48640
rect 28500 48628 28506 48680
rect 31110 48668 31116 48680
rect 31071 48640 31116 48668
rect 31110 48628 31116 48640
rect 31168 48628 31174 48680
rect 33060 48677 33088 48708
rect 34330 48696 34336 48748
rect 34388 48736 34394 48748
rect 34885 48739 34943 48745
rect 34885 48736 34897 48739
rect 34388 48708 34897 48736
rect 34388 48696 34394 48708
rect 34885 48705 34897 48708
rect 34931 48705 34943 48739
rect 34885 48699 34943 48705
rect 33318 48677 33324 48680
rect 31849 48671 31907 48677
rect 31849 48668 31861 48671
rect 31726 48640 31861 48668
rect 18414 48609 18420 48612
rect 18408 48563 18420 48609
rect 18472 48600 18478 48612
rect 20257 48603 20315 48609
rect 20257 48600 20269 48603
rect 18472 48572 18508 48600
rect 19536 48572 20269 48600
rect 18414 48560 18420 48563
rect 18472 48560 18478 48572
rect 19334 48492 19340 48544
rect 19392 48532 19398 48544
rect 19536 48541 19564 48572
rect 20257 48569 20269 48572
rect 20303 48600 20315 48603
rect 20346 48600 20352 48612
rect 20303 48572 20352 48600
rect 20303 48569 20315 48572
rect 20257 48563 20315 48569
rect 20346 48560 20352 48572
rect 20404 48560 20410 48612
rect 20530 48609 20536 48612
rect 20473 48603 20536 48609
rect 20473 48569 20485 48603
rect 20519 48569 20536 48603
rect 20473 48563 20536 48569
rect 20530 48560 20536 48563
rect 20588 48560 20594 48612
rect 25501 48603 25559 48609
rect 25501 48569 25513 48603
rect 25547 48600 25559 48603
rect 26510 48600 26516 48612
rect 25547 48572 26516 48600
rect 25547 48569 25559 48572
rect 25501 48563 25559 48569
rect 26510 48560 26516 48572
rect 26568 48560 26574 48612
rect 29356 48603 29414 48609
rect 29356 48569 29368 48603
rect 29402 48600 29414 48603
rect 30929 48603 30987 48609
rect 30929 48600 30941 48603
rect 29402 48572 30941 48600
rect 29402 48569 29414 48572
rect 29356 48563 29414 48569
rect 30929 48569 30941 48572
rect 30975 48569 30987 48603
rect 31128 48600 31156 48628
rect 31726 48600 31754 48640
rect 31849 48637 31861 48640
rect 31895 48637 31907 48671
rect 31849 48631 31907 48637
rect 33045 48671 33103 48677
rect 33045 48637 33057 48671
rect 33091 48637 33103 48671
rect 33312 48668 33324 48677
rect 33279 48640 33324 48668
rect 33045 48631 33103 48637
rect 33312 48631 33324 48640
rect 31128 48572 31754 48600
rect 33060 48600 33088 48631
rect 33318 48628 33324 48631
rect 33376 48628 33382 48680
rect 34348 48600 34376 48696
rect 56502 48628 56508 48680
rect 56560 48668 56566 48680
rect 56597 48671 56655 48677
rect 56597 48668 56609 48671
rect 56560 48640 56609 48668
rect 56560 48628 56566 48640
rect 56597 48637 56609 48640
rect 56643 48637 56655 48671
rect 56597 48631 56655 48637
rect 33060 48572 34376 48600
rect 30929 48563 30987 48569
rect 34606 48560 34612 48612
rect 34664 48600 34670 48612
rect 35130 48603 35188 48609
rect 35130 48600 35142 48603
rect 34664 48572 35142 48600
rect 34664 48560 34670 48572
rect 35130 48569 35142 48572
rect 35176 48569 35188 48603
rect 57974 48600 57980 48612
rect 57935 48572 57980 48600
rect 35130 48563 35188 48569
rect 57974 48560 57980 48572
rect 58032 48560 58038 48612
rect 19521 48535 19579 48541
rect 19521 48532 19533 48535
rect 19392 48504 19533 48532
rect 19392 48492 19398 48504
rect 19521 48501 19533 48504
rect 19567 48501 19579 48535
rect 21174 48532 21180 48544
rect 21135 48504 21180 48532
rect 19521 48495 19579 48501
rect 21174 48492 21180 48504
rect 21232 48492 21238 48544
rect 26602 48492 26608 48544
rect 26660 48532 26666 48544
rect 26789 48535 26847 48541
rect 26789 48532 26801 48535
rect 26660 48504 26801 48532
rect 26660 48492 26666 48504
rect 26789 48501 26801 48504
rect 26835 48501 26847 48535
rect 26789 48495 26847 48501
rect 27706 48492 27712 48544
rect 27764 48532 27770 48544
rect 27893 48535 27951 48541
rect 27893 48532 27905 48535
rect 27764 48504 27905 48532
rect 27764 48492 27770 48504
rect 27893 48501 27905 48504
rect 27939 48501 27951 48535
rect 28534 48532 28540 48544
rect 28495 48504 28540 48532
rect 27893 48495 27951 48501
rect 28534 48492 28540 48504
rect 28592 48492 28598 48544
rect 57882 48492 57888 48544
rect 57940 48532 57946 48544
rect 58069 48535 58127 48541
rect 58069 48532 58081 48535
rect 57940 48504 58081 48532
rect 57940 48492 57946 48504
rect 58069 48501 58081 48504
rect 58115 48501 58127 48535
rect 58069 48495 58127 48501
rect 1104 48442 58880 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 50326 48442
rect 50378 48390 50390 48442
rect 50442 48390 50454 48442
rect 50506 48390 50518 48442
rect 50570 48390 58880 48442
rect 1104 48368 58880 48390
rect 15197 48331 15255 48337
rect 15197 48297 15209 48331
rect 15243 48297 15255 48331
rect 18414 48328 18420 48340
rect 18375 48300 18420 48328
rect 15197 48291 15255 48297
rect 15212 48260 15240 48291
rect 18414 48288 18420 48300
rect 18472 48288 18478 48340
rect 18601 48331 18659 48337
rect 18601 48297 18613 48331
rect 18647 48297 18659 48331
rect 31294 48328 31300 48340
rect 31255 48300 31300 48328
rect 18601 48291 18659 48297
rect 16482 48269 16488 48272
rect 16209 48263 16267 48269
rect 16209 48260 16221 48263
rect 15120 48232 15240 48260
rect 15764 48232 16221 48260
rect 1394 48192 1400 48204
rect 1355 48164 1400 48192
rect 1394 48152 1400 48164
rect 1452 48152 1458 48204
rect 15120 48124 15148 48232
rect 15194 48195 15252 48201
rect 15194 48161 15206 48195
rect 15240 48192 15252 48195
rect 15764 48192 15792 48232
rect 16209 48229 16221 48232
rect 16255 48229 16267 48263
rect 16209 48223 16267 48229
rect 16425 48263 16488 48269
rect 16425 48229 16437 48263
rect 16471 48229 16488 48263
rect 16425 48223 16488 48229
rect 16482 48220 16488 48223
rect 16540 48220 16546 48272
rect 18616 48260 18644 48291
rect 31294 48288 31300 48300
rect 31352 48288 31358 48340
rect 33686 48328 33692 48340
rect 33647 48300 33692 48328
rect 33686 48288 33692 48300
rect 33744 48288 33750 48340
rect 34422 48328 34428 48340
rect 34383 48300 34428 48328
rect 34422 48288 34428 48300
rect 34480 48288 34486 48340
rect 57974 48288 57980 48340
rect 58032 48328 58038 48340
rect 58161 48331 58219 48337
rect 58161 48328 58173 48331
rect 58032 48300 58173 48328
rect 58032 48288 58038 48300
rect 58161 48297 58173 48300
rect 58207 48297 58219 48331
rect 58161 48291 58219 48297
rect 18524 48232 18644 48260
rect 20800 48263 20858 48269
rect 15240 48164 15792 48192
rect 15240 48161 15252 48164
rect 15194 48155 15252 48161
rect 15764 48136 15792 48164
rect 16114 48152 16120 48204
rect 16172 48192 16178 48204
rect 17037 48195 17095 48201
rect 17037 48192 17049 48195
rect 16172 48164 17049 48192
rect 16172 48152 16178 48164
rect 17037 48161 17049 48164
rect 17083 48161 17095 48195
rect 17037 48155 17095 48161
rect 17221 48195 17279 48201
rect 17221 48161 17233 48195
rect 17267 48192 17279 48195
rect 17954 48192 17960 48204
rect 17267 48164 17960 48192
rect 17267 48161 17279 48164
rect 17221 48155 17279 48161
rect 15565 48127 15623 48133
rect 15565 48124 15577 48127
rect 15120 48096 15577 48124
rect 15565 48093 15577 48096
rect 15611 48093 15623 48127
rect 15565 48087 15623 48093
rect 15657 48127 15715 48133
rect 15657 48093 15669 48127
rect 15703 48124 15715 48127
rect 15746 48124 15752 48136
rect 15703 48096 15752 48124
rect 15703 48093 15715 48096
rect 15657 48087 15715 48093
rect 15010 47988 15016 48000
rect 14971 47960 15016 47988
rect 15010 47948 15016 47960
rect 15068 47948 15074 48000
rect 15580 47988 15608 48087
rect 15746 48084 15752 48096
rect 15804 48084 15810 48136
rect 16577 48059 16635 48065
rect 16577 48025 16589 48059
rect 16623 48056 16635 48059
rect 17236 48056 17264 48155
rect 17954 48152 17960 48164
rect 18012 48152 18018 48204
rect 18524 48124 18552 48232
rect 20800 48229 20812 48263
rect 20846 48260 20858 48263
rect 21174 48260 21180 48272
rect 20846 48232 21180 48260
rect 20846 48229 20858 48232
rect 20800 48223 20858 48229
rect 21174 48220 21180 48232
rect 21232 48220 21238 48272
rect 27522 48260 27528 48272
rect 25608 48232 27528 48260
rect 18598 48195 18656 48201
rect 18598 48161 18610 48195
rect 18644 48192 18656 48195
rect 19061 48195 19119 48201
rect 19061 48192 19073 48195
rect 18644 48164 19073 48192
rect 18644 48161 18656 48164
rect 18598 48155 18656 48161
rect 19061 48161 19073 48164
rect 19107 48192 19119 48195
rect 19334 48192 19340 48204
rect 19107 48164 19340 48192
rect 19107 48161 19119 48164
rect 19061 48155 19119 48161
rect 19334 48152 19340 48164
rect 19392 48152 19398 48204
rect 23661 48195 23719 48201
rect 23661 48161 23673 48195
rect 23707 48161 23719 48195
rect 23661 48155 23719 48161
rect 24121 48195 24179 48201
rect 24121 48161 24133 48195
rect 24167 48192 24179 48195
rect 24210 48192 24216 48204
rect 24167 48164 24216 48192
rect 24167 48161 24179 48164
rect 24121 48155 24179 48161
rect 18524 48096 19012 48124
rect 18984 48065 19012 48096
rect 19426 48084 19432 48136
rect 19484 48124 19490 48136
rect 20533 48127 20591 48133
rect 20533 48124 20545 48127
rect 19484 48096 20545 48124
rect 19484 48084 19490 48096
rect 20533 48093 20545 48096
rect 20579 48093 20591 48127
rect 23676 48124 23704 48155
rect 24210 48152 24216 48164
rect 24268 48152 24274 48204
rect 24305 48195 24363 48201
rect 24305 48161 24317 48195
rect 24351 48192 24363 48195
rect 25314 48192 25320 48204
rect 24351 48164 25320 48192
rect 24351 48161 24363 48164
rect 24305 48155 24363 48161
rect 25314 48152 25320 48164
rect 25372 48152 25378 48204
rect 25608 48201 25636 48232
rect 27522 48220 27528 48232
rect 27580 48220 27586 48272
rect 28534 48220 28540 48272
rect 28592 48260 28598 48272
rect 28629 48263 28687 48269
rect 28629 48260 28641 48263
rect 28592 48232 28641 48260
rect 28592 48220 28598 48232
rect 28629 48229 28641 48232
rect 28675 48229 28687 48263
rect 28629 48223 28687 48229
rect 30926 48220 30932 48272
rect 30984 48260 30990 48272
rect 32309 48263 32367 48269
rect 32309 48260 32321 48263
rect 30984 48232 32321 48260
rect 30984 48220 30990 48232
rect 32309 48229 32321 48232
rect 32355 48229 32367 48263
rect 33704 48260 33732 48288
rect 34241 48263 34299 48269
rect 33704 48232 34100 48260
rect 32309 48223 32367 48229
rect 25593 48195 25651 48201
rect 25593 48161 25605 48195
rect 25639 48161 25651 48195
rect 25593 48155 25651 48161
rect 25860 48195 25918 48201
rect 25860 48161 25872 48195
rect 25906 48192 25918 48195
rect 26326 48192 26332 48204
rect 25906 48164 26332 48192
rect 25906 48161 25918 48164
rect 25860 48155 25918 48161
rect 26326 48152 26332 48164
rect 26384 48152 26390 48204
rect 27893 48195 27951 48201
rect 27893 48161 27905 48195
rect 27939 48192 27951 48195
rect 28552 48192 28580 48220
rect 27939 48164 28580 48192
rect 28813 48195 28871 48201
rect 27939 48161 27951 48164
rect 27893 48155 27951 48161
rect 28813 48161 28825 48195
rect 28859 48161 28871 48195
rect 28813 48155 28871 48161
rect 30469 48195 30527 48201
rect 30469 48161 30481 48195
rect 30515 48161 30527 48195
rect 31478 48192 31484 48204
rect 31439 48164 31484 48192
rect 30469 48155 30527 48161
rect 25130 48124 25136 48136
rect 23676 48096 25136 48124
rect 20533 48087 20591 48093
rect 25130 48084 25136 48096
rect 25188 48084 25194 48136
rect 27706 48084 27712 48136
rect 27764 48124 27770 48136
rect 28169 48127 28227 48133
rect 28169 48124 28181 48127
rect 27764 48096 28181 48124
rect 27764 48084 27770 48096
rect 28169 48093 28181 48096
rect 28215 48124 28227 48127
rect 28828 48124 28856 48155
rect 28215 48096 28856 48124
rect 30484 48124 30512 48155
rect 31478 48152 31484 48164
rect 31536 48152 31542 48204
rect 31662 48192 31668 48204
rect 31623 48164 31668 48192
rect 31662 48152 31668 48164
rect 31720 48152 31726 48204
rect 31754 48152 31760 48204
rect 31812 48192 31818 48204
rect 32214 48192 32220 48204
rect 31812 48164 31857 48192
rect 32175 48164 32220 48192
rect 31812 48152 31818 48164
rect 32214 48152 32220 48164
rect 32272 48152 32278 48204
rect 33042 48192 33048 48204
rect 33003 48164 33048 48192
rect 33042 48152 33048 48164
rect 33100 48152 33106 48204
rect 33597 48195 33655 48201
rect 33597 48161 33609 48195
rect 33643 48192 33655 48195
rect 33686 48192 33692 48204
rect 33643 48164 33692 48192
rect 33643 48161 33655 48164
rect 33597 48155 33655 48161
rect 33686 48152 33692 48164
rect 33744 48152 33750 48204
rect 34072 48192 34100 48232
rect 34241 48229 34253 48263
rect 34287 48260 34299 48263
rect 35250 48260 35256 48272
rect 34287 48232 35256 48260
rect 34287 48229 34299 48232
rect 34241 48223 34299 48229
rect 35250 48220 35256 48232
rect 35308 48220 35314 48272
rect 34517 48195 34575 48201
rect 34517 48192 34529 48195
rect 34072 48164 34529 48192
rect 34517 48161 34529 48164
rect 34563 48161 34575 48195
rect 34517 48155 34575 48161
rect 31846 48124 31852 48136
rect 30484 48096 31852 48124
rect 28215 48093 28227 48096
rect 28169 48087 28227 48093
rect 31846 48084 31852 48096
rect 31904 48084 31910 48136
rect 57057 48127 57115 48133
rect 57057 48093 57069 48127
rect 57103 48124 57115 48127
rect 57517 48127 57575 48133
rect 57517 48124 57529 48127
rect 57103 48096 57529 48124
rect 57103 48093 57115 48096
rect 57057 48087 57115 48093
rect 57517 48093 57529 48096
rect 57563 48093 57575 48127
rect 57698 48124 57704 48136
rect 57659 48096 57704 48124
rect 57517 48087 57575 48093
rect 57698 48084 57704 48096
rect 57756 48084 57762 48136
rect 16623 48028 17264 48056
rect 18969 48059 19027 48065
rect 16623 48025 16635 48028
rect 16577 48019 16635 48025
rect 18969 48025 18981 48059
rect 19015 48056 19027 48059
rect 20438 48056 20444 48068
rect 19015 48028 20444 48056
rect 19015 48025 19027 48028
rect 18969 48019 19027 48025
rect 20438 48016 20444 48028
rect 20496 48016 20502 48068
rect 23474 48056 23480 48068
rect 23435 48028 23480 48056
rect 23474 48016 23480 48028
rect 23532 48016 23538 48068
rect 26973 48059 27031 48065
rect 26973 48025 26985 48059
rect 27019 48056 27031 48059
rect 27798 48056 27804 48068
rect 27019 48028 27804 48056
rect 27019 48025 27031 48028
rect 26973 48019 27031 48025
rect 27798 48016 27804 48028
rect 27856 48016 27862 48068
rect 29270 48056 29276 48068
rect 28000 48028 29276 48056
rect 16390 47988 16396 48000
rect 15580 47960 16396 47988
rect 16390 47948 16396 47960
rect 16448 47948 16454 48000
rect 17037 47991 17095 47997
rect 17037 47957 17049 47991
rect 17083 47988 17095 47991
rect 17402 47988 17408 48000
rect 17083 47960 17408 47988
rect 17083 47957 17095 47960
rect 17037 47951 17095 47957
rect 17402 47948 17408 47960
rect 17460 47948 17466 48000
rect 20530 47948 20536 48000
rect 20588 47988 20594 48000
rect 21913 47991 21971 47997
rect 21913 47988 21925 47991
rect 20588 47960 21925 47988
rect 20588 47948 20594 47960
rect 21913 47957 21925 47960
rect 21959 47957 21971 47991
rect 21913 47951 21971 47957
rect 24213 47991 24271 47997
rect 24213 47957 24225 47991
rect 24259 47988 24271 47991
rect 24854 47988 24860 48000
rect 24259 47960 24860 47988
rect 24259 47957 24271 47960
rect 24213 47951 24271 47957
rect 24854 47948 24860 47960
rect 24912 47988 24918 48000
rect 25406 47988 25412 48000
rect 24912 47960 25412 47988
rect 24912 47948 24918 47960
rect 25406 47948 25412 47960
rect 25464 47948 25470 48000
rect 27709 47991 27767 47997
rect 27709 47957 27721 47991
rect 27755 47988 27767 47991
rect 28000 47988 28028 48028
rect 29270 48016 29276 48028
rect 29328 48016 29334 48068
rect 34238 48056 34244 48068
rect 34199 48028 34244 48056
rect 34238 48016 34244 48028
rect 34296 48016 34302 48068
rect 27755 47960 28028 47988
rect 27755 47957 27767 47960
rect 27709 47951 27767 47957
rect 28074 47948 28080 48000
rect 28132 47988 28138 48000
rect 28132 47960 28177 47988
rect 28132 47948 28138 47960
rect 28258 47948 28264 48000
rect 28316 47988 28322 48000
rect 28997 47991 29055 47997
rect 28997 47988 29009 47991
rect 28316 47960 29009 47988
rect 28316 47948 28322 47960
rect 28997 47957 29009 47960
rect 29043 47957 29055 47991
rect 28997 47951 29055 47957
rect 29914 47948 29920 48000
rect 29972 47988 29978 48000
rect 30561 47991 30619 47997
rect 30561 47988 30573 47991
rect 29972 47960 30573 47988
rect 29972 47948 29978 47960
rect 30561 47957 30573 47960
rect 30607 47957 30619 47991
rect 30561 47951 30619 47957
rect 31754 47948 31760 48000
rect 31812 47988 31818 48000
rect 31938 47988 31944 48000
rect 31812 47960 31944 47988
rect 31812 47948 31818 47960
rect 31938 47948 31944 47960
rect 31996 47988 32002 48000
rect 32861 47991 32919 47997
rect 32861 47988 32873 47991
rect 31996 47960 32873 47988
rect 31996 47948 32002 47960
rect 32861 47957 32873 47960
rect 32907 47957 32919 47991
rect 32861 47951 32919 47957
rect 1104 47898 58880 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 58880 47898
rect 1104 47824 58880 47846
rect 16482 47744 16488 47796
rect 16540 47784 16546 47796
rect 18693 47787 18751 47793
rect 18693 47784 18705 47787
rect 16540 47756 18705 47784
rect 16540 47744 16546 47756
rect 18693 47753 18705 47756
rect 18739 47753 18751 47787
rect 18693 47747 18751 47753
rect 20165 47787 20223 47793
rect 20165 47753 20177 47787
rect 20211 47784 20223 47787
rect 21082 47784 21088 47796
rect 20211 47756 21088 47784
rect 20211 47753 20223 47756
rect 20165 47747 20223 47753
rect 21082 47744 21088 47756
rect 21140 47744 21146 47796
rect 25314 47784 25320 47796
rect 25275 47756 25320 47784
rect 25314 47744 25320 47756
rect 25372 47744 25378 47796
rect 26326 47784 26332 47796
rect 26287 47756 26332 47784
rect 26326 47744 26332 47756
rect 26384 47744 26390 47796
rect 26694 47744 26700 47796
rect 26752 47784 26758 47796
rect 26789 47787 26847 47793
rect 26789 47784 26801 47787
rect 26752 47756 26801 47784
rect 26752 47744 26758 47756
rect 26789 47753 26801 47756
rect 26835 47784 26847 47787
rect 28074 47784 28080 47796
rect 26835 47756 28080 47784
rect 26835 47753 26847 47756
rect 26789 47747 26847 47753
rect 28074 47744 28080 47756
rect 28132 47784 28138 47796
rect 29914 47784 29920 47796
rect 28132 47756 28304 47784
rect 29875 47756 29920 47784
rect 28132 47744 28138 47756
rect 27798 47716 27804 47728
rect 26620 47688 27804 47716
rect 18782 47608 18788 47660
rect 18840 47648 18846 47660
rect 19245 47651 19303 47657
rect 19245 47648 19257 47651
rect 18840 47620 19257 47648
rect 18840 47608 18846 47620
rect 19245 47617 19257 47620
rect 19291 47648 19303 47651
rect 26620 47648 26648 47688
rect 27798 47676 27804 47688
rect 27856 47676 27862 47728
rect 28276 47657 28304 47756
rect 29914 47744 29920 47756
rect 29972 47744 29978 47796
rect 32214 47784 32220 47796
rect 30024 47756 32220 47784
rect 19291 47620 20944 47648
rect 19291 47617 19303 47620
rect 19245 47611 19303 47617
rect 1394 47580 1400 47592
rect 1355 47552 1400 47580
rect 1394 47540 1400 47552
rect 1452 47540 1458 47592
rect 13906 47540 13912 47592
rect 13964 47580 13970 47592
rect 14369 47583 14427 47589
rect 14369 47580 14381 47583
rect 13964 47552 14381 47580
rect 13964 47540 13970 47552
rect 14369 47549 14381 47552
rect 14415 47549 14427 47583
rect 14369 47543 14427 47549
rect 14636 47583 14694 47589
rect 14636 47549 14648 47583
rect 14682 47580 14694 47583
rect 15010 47580 15016 47592
rect 14682 47552 15016 47580
rect 14682 47549 14694 47552
rect 14636 47543 14694 47549
rect 15010 47540 15016 47552
rect 15068 47540 15074 47592
rect 17313 47583 17371 47589
rect 17313 47549 17325 47583
rect 17359 47549 17371 47583
rect 17313 47543 17371 47549
rect 17328 47512 17356 47543
rect 17402 47540 17408 47592
rect 17460 47580 17466 47592
rect 17569 47583 17627 47589
rect 17569 47580 17581 47583
rect 17460 47552 17581 47580
rect 17460 47540 17466 47552
rect 17569 47549 17581 47552
rect 17615 47549 17627 47583
rect 19150 47580 19156 47592
rect 19111 47552 19156 47580
rect 17569 47543 17627 47549
rect 19150 47540 19156 47552
rect 19208 47540 19214 47592
rect 19334 47580 19340 47592
rect 19295 47552 19340 47580
rect 19334 47540 19340 47552
rect 19392 47540 19398 47592
rect 20346 47580 20352 47592
rect 20307 47552 20352 47580
rect 20346 47540 20352 47552
rect 20404 47540 20410 47592
rect 20438 47540 20444 47592
rect 20496 47580 20502 47592
rect 20916 47589 20944 47620
rect 26528 47620 26648 47648
rect 28261 47651 28319 47657
rect 20901 47583 20959 47589
rect 20496 47552 20668 47580
rect 20496 47540 20502 47552
rect 18138 47512 18144 47524
rect 17328 47484 18144 47512
rect 18138 47472 18144 47484
rect 18196 47512 18202 47524
rect 19426 47512 19432 47524
rect 18196 47484 19432 47512
rect 18196 47472 18202 47484
rect 19426 47472 19432 47484
rect 19484 47472 19490 47524
rect 20165 47515 20223 47521
rect 20165 47481 20177 47515
rect 20211 47512 20223 47515
rect 20530 47512 20536 47524
rect 20211 47484 20536 47512
rect 20211 47481 20223 47484
rect 20165 47475 20223 47481
rect 20530 47472 20536 47484
rect 20588 47472 20594 47524
rect 20640 47512 20668 47552
rect 20901 47549 20913 47583
rect 20947 47549 20959 47583
rect 20901 47543 20959 47549
rect 23566 47540 23572 47592
rect 23624 47580 23630 47592
rect 26528 47589 26556 47620
rect 28261 47617 28273 47651
rect 28307 47617 28319 47651
rect 30024 47648 30052 47756
rect 32214 47744 32220 47756
rect 32272 47744 32278 47796
rect 57241 47787 57299 47793
rect 57241 47753 57253 47787
rect 57287 47784 57299 47787
rect 57698 47784 57704 47796
rect 57287 47756 57704 47784
rect 57287 47753 57299 47756
rect 57241 47747 57299 47753
rect 57698 47744 57704 47756
rect 57756 47744 57762 47796
rect 28261 47611 28319 47617
rect 29748 47620 30052 47648
rect 29748 47592 29776 47620
rect 23937 47583 23995 47589
rect 23937 47580 23949 47583
rect 23624 47552 23949 47580
rect 23624 47540 23630 47552
rect 23937 47549 23949 47552
rect 23983 47549 23995 47583
rect 23937 47543 23995 47549
rect 26513 47583 26571 47589
rect 26513 47549 26525 47583
rect 26559 47549 26571 47583
rect 26513 47543 26571 47549
rect 26602 47540 26608 47592
rect 26660 47580 26666 47592
rect 26881 47583 26939 47589
rect 26660 47552 26705 47580
rect 26660 47540 26666 47552
rect 26881 47549 26893 47583
rect 26927 47580 26939 47583
rect 27706 47580 27712 47592
rect 26927 47552 27712 47580
rect 26927 47549 26939 47552
rect 26881 47543 26939 47549
rect 27706 47540 27712 47552
rect 27764 47540 27770 47592
rect 27801 47583 27859 47589
rect 27801 47549 27813 47583
rect 27847 47549 27859 47583
rect 27801 47543 27859 47549
rect 20993 47515 21051 47521
rect 20993 47512 21005 47515
rect 20640 47484 21005 47512
rect 20993 47481 21005 47484
rect 21039 47481 21051 47515
rect 20993 47475 21051 47481
rect 24204 47515 24262 47521
rect 24204 47481 24216 47515
rect 24250 47512 24262 47515
rect 25222 47512 25228 47524
rect 24250 47484 25228 47512
rect 24250 47481 24262 47484
rect 24204 47475 24262 47481
rect 25222 47472 25228 47484
rect 25280 47472 25286 47524
rect 15746 47444 15752 47456
rect 15707 47416 15752 47444
rect 15746 47404 15752 47416
rect 15804 47404 15810 47456
rect 27816 47444 27844 47543
rect 27890 47540 27896 47592
rect 27948 47580 27954 47592
rect 28077 47583 28135 47589
rect 27948 47552 27993 47580
rect 27948 47540 27954 47552
rect 28077 47549 28089 47583
rect 28123 47549 28135 47583
rect 29730 47580 29736 47592
rect 29643 47552 29736 47580
rect 28077 47543 28135 47549
rect 27982 47472 27988 47524
rect 28040 47512 28046 47524
rect 28092 47512 28120 47543
rect 29730 47540 29736 47552
rect 29788 47540 29794 47592
rect 30009 47583 30067 47589
rect 30009 47549 30021 47583
rect 30055 47580 30067 47583
rect 30282 47580 30288 47592
rect 30055 47552 30288 47580
rect 30055 47549 30067 47552
rect 30009 47543 30067 47549
rect 30282 47540 30288 47552
rect 30340 47540 30346 47592
rect 30466 47540 30472 47592
rect 30524 47580 30530 47592
rect 30650 47580 30656 47592
rect 30524 47552 30656 47580
rect 30524 47540 30530 47552
rect 30650 47540 30656 47552
rect 30708 47540 30714 47592
rect 33321 47583 33379 47589
rect 33321 47549 33333 47583
rect 33367 47549 33379 47583
rect 33502 47580 33508 47592
rect 33463 47552 33508 47580
rect 33321 47543 33379 47549
rect 28040 47484 28120 47512
rect 30920 47515 30978 47521
rect 28040 47472 28046 47484
rect 30920 47481 30932 47515
rect 30966 47512 30978 47515
rect 31018 47512 31024 47524
rect 30966 47484 31024 47512
rect 30966 47481 30978 47484
rect 30920 47475 30978 47481
rect 31018 47472 31024 47484
rect 31076 47472 31082 47524
rect 33336 47512 33364 47543
rect 33502 47540 33508 47552
rect 33560 47540 33566 47592
rect 33597 47583 33655 47589
rect 33597 47549 33609 47583
rect 33643 47580 33655 47583
rect 34330 47580 34336 47592
rect 33643 47552 34336 47580
rect 33643 47549 33655 47552
rect 33597 47543 33655 47549
rect 34330 47540 34336 47552
rect 34388 47540 34394 47592
rect 57425 47583 57483 47589
rect 57425 47549 57437 47583
rect 57471 47580 57483 47583
rect 57514 47580 57520 47592
rect 57471 47552 57520 47580
rect 57471 47549 57483 47552
rect 57425 47543 57483 47549
rect 57514 47540 57520 47552
rect 57572 47580 57578 47592
rect 57698 47580 57704 47592
rect 57572 47552 57704 47580
rect 57572 47540 57578 47552
rect 57698 47540 57704 47552
rect 57756 47540 57762 47592
rect 33686 47512 33692 47524
rect 33336 47484 33692 47512
rect 33686 47472 33692 47484
rect 33744 47512 33750 47524
rect 34238 47512 34244 47524
rect 33744 47484 34244 47512
rect 33744 47472 33750 47484
rect 34238 47472 34244 47484
rect 34296 47472 34302 47524
rect 55674 47472 55680 47524
rect 55732 47512 55738 47524
rect 57977 47515 58035 47521
rect 57977 47512 57989 47515
rect 55732 47484 57989 47512
rect 55732 47472 55738 47484
rect 57977 47481 57989 47484
rect 58023 47481 58035 47515
rect 58158 47512 58164 47524
rect 58119 47484 58164 47512
rect 57977 47475 58035 47481
rect 58158 47472 58164 47484
rect 58216 47472 58222 47524
rect 28442 47444 28448 47456
rect 27816 47416 28448 47444
rect 28442 47404 28448 47416
rect 28500 47404 28506 47456
rect 29546 47444 29552 47456
rect 29507 47416 29552 47444
rect 29546 47404 29552 47416
rect 29604 47404 29610 47456
rect 32030 47444 32036 47456
rect 31991 47416 32036 47444
rect 32030 47404 32036 47416
rect 32088 47404 32094 47456
rect 33134 47444 33140 47456
rect 33095 47416 33140 47444
rect 33134 47404 33140 47416
rect 33192 47404 33198 47456
rect 1104 47354 58880 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 50326 47354
rect 50378 47302 50390 47354
rect 50442 47302 50454 47354
rect 50506 47302 50518 47354
rect 50570 47302 58880 47354
rect 1104 47280 58880 47302
rect 15746 47200 15752 47252
rect 15804 47240 15810 47252
rect 16301 47243 16359 47249
rect 16301 47240 16313 47243
rect 15804 47212 16313 47240
rect 15804 47200 15810 47212
rect 16301 47209 16313 47212
rect 16347 47209 16359 47243
rect 24210 47240 24216 47252
rect 24171 47212 24216 47240
rect 16301 47203 16359 47209
rect 24210 47200 24216 47212
rect 24268 47200 24274 47252
rect 25222 47240 25228 47252
rect 25183 47212 25228 47240
rect 25222 47200 25228 47212
rect 25280 47200 25286 47252
rect 28261 47243 28319 47249
rect 28261 47209 28273 47243
rect 28307 47240 28319 47243
rect 28350 47240 28356 47252
rect 28307 47212 28356 47240
rect 28307 47209 28319 47212
rect 28261 47203 28319 47209
rect 28350 47200 28356 47212
rect 28408 47200 28414 47252
rect 29549 47243 29607 47249
rect 29549 47209 29561 47243
rect 29595 47240 29607 47243
rect 29730 47240 29736 47252
rect 29595 47212 29736 47240
rect 29595 47209 29607 47212
rect 29549 47203 29607 47209
rect 29730 47200 29736 47212
rect 29788 47200 29794 47252
rect 31018 47240 31024 47252
rect 30979 47212 31024 47240
rect 31018 47200 31024 47212
rect 31076 47200 31082 47252
rect 33502 47200 33508 47252
rect 33560 47240 33566 47252
rect 33689 47243 33747 47249
rect 33689 47240 33701 47243
rect 33560 47212 33701 47240
rect 33560 47200 33566 47212
rect 33689 47209 33701 47212
rect 33735 47209 33747 47243
rect 34238 47240 34244 47252
rect 34199 47212 34244 47240
rect 33689 47203 33747 47209
rect 16117 47175 16175 47181
rect 16117 47141 16129 47175
rect 16163 47172 16175 47175
rect 16482 47172 16488 47184
rect 16163 47144 16488 47172
rect 16163 47141 16175 47144
rect 16117 47135 16175 47141
rect 16482 47132 16488 47144
rect 16540 47132 16546 47184
rect 14921 47107 14979 47113
rect 14921 47073 14933 47107
rect 14967 47104 14979 47107
rect 15378 47104 15384 47116
rect 14967 47076 15384 47104
rect 14967 47073 14979 47076
rect 14921 47067 14979 47073
rect 15378 47064 15384 47076
rect 15436 47064 15442 47116
rect 16390 47104 16396 47116
rect 16351 47076 16396 47104
rect 16390 47064 16396 47076
rect 16448 47064 16454 47116
rect 16853 47107 16911 47113
rect 16853 47073 16865 47107
rect 16899 47073 16911 47107
rect 17034 47104 17040 47116
rect 16995 47076 17040 47104
rect 16853 47067 16911 47073
rect 15197 47039 15255 47045
rect 15197 47005 15209 47039
rect 15243 47036 15255 47039
rect 15286 47036 15292 47048
rect 15243 47008 15292 47036
rect 15243 47005 15255 47008
rect 15197 46999 15255 47005
rect 15286 46996 15292 47008
rect 15344 46996 15350 47048
rect 16868 47036 16896 47067
rect 17034 47064 17040 47076
rect 17092 47064 17098 47116
rect 18782 47104 18788 47116
rect 18743 47076 18788 47104
rect 18782 47064 18788 47076
rect 18840 47064 18846 47116
rect 18969 47107 19027 47113
rect 18969 47073 18981 47107
rect 19015 47104 19027 47107
rect 19150 47104 19156 47116
rect 19015 47076 19156 47104
rect 19015 47073 19027 47076
rect 18969 47067 19027 47073
rect 19150 47064 19156 47076
rect 19208 47064 19214 47116
rect 19981 47107 20039 47113
rect 19981 47073 19993 47107
rect 20027 47104 20039 47107
rect 20162 47104 20168 47116
rect 20027 47076 20168 47104
rect 20027 47073 20039 47076
rect 19981 47067 20039 47073
rect 17954 47036 17960 47048
rect 16868 47008 17960 47036
rect 17954 46996 17960 47008
rect 18012 46996 18018 47048
rect 19061 47039 19119 47045
rect 19061 47005 19073 47039
rect 19107 47036 19119 47039
rect 19334 47036 19340 47048
rect 19107 47008 19340 47036
rect 19107 47005 19119 47008
rect 19061 46999 19119 47005
rect 19334 46996 19340 47008
rect 19392 47036 19398 47048
rect 19996 47036 20024 47067
rect 20162 47064 20168 47076
rect 20220 47064 20226 47116
rect 21168 47107 21226 47113
rect 21168 47073 21180 47107
rect 21214 47104 21226 47107
rect 21450 47104 21456 47116
rect 21214 47076 21456 47104
rect 21214 47073 21226 47076
rect 21168 47067 21226 47073
rect 21450 47064 21456 47076
rect 21508 47064 21514 47116
rect 22925 47107 22983 47113
rect 22925 47073 22937 47107
rect 22971 47104 22983 47107
rect 23474 47104 23480 47116
rect 22971 47076 23480 47104
rect 22971 47073 22983 47076
rect 22925 47067 22983 47073
rect 23474 47064 23480 47076
rect 23532 47064 23538 47116
rect 23661 47107 23719 47113
rect 23661 47073 23673 47107
rect 23707 47073 23719 47107
rect 23661 47067 23719 47073
rect 24121 47107 24179 47113
rect 24121 47073 24133 47107
rect 24167 47073 24179 47107
rect 24121 47067 24179 47073
rect 19392 47008 20024 47036
rect 19392 46996 19398 47008
rect 20622 46996 20628 47048
rect 20680 47036 20686 47048
rect 20901 47039 20959 47045
rect 20901 47036 20913 47039
rect 20680 47008 20913 47036
rect 20680 46996 20686 47008
rect 20901 47005 20913 47008
rect 20947 47005 20959 47039
rect 23676 47036 23704 47067
rect 20901 46999 20959 47005
rect 22756 47008 23704 47036
rect 22756 46980 22784 47008
rect 16114 46968 16120 46980
rect 16075 46940 16120 46968
rect 16114 46928 16120 46940
rect 16172 46928 16178 46980
rect 22738 46968 22744 46980
rect 22699 46940 22744 46968
rect 22738 46928 22744 46940
rect 22796 46928 22802 46980
rect 23474 46968 23480 46980
rect 23435 46940 23480 46968
rect 23474 46928 23480 46940
rect 23532 46928 23538 46980
rect 24136 46968 24164 47067
rect 24228 47036 24256 47200
rect 25314 47132 25320 47184
rect 25372 47172 25378 47184
rect 29914 47172 29920 47184
rect 25372 47144 25728 47172
rect 25372 47132 25378 47144
rect 25406 47104 25412 47116
rect 25367 47076 25412 47104
rect 25406 47064 25412 47076
rect 25464 47064 25470 47116
rect 25700 47113 25728 47144
rect 29380 47144 29920 47172
rect 25685 47107 25743 47113
rect 25685 47073 25697 47107
rect 25731 47073 25743 47107
rect 25685 47067 25743 47073
rect 26694 47064 26700 47116
rect 26752 47104 26758 47116
rect 26789 47107 26847 47113
rect 26789 47104 26801 47107
rect 26752 47076 26801 47104
rect 26752 47064 26758 47076
rect 26789 47073 26801 47076
rect 26835 47073 26847 47107
rect 26789 47067 26847 47073
rect 27801 47107 27859 47113
rect 27801 47073 27813 47107
rect 27847 47073 27859 47107
rect 27801 47067 27859 47073
rect 25593 47039 25651 47045
rect 25593 47036 25605 47039
rect 24228 47008 25605 47036
rect 25593 47005 25605 47008
rect 25639 47005 25651 47039
rect 25593 46999 25651 47005
rect 27065 47039 27123 47045
rect 27065 47005 27077 47039
rect 27111 47036 27123 47039
rect 27614 47036 27620 47048
rect 27111 47008 27620 47036
rect 27111 47005 27123 47008
rect 27065 46999 27123 47005
rect 27614 46996 27620 47008
rect 27672 46996 27678 47048
rect 27816 47036 27844 47067
rect 27890 47064 27896 47116
rect 27948 47104 27954 47116
rect 27985 47107 28043 47113
rect 27985 47104 27997 47107
rect 27948 47076 27997 47104
rect 27948 47064 27954 47076
rect 27985 47073 27997 47076
rect 28031 47073 28043 47107
rect 28258 47104 28264 47116
rect 28219 47076 28264 47104
rect 27985 47067 28043 47073
rect 28258 47064 28264 47076
rect 28316 47064 28322 47116
rect 28442 47104 28448 47116
rect 28403 47076 28448 47104
rect 28442 47064 28448 47076
rect 28500 47064 28506 47116
rect 29380 47113 29408 47144
rect 29914 47132 29920 47144
rect 29972 47132 29978 47184
rect 30466 47132 30472 47184
rect 30524 47172 30530 47184
rect 32576 47175 32634 47181
rect 30524 47144 32352 47172
rect 30524 47132 30530 47144
rect 29365 47107 29423 47113
rect 29365 47073 29377 47107
rect 29411 47073 29423 47107
rect 29365 47067 29423 47073
rect 29549 47107 29607 47113
rect 29549 47073 29561 47107
rect 29595 47104 29607 47107
rect 30282 47104 30288 47116
rect 29595 47076 30288 47104
rect 29595 47073 29607 47076
rect 29549 47067 29607 47073
rect 30282 47064 30288 47076
rect 30340 47064 30346 47116
rect 31205 47107 31263 47113
rect 31205 47073 31217 47107
rect 31251 47073 31263 47107
rect 31205 47067 31263 47073
rect 31481 47107 31539 47113
rect 31481 47073 31493 47107
rect 31527 47104 31539 47107
rect 32030 47104 32036 47116
rect 31527 47076 32036 47104
rect 31527 47073 31539 47076
rect 31481 47067 31539 47073
rect 31220 47036 31248 47067
rect 32030 47064 32036 47076
rect 32088 47064 32094 47116
rect 32324 47048 32352 47144
rect 32576 47141 32588 47175
rect 32622 47172 32634 47175
rect 33134 47172 33140 47184
rect 32622 47144 33140 47172
rect 32622 47141 32634 47144
rect 32576 47135 32634 47141
rect 33134 47132 33140 47144
rect 33192 47132 33198 47184
rect 33704 47104 33732 47203
rect 34238 47200 34244 47212
rect 34296 47200 34302 47252
rect 57698 47240 57704 47252
rect 57659 47212 57704 47240
rect 57698 47200 57704 47212
rect 57756 47200 57762 47252
rect 34149 47107 34207 47113
rect 34149 47104 34161 47107
rect 33704 47076 34161 47104
rect 34149 47073 34161 47076
rect 34195 47073 34207 47107
rect 34330 47104 34336 47116
rect 34291 47076 34336 47104
rect 34149 47067 34207 47073
rect 34330 47064 34336 47076
rect 34388 47064 34394 47116
rect 56870 47104 56876 47116
rect 56831 47076 56876 47104
rect 56870 47064 56876 47076
rect 56928 47064 56934 47116
rect 57517 47107 57575 47113
rect 57517 47073 57529 47107
rect 57563 47104 57575 47107
rect 57606 47104 57612 47116
rect 57563 47076 57612 47104
rect 57563 47073 57575 47076
rect 57517 47067 57575 47073
rect 57606 47064 57612 47076
rect 57664 47064 57670 47116
rect 31846 47036 31852 47048
rect 27816 47008 28028 47036
rect 31220 47008 31852 47036
rect 28000 46980 28028 47008
rect 31846 46996 31852 47008
rect 31904 46996 31910 47048
rect 32306 47036 32312 47048
rect 32267 47008 32312 47036
rect 32306 46996 32312 47008
rect 32364 46996 32370 47048
rect 24762 46968 24768 46980
rect 24136 46940 24768 46968
rect 24762 46928 24768 46940
rect 24820 46928 24826 46980
rect 26973 46971 27031 46977
rect 26973 46937 26985 46971
rect 27019 46968 27031 46971
rect 27798 46968 27804 46980
rect 27019 46940 27804 46968
rect 27019 46937 27031 46940
rect 26973 46931 27031 46937
rect 27798 46928 27804 46940
rect 27856 46928 27862 46980
rect 27982 46928 27988 46980
rect 28040 46928 28046 46980
rect 31389 46971 31447 46977
rect 31389 46937 31401 46971
rect 31435 46968 31447 46971
rect 31938 46968 31944 46980
rect 31435 46940 31944 46968
rect 31435 46937 31447 46940
rect 31389 46931 31447 46937
rect 31938 46928 31944 46940
rect 31996 46928 32002 46980
rect 14734 46900 14740 46912
rect 14695 46872 14740 46900
rect 14734 46860 14740 46872
rect 14792 46860 14798 46912
rect 15102 46900 15108 46912
rect 15063 46872 15108 46900
rect 15102 46860 15108 46872
rect 15160 46860 15166 46912
rect 16945 46903 17003 46909
rect 16945 46869 16957 46903
rect 16991 46900 17003 46903
rect 17770 46900 17776 46912
rect 16991 46872 17776 46900
rect 16991 46869 17003 46872
rect 16945 46863 17003 46869
rect 17770 46860 17776 46872
rect 17828 46860 17834 46912
rect 18598 46900 18604 46912
rect 18559 46872 18604 46900
rect 18598 46860 18604 46872
rect 18656 46860 18662 46912
rect 20070 46900 20076 46912
rect 20031 46872 20076 46900
rect 20070 46860 20076 46872
rect 20128 46860 20134 46912
rect 22281 46903 22339 46909
rect 22281 46869 22293 46903
rect 22327 46900 22339 46903
rect 22554 46900 22560 46912
rect 22327 46872 22560 46900
rect 22327 46869 22339 46872
rect 22281 46863 22339 46869
rect 22554 46860 22560 46872
rect 22612 46860 22618 46912
rect 26602 46900 26608 46912
rect 26563 46872 26608 46900
rect 26602 46860 26608 46872
rect 26660 46860 26666 46912
rect 1104 46810 58880 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 58880 46810
rect 1104 46736 58880 46758
rect 14829 46699 14887 46705
rect 14829 46665 14841 46699
rect 14875 46696 14887 46699
rect 15102 46696 15108 46708
rect 14875 46668 15108 46696
rect 14875 46665 14887 46668
rect 14829 46659 14887 46665
rect 15102 46656 15108 46668
rect 15160 46656 15166 46708
rect 15378 46696 15384 46708
rect 15339 46668 15384 46696
rect 15378 46656 15384 46668
rect 15436 46656 15442 46708
rect 16025 46699 16083 46705
rect 16025 46665 16037 46699
rect 16071 46696 16083 46699
rect 16390 46696 16396 46708
rect 16071 46668 16396 46696
rect 16071 46665 16083 46668
rect 16025 46659 16083 46665
rect 16390 46656 16396 46668
rect 16448 46656 16454 46708
rect 18969 46699 19027 46705
rect 18969 46665 18981 46699
rect 19015 46696 19027 46699
rect 19150 46696 19156 46708
rect 19015 46668 19156 46696
rect 19015 46665 19027 46668
rect 18969 46659 19027 46665
rect 19150 46656 19156 46668
rect 19208 46656 19214 46708
rect 20162 46656 20168 46708
rect 20220 46696 20226 46708
rect 20809 46699 20867 46705
rect 20809 46696 20821 46699
rect 20220 46668 20821 46696
rect 20220 46656 20226 46668
rect 20809 46665 20821 46668
rect 20855 46665 20867 46699
rect 20809 46659 20867 46665
rect 22462 46656 22468 46708
rect 22520 46696 22526 46708
rect 22741 46699 22799 46705
rect 22741 46696 22753 46699
rect 22520 46668 22753 46696
rect 22520 46656 22526 46668
rect 22741 46665 22753 46668
rect 22787 46665 22799 46699
rect 27798 46696 27804 46708
rect 27759 46668 27804 46696
rect 22741 46659 22799 46665
rect 27798 46656 27804 46668
rect 27856 46656 27862 46708
rect 30282 46696 30288 46708
rect 30243 46668 30288 46696
rect 30282 46656 30288 46668
rect 30340 46656 30346 46708
rect 31846 46656 31852 46708
rect 31904 46696 31910 46708
rect 32033 46699 32091 46705
rect 32033 46696 32045 46699
rect 31904 46668 32045 46696
rect 31904 46656 31910 46668
rect 32033 46665 32045 46668
rect 32079 46665 32091 46699
rect 32033 46659 32091 46665
rect 15396 46560 15424 46656
rect 31205 46631 31263 46637
rect 31205 46597 31217 46631
rect 31251 46628 31263 46631
rect 32398 46628 32404 46640
rect 31251 46600 32404 46628
rect 31251 46597 31263 46600
rect 31205 46591 31263 46597
rect 32398 46588 32404 46600
rect 32456 46588 32462 46640
rect 19426 46560 19432 46572
rect 15396 46532 15976 46560
rect 19387 46532 19432 46560
rect 1394 46492 1400 46504
rect 1355 46464 1400 46492
rect 1394 46452 1400 46464
rect 1452 46452 1458 46504
rect 13449 46495 13507 46501
rect 13449 46461 13461 46495
rect 13495 46461 13507 46495
rect 13449 46455 13507 46461
rect 13716 46495 13774 46501
rect 13716 46461 13728 46495
rect 13762 46492 13774 46495
rect 14734 46492 14740 46504
rect 13762 46464 14740 46492
rect 13762 46461 13774 46464
rect 13716 46455 13774 46461
rect 13464 46424 13492 46455
rect 14734 46452 14740 46464
rect 14792 46452 14798 46504
rect 15102 46452 15108 46504
rect 15160 46492 15166 46504
rect 15289 46495 15347 46501
rect 15289 46492 15301 46495
rect 15160 46464 15301 46492
rect 15160 46452 15166 46464
rect 15289 46461 15301 46464
rect 15335 46461 15347 46495
rect 15289 46455 15347 46461
rect 15378 46452 15384 46504
rect 15436 46492 15442 46504
rect 15948 46501 15976 46532
rect 19426 46520 19432 46532
rect 19484 46520 19490 46572
rect 24670 46520 24676 46572
rect 24728 46560 24734 46572
rect 25501 46563 25559 46569
rect 25501 46560 25513 46563
rect 24728 46532 25513 46560
rect 24728 46520 24734 46532
rect 25501 46529 25513 46532
rect 25547 46529 25559 46563
rect 31754 46560 31760 46572
rect 25501 46523 25559 46529
rect 30300 46532 31760 46560
rect 15473 46495 15531 46501
rect 15473 46492 15485 46495
rect 15436 46464 15485 46492
rect 15436 46452 15442 46464
rect 15473 46461 15485 46464
rect 15519 46461 15531 46495
rect 15473 46455 15531 46461
rect 15933 46495 15991 46501
rect 15933 46461 15945 46495
rect 15979 46461 15991 46495
rect 15933 46455 15991 46461
rect 16758 46452 16764 46504
rect 16816 46492 16822 46504
rect 17589 46495 17647 46501
rect 17589 46492 17601 46495
rect 16816 46464 17601 46492
rect 16816 46452 16822 46464
rect 17589 46461 17601 46464
rect 17635 46461 17647 46495
rect 17589 46455 17647 46461
rect 17856 46495 17914 46501
rect 17856 46461 17868 46495
rect 17902 46492 17914 46495
rect 18598 46492 18604 46504
rect 17902 46464 18604 46492
rect 17902 46461 17914 46464
rect 17856 46455 17914 46461
rect 18598 46452 18604 46464
rect 18656 46452 18662 46504
rect 19696 46495 19754 46501
rect 19696 46461 19708 46495
rect 19742 46492 19754 46495
rect 20070 46492 20076 46504
rect 19742 46464 20076 46492
rect 19742 46461 19754 46464
rect 19696 46455 19754 46461
rect 20070 46452 20076 46464
rect 20128 46452 20134 46504
rect 20898 46452 20904 46504
rect 20956 46492 20962 46504
rect 21453 46495 21511 46501
rect 21453 46492 21465 46495
rect 20956 46464 21465 46492
rect 20956 46452 20962 46464
rect 21453 46461 21465 46464
rect 21499 46461 21511 46495
rect 23382 46492 23388 46504
rect 23343 46464 23388 46492
rect 21453 46455 21511 46461
rect 23382 46452 23388 46464
rect 23440 46452 23446 46504
rect 23569 46495 23627 46501
rect 23569 46461 23581 46495
rect 23615 46461 23627 46495
rect 24762 46492 24768 46504
rect 24723 46464 24768 46492
rect 23569 46455 23627 46461
rect 13906 46424 13912 46436
rect 13464 46396 13912 46424
rect 13906 46384 13912 46396
rect 13964 46384 13970 46436
rect 22554 46424 22560 46436
rect 22515 46396 22560 46424
rect 22554 46384 22560 46396
rect 22612 46384 22618 46436
rect 22830 46433 22836 46436
rect 22773 46427 22836 46433
rect 22773 46424 22785 46427
rect 22664 46396 22785 46424
rect 21545 46359 21603 46365
rect 21545 46325 21557 46359
rect 21591 46356 21603 46359
rect 22094 46356 22100 46368
rect 21591 46328 22100 46356
rect 21591 46325 21603 46328
rect 21545 46319 21603 46325
rect 22094 46316 22100 46328
rect 22152 46356 22158 46368
rect 22664 46356 22692 46396
rect 22773 46393 22785 46396
rect 22819 46393 22836 46427
rect 22773 46387 22836 46393
rect 22830 46384 22836 46387
rect 22888 46384 22894 46436
rect 23584 46424 23612 46455
rect 24762 46452 24768 46464
rect 24820 46452 24826 46504
rect 24946 46492 24952 46504
rect 24907 46464 24952 46492
rect 24946 46452 24952 46464
rect 25004 46452 25010 46504
rect 25038 46452 25044 46504
rect 25096 46492 25102 46504
rect 25768 46495 25826 46501
rect 25096 46464 25141 46492
rect 25096 46452 25102 46464
rect 25768 46461 25780 46495
rect 25814 46492 25826 46495
rect 26602 46492 26608 46504
rect 25814 46464 26608 46492
rect 25814 46461 25826 46464
rect 25768 46455 25826 46461
rect 26602 46452 26608 46464
rect 26660 46452 26666 46504
rect 27801 46495 27859 46501
rect 27801 46461 27813 46495
rect 27847 46461 27859 46495
rect 27982 46492 27988 46504
rect 27943 46464 27988 46492
rect 27801 46455 27859 46461
rect 22940 46396 23612 46424
rect 27816 46424 27844 46455
rect 27982 46452 27988 46464
rect 28040 46452 28046 46504
rect 28905 46495 28963 46501
rect 28905 46461 28917 46495
rect 28951 46492 28963 46495
rect 30300 46492 30328 46532
rect 31754 46520 31760 46532
rect 31812 46520 31818 46572
rect 32306 46520 32312 46572
rect 32364 46560 32370 46572
rect 33045 46563 33103 46569
rect 33045 46560 33057 46563
rect 32364 46532 33057 46560
rect 32364 46520 32370 46532
rect 33045 46529 33057 46532
rect 33091 46529 33103 46563
rect 58158 46560 58164 46572
rect 58119 46532 58164 46560
rect 33045 46523 33103 46529
rect 58158 46520 58164 46532
rect 58216 46520 58222 46572
rect 31478 46492 31484 46504
rect 28951 46464 30328 46492
rect 31439 46464 31484 46492
rect 28951 46461 28963 46464
rect 28905 46455 28963 46461
rect 31478 46452 31484 46464
rect 31536 46452 31542 46504
rect 31938 46492 31944 46504
rect 31899 46464 31944 46492
rect 31938 46452 31944 46464
rect 31996 46452 32002 46504
rect 32030 46452 32036 46504
rect 32088 46492 32094 46504
rect 32125 46495 32183 46501
rect 32125 46492 32137 46495
rect 32088 46464 32137 46492
rect 32088 46452 32094 46464
rect 32125 46461 32137 46464
rect 32171 46461 32183 46495
rect 32125 46455 32183 46461
rect 28442 46424 28448 46436
rect 27816 46396 28448 46424
rect 22940 46368 22968 46396
rect 28442 46384 28448 46396
rect 28500 46384 28506 46436
rect 29172 46427 29230 46433
rect 29172 46393 29184 46427
rect 29218 46424 29230 46427
rect 29546 46424 29552 46436
rect 29218 46396 29552 46424
rect 29218 46393 29230 46396
rect 29172 46387 29230 46393
rect 29546 46384 29552 46396
rect 29604 46384 29610 46436
rect 31202 46424 31208 46436
rect 31163 46396 31208 46424
rect 31202 46384 31208 46396
rect 31260 46384 31266 46436
rect 33312 46427 33370 46433
rect 33312 46393 33324 46427
rect 33358 46424 33370 46427
rect 33502 46424 33508 46436
rect 33358 46396 33508 46424
rect 33358 46393 33370 46396
rect 33312 46387 33370 46393
rect 33502 46384 33508 46396
rect 33560 46384 33566 46436
rect 57974 46424 57980 46436
rect 57935 46396 57980 46424
rect 57974 46384 57980 46396
rect 58032 46384 58038 46436
rect 22922 46356 22928 46368
rect 22152 46328 22692 46356
rect 22883 46328 22928 46356
rect 22152 46316 22158 46328
rect 22922 46316 22928 46328
rect 22980 46316 22986 46368
rect 23014 46316 23020 46368
rect 23072 46356 23078 46368
rect 23477 46359 23535 46365
rect 23477 46356 23489 46359
rect 23072 46328 23489 46356
rect 23072 46316 23078 46328
rect 23477 46325 23489 46328
rect 23523 46325 23535 46359
rect 24578 46356 24584 46368
rect 24539 46328 24584 46356
rect 23477 46319 23535 46325
rect 24578 46316 24584 46328
rect 24636 46316 24642 46368
rect 26881 46359 26939 46365
rect 26881 46325 26893 46359
rect 26927 46356 26939 46359
rect 27614 46356 27620 46368
rect 26927 46328 27620 46356
rect 26927 46325 26939 46328
rect 26881 46319 26939 46325
rect 27614 46316 27620 46328
rect 27672 46316 27678 46368
rect 31386 46356 31392 46368
rect 31347 46328 31392 46356
rect 31386 46316 31392 46328
rect 31444 46316 31450 46368
rect 33410 46316 33416 46368
rect 33468 46356 33474 46368
rect 34330 46356 34336 46368
rect 33468 46328 34336 46356
rect 33468 46316 33474 46328
rect 34330 46316 34336 46328
rect 34388 46356 34394 46368
rect 34425 46359 34483 46365
rect 34425 46356 34437 46359
rect 34388 46328 34437 46356
rect 34388 46316 34394 46328
rect 34425 46325 34437 46328
rect 34471 46325 34483 46359
rect 34425 46319 34483 46325
rect 1104 46266 58880 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 50326 46266
rect 50378 46214 50390 46266
rect 50442 46214 50454 46266
rect 50506 46214 50518 46266
rect 50570 46214 58880 46266
rect 1104 46192 58880 46214
rect 17034 46112 17040 46164
rect 17092 46152 17098 46164
rect 17129 46155 17187 46161
rect 17129 46152 17141 46155
rect 17092 46124 17141 46152
rect 17092 46112 17098 46124
rect 17129 46121 17141 46124
rect 17175 46121 17187 46155
rect 17129 46115 17187 46121
rect 19426 46112 19432 46164
rect 19484 46152 19490 46164
rect 20622 46152 20628 46164
rect 19484 46124 20628 46152
rect 19484 46112 19490 46124
rect 20622 46112 20628 46124
rect 20680 46112 20686 46164
rect 21450 46152 21456 46164
rect 21411 46124 21456 46152
rect 21450 46112 21456 46124
rect 21508 46112 21514 46164
rect 21637 46155 21695 46161
rect 21637 46121 21649 46155
rect 21683 46152 21695 46155
rect 22094 46152 22100 46164
rect 21683 46124 22100 46152
rect 21683 46121 21695 46124
rect 21637 46115 21695 46121
rect 22094 46112 22100 46124
rect 22152 46112 22158 46164
rect 25038 46112 25044 46164
rect 25096 46152 25102 46164
rect 26605 46155 26663 46161
rect 26605 46152 26617 46155
rect 25096 46124 26617 46152
rect 25096 46112 25102 46124
rect 26605 46121 26617 46124
rect 26651 46121 26663 46155
rect 26605 46115 26663 46121
rect 30469 46155 30527 46161
rect 30469 46121 30481 46155
rect 30515 46121 30527 46155
rect 30469 46115 30527 46121
rect 22738 46084 22744 46096
rect 20824 46056 22744 46084
rect 14737 46019 14795 46025
rect 14737 45985 14749 46019
rect 14783 46016 14795 46019
rect 15378 46016 15384 46028
rect 14783 45988 15384 46016
rect 14783 45985 14795 45988
rect 14737 45979 14795 45985
rect 15378 45976 15384 45988
rect 15436 45976 15442 46028
rect 16016 46019 16074 46025
rect 16016 45985 16028 46019
rect 16062 46016 16074 46019
rect 17589 46019 17647 46025
rect 17589 46016 17601 46019
rect 16062 45988 17601 46016
rect 16062 45985 16074 45988
rect 16016 45979 16074 45985
rect 17589 45985 17601 45988
rect 17635 45985 17647 46019
rect 17770 46016 17776 46028
rect 17731 45988 17776 46016
rect 17589 45979 17647 45985
rect 17770 45976 17776 45988
rect 17828 46016 17834 46028
rect 18509 46019 18567 46025
rect 18509 46016 18521 46019
rect 17828 45988 18521 46016
rect 17828 45976 17834 45988
rect 18509 45985 18521 45988
rect 18555 45985 18567 46019
rect 18509 45979 18567 45985
rect 19886 45976 19892 46028
rect 19944 46016 19950 46028
rect 19981 46019 20039 46025
rect 19981 46016 19993 46019
rect 19944 45988 19993 46016
rect 19944 45976 19950 45988
rect 19981 45985 19993 45988
rect 20027 45985 20039 46019
rect 20162 46016 20168 46028
rect 20123 45988 20168 46016
rect 19981 45979 20039 45985
rect 20162 45976 20168 45988
rect 20220 45976 20226 46028
rect 20824 46025 20852 46056
rect 22738 46044 22744 46056
rect 22796 46044 22802 46096
rect 23014 46093 23020 46096
rect 23008 46084 23020 46093
rect 22975 46056 23020 46084
rect 23008 46047 23020 46056
rect 23014 46044 23020 46047
rect 23072 46044 23078 46096
rect 24578 46044 24584 46096
rect 24636 46084 24642 46096
rect 25470 46087 25528 46093
rect 25470 46084 25482 46087
rect 24636 46056 25482 46084
rect 24636 46044 24642 46056
rect 25470 46053 25482 46056
rect 25516 46053 25528 46087
rect 26620 46084 26648 46115
rect 29270 46084 29276 46096
rect 26620 46056 27292 46084
rect 25470 46047 25528 46053
rect 20809 46019 20867 46025
rect 20809 45985 20821 46019
rect 20855 45985 20867 46019
rect 20809 45979 20867 45985
rect 21634 46019 21692 46025
rect 21634 45985 21646 46019
rect 21680 46016 21692 46019
rect 22097 46019 22155 46025
rect 22097 46016 22109 46019
rect 21680 45988 22109 46016
rect 21680 45985 21692 45988
rect 21634 45979 21692 45985
rect 22097 45985 22109 45988
rect 22143 46016 22155 46019
rect 22554 46016 22560 46028
rect 22143 45988 22560 46016
rect 22143 45985 22155 45988
rect 22097 45979 22155 45985
rect 22554 45976 22560 45988
rect 22612 45976 22618 46028
rect 23474 46016 23480 46028
rect 22756 45988 23480 46016
rect 13906 45908 13912 45960
rect 13964 45948 13970 45960
rect 15749 45951 15807 45957
rect 15749 45948 15761 45951
rect 13964 45920 15761 45948
rect 13964 45908 13970 45920
rect 15749 45917 15761 45920
rect 15795 45917 15807 45951
rect 15749 45911 15807 45917
rect 17034 45908 17040 45960
rect 17092 45948 17098 45960
rect 22756 45957 22784 45988
rect 23474 45976 23480 45988
rect 23532 46016 23538 46028
rect 23532 45988 23796 46016
rect 23532 45976 23538 45988
rect 18049 45951 18107 45957
rect 18049 45948 18061 45951
rect 17092 45920 18061 45948
rect 17092 45908 17098 45920
rect 18049 45917 18061 45920
rect 18095 45917 18107 45951
rect 18049 45911 18107 45917
rect 22005 45951 22063 45957
rect 22005 45917 22017 45951
rect 22051 45948 22063 45951
rect 22741 45951 22799 45957
rect 22051 45920 22140 45948
rect 22051 45917 22063 45920
rect 22005 45911 22063 45917
rect 22112 45892 22140 45920
rect 22741 45917 22753 45951
rect 22787 45917 22799 45951
rect 23768 45948 23796 45988
rect 24946 45976 24952 46028
rect 25004 46016 25010 46028
rect 27264 46025 27292 46056
rect 27724 46056 29276 46084
rect 27065 46019 27123 46025
rect 27065 46016 27077 46019
rect 25004 45988 27077 46016
rect 25004 45976 25010 45988
rect 27065 45985 27077 45988
rect 27111 45985 27123 46019
rect 27065 45979 27123 45985
rect 27249 46019 27307 46025
rect 27249 45985 27261 46019
rect 27295 45985 27307 46019
rect 27249 45979 27307 45985
rect 27430 45976 27436 46028
rect 27488 46016 27494 46028
rect 27724 46025 27752 46056
rect 29270 46044 29276 46056
rect 29328 46044 29334 46096
rect 30484 46084 30512 46115
rect 31202 46112 31208 46164
rect 31260 46152 31266 46164
rect 32493 46155 32551 46161
rect 32493 46152 32505 46155
rect 31260 46124 32505 46152
rect 31260 46112 31266 46124
rect 32493 46121 32505 46124
rect 32539 46121 32551 46155
rect 33502 46152 33508 46164
rect 33463 46124 33508 46152
rect 32493 46115 32551 46121
rect 33502 46112 33508 46124
rect 33560 46112 33566 46164
rect 57974 46112 57980 46164
rect 58032 46152 58038 46164
rect 58161 46155 58219 46161
rect 58161 46152 58173 46155
rect 58032 46124 58173 46152
rect 58032 46112 58038 46124
rect 58161 46121 58173 46124
rect 58207 46121 58219 46155
rect 58161 46115 58219 46121
rect 33042 46084 33048 46096
rect 30484 46056 33048 46084
rect 33042 46044 33048 46056
rect 33100 46044 33106 46096
rect 27709 46019 27767 46025
rect 27709 46016 27721 46019
rect 27488 45988 27721 46016
rect 27488 45976 27494 45988
rect 27709 45985 27721 45988
rect 27755 45985 27767 46019
rect 27709 45979 27767 45985
rect 27798 45976 27804 46028
rect 27856 46016 27862 46028
rect 27965 46019 28023 46025
rect 27965 46016 27977 46019
rect 27856 45988 27977 46016
rect 27856 45976 27862 45988
rect 27965 45985 27977 45988
rect 28011 45985 28023 46019
rect 29288 46016 29316 46044
rect 30466 46016 30472 46028
rect 29288 45988 30472 46016
rect 27965 45979 28023 45985
rect 30466 45976 30472 45988
rect 30524 45976 30530 46028
rect 30650 46016 30656 46028
rect 30611 45988 30656 46016
rect 30650 45976 30656 45988
rect 30708 45976 30714 46028
rect 31380 46019 31438 46025
rect 31380 45985 31392 46019
rect 31426 46016 31438 46019
rect 32950 46016 32956 46028
rect 31426 45988 32956 46016
rect 31426 45985 31438 45988
rect 31380 45979 31438 45985
rect 32950 45976 32956 45988
rect 33008 45976 33014 46028
rect 33410 46016 33416 46028
rect 33371 45988 33416 46016
rect 33410 45976 33416 45988
rect 33468 45976 33474 46028
rect 24670 45948 24676 45960
rect 23768 45920 24676 45948
rect 22741 45911 22799 45917
rect 17954 45880 17960 45892
rect 17915 45852 17960 45880
rect 17954 45840 17960 45852
rect 18012 45840 18018 45892
rect 22094 45840 22100 45892
rect 22152 45840 22158 45892
rect 22554 45840 22560 45892
rect 22612 45880 22618 45892
rect 22756 45880 22784 45911
rect 24670 45908 24676 45920
rect 24728 45948 24734 45960
rect 25225 45951 25283 45957
rect 25225 45948 25237 45951
rect 24728 45920 25237 45948
rect 24728 45908 24734 45920
rect 25225 45917 25237 45920
rect 25271 45917 25283 45951
rect 30484 45948 30512 45976
rect 31113 45951 31171 45957
rect 31113 45948 31125 45951
rect 30484 45920 31125 45948
rect 25225 45911 25283 45917
rect 31113 45917 31125 45920
rect 31159 45917 31171 45951
rect 31113 45911 31171 45917
rect 57057 45951 57115 45957
rect 57057 45917 57069 45951
rect 57103 45948 57115 45951
rect 57517 45951 57575 45957
rect 57517 45948 57529 45951
rect 57103 45920 57529 45948
rect 57103 45917 57115 45920
rect 57057 45911 57115 45917
rect 57517 45917 57529 45920
rect 57563 45917 57575 45951
rect 57698 45948 57704 45960
rect 57659 45920 57704 45948
rect 57517 45911 57575 45917
rect 57698 45908 57704 45920
rect 57756 45908 57762 45960
rect 22612 45852 22784 45880
rect 22612 45840 22618 45852
rect 14826 45812 14832 45824
rect 14787 45784 14832 45812
rect 14826 45772 14832 45784
rect 14884 45772 14890 45824
rect 18598 45812 18604 45824
rect 18559 45784 18604 45812
rect 18598 45772 18604 45784
rect 18656 45772 18662 45824
rect 20070 45812 20076 45824
rect 20031 45784 20076 45812
rect 20070 45772 20076 45784
rect 20128 45772 20134 45824
rect 22462 45772 22468 45824
rect 22520 45812 22526 45824
rect 24121 45815 24179 45821
rect 24121 45812 24133 45815
rect 22520 45784 24133 45812
rect 22520 45772 22526 45784
rect 24121 45781 24133 45784
rect 24167 45781 24179 45815
rect 24121 45775 24179 45781
rect 24762 45772 24768 45824
rect 24820 45812 24826 45824
rect 27157 45815 27215 45821
rect 27157 45812 27169 45815
rect 24820 45784 27169 45812
rect 24820 45772 24826 45784
rect 27157 45781 27169 45784
rect 27203 45781 27215 45815
rect 29086 45812 29092 45824
rect 29047 45784 29092 45812
rect 27157 45775 27215 45781
rect 29086 45772 29092 45784
rect 29144 45772 29150 45824
rect 1104 45722 58880 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 58880 45722
rect 1104 45648 58880 45670
rect 15378 45608 15384 45620
rect 15339 45580 15384 45608
rect 15378 45568 15384 45580
rect 15436 45568 15442 45620
rect 22557 45611 22615 45617
rect 22557 45577 22569 45611
rect 22603 45608 22615 45611
rect 23382 45608 23388 45620
rect 22603 45580 23388 45608
rect 22603 45577 22615 45580
rect 22557 45571 22615 45577
rect 23382 45568 23388 45580
rect 23440 45568 23446 45620
rect 24946 45568 24952 45620
rect 25004 45608 25010 45620
rect 25133 45611 25191 45617
rect 25133 45608 25145 45611
rect 25004 45580 25145 45608
rect 25004 45568 25010 45580
rect 25133 45577 25145 45580
rect 25179 45577 25191 45611
rect 27798 45608 27804 45620
rect 27759 45580 27804 45608
rect 25133 45571 25191 45577
rect 27798 45568 27804 45580
rect 27856 45568 27862 45620
rect 31202 45568 31208 45620
rect 31260 45608 31266 45620
rect 31481 45611 31539 45617
rect 31481 45608 31493 45611
rect 31260 45580 31493 45608
rect 31260 45568 31266 45580
rect 31481 45577 31493 45580
rect 31527 45577 31539 45611
rect 31481 45571 31539 45577
rect 57241 45611 57299 45617
rect 57241 45577 57253 45611
rect 57287 45608 57299 45611
rect 57698 45608 57704 45620
rect 57287 45580 57704 45608
rect 57287 45577 57299 45580
rect 57241 45571 57299 45577
rect 57698 45568 57704 45580
rect 57756 45568 57762 45620
rect 17773 45543 17831 45549
rect 17773 45509 17785 45543
rect 17819 45540 17831 45543
rect 17954 45540 17960 45552
rect 17819 45512 17960 45540
rect 17819 45509 17831 45512
rect 17773 45503 17831 45509
rect 17954 45500 17960 45512
rect 18012 45540 18018 45552
rect 18598 45540 18604 45552
rect 18012 45512 18604 45540
rect 18012 45500 18018 45512
rect 18598 45500 18604 45512
rect 18656 45500 18662 45552
rect 31665 45543 31723 45549
rect 31665 45509 31677 45543
rect 31711 45540 31723 45543
rect 31938 45540 31944 45552
rect 31711 45512 31944 45540
rect 31711 45509 31723 45512
rect 31665 45503 31723 45509
rect 31938 45500 31944 45512
rect 31996 45540 32002 45552
rect 58158 45540 58164 45552
rect 31996 45512 33272 45540
rect 58119 45512 58164 45540
rect 31996 45500 32002 45512
rect 13998 45472 14004 45484
rect 13959 45444 14004 45472
rect 13998 45432 14004 45444
rect 14056 45432 14062 45484
rect 24302 45432 24308 45484
rect 24360 45472 24366 45484
rect 29270 45472 29276 45484
rect 24360 45444 24624 45472
rect 24360 45432 24366 45444
rect 1394 45404 1400 45416
rect 1355 45376 1400 45404
rect 1394 45364 1400 45376
rect 1452 45364 1458 45416
rect 14268 45407 14326 45413
rect 14268 45373 14280 45407
rect 14314 45404 14326 45407
rect 14826 45404 14832 45416
rect 14314 45376 14832 45404
rect 14314 45373 14326 45376
rect 14268 45367 14326 45373
rect 14826 45364 14832 45376
rect 14884 45364 14890 45416
rect 17586 45404 17592 45416
rect 17547 45376 17592 45404
rect 17586 45364 17592 45376
rect 17644 45364 17650 45416
rect 17865 45407 17923 45413
rect 17865 45373 17877 45407
rect 17911 45404 17923 45407
rect 18138 45404 18144 45416
rect 17911 45376 18144 45404
rect 17911 45373 17923 45376
rect 17865 45367 17923 45373
rect 18138 45364 18144 45376
rect 18196 45364 18202 45416
rect 18601 45407 18659 45413
rect 18601 45373 18613 45407
rect 18647 45404 18659 45407
rect 19426 45404 19432 45416
rect 18647 45376 19432 45404
rect 18647 45373 18659 45376
rect 18601 45367 18659 45373
rect 19426 45364 19432 45376
rect 19484 45364 19490 45416
rect 20898 45404 20904 45416
rect 20859 45376 20904 45404
rect 20898 45364 20904 45376
rect 20956 45364 20962 45416
rect 20990 45364 20996 45416
rect 21048 45404 21054 45416
rect 21085 45407 21143 45413
rect 21085 45404 21097 45407
rect 21048 45376 21097 45404
rect 21048 45364 21054 45376
rect 21085 45373 21097 45376
rect 21131 45373 21143 45407
rect 21085 45367 21143 45373
rect 21177 45407 21235 45413
rect 21177 45373 21189 45407
rect 21223 45404 21235 45407
rect 21634 45404 21640 45416
rect 21223 45376 21640 45404
rect 21223 45373 21235 45376
rect 21177 45367 21235 45373
rect 21634 45364 21640 45376
rect 21692 45364 21698 45416
rect 22462 45364 22468 45416
rect 22520 45404 22526 45416
rect 22557 45407 22615 45413
rect 22557 45404 22569 45407
rect 22520 45376 22569 45404
rect 22520 45364 22526 45376
rect 22557 45373 22569 45376
rect 22603 45373 22615 45407
rect 22830 45404 22836 45416
rect 22791 45376 22836 45404
rect 22557 45367 22615 45373
rect 22830 45364 22836 45376
rect 22888 45364 22894 45416
rect 22922 45364 22928 45416
rect 22980 45404 22986 45416
rect 23293 45407 23351 45413
rect 23293 45404 23305 45407
rect 22980 45376 23305 45404
rect 22980 45364 22986 45376
rect 23293 45373 23305 45376
rect 23339 45373 23351 45407
rect 23293 45367 23351 45373
rect 23477 45407 23535 45413
rect 23477 45373 23489 45407
rect 23523 45404 23535 45407
rect 23934 45404 23940 45416
rect 23523 45376 23940 45404
rect 23523 45373 23535 45376
rect 23477 45367 23535 45373
rect 23934 45364 23940 45376
rect 23992 45364 23998 45416
rect 24210 45364 24216 45416
rect 24268 45404 24274 45416
rect 24596 45413 24624 45444
rect 26068 45444 28120 45472
rect 29231 45444 29276 45472
rect 26068 45413 26096 45444
rect 24397 45407 24455 45413
rect 24397 45404 24409 45407
rect 24268 45376 24409 45404
rect 24268 45364 24274 45376
rect 24397 45373 24409 45376
rect 24443 45373 24455 45407
rect 24397 45367 24455 45373
rect 24581 45407 24639 45413
rect 24581 45373 24593 45407
rect 24627 45373 24639 45407
rect 24581 45367 24639 45373
rect 25041 45407 25099 45413
rect 25041 45373 25053 45407
rect 25087 45373 25099 45407
rect 25041 45367 25099 45373
rect 26053 45407 26111 45413
rect 26053 45373 26065 45407
rect 26099 45373 26111 45407
rect 26234 45404 26240 45416
rect 26195 45376 26240 45404
rect 26053 45367 26111 45373
rect 18690 45296 18696 45348
rect 18748 45336 18754 45348
rect 18846 45339 18904 45345
rect 18846 45336 18858 45339
rect 18748 45308 18858 45336
rect 18748 45296 18754 45308
rect 18846 45305 18858 45308
rect 18892 45305 18904 45339
rect 18846 45299 18904 45305
rect 22646 45296 22652 45348
rect 22704 45336 22710 45348
rect 22741 45339 22799 45345
rect 22741 45336 22753 45339
rect 22704 45308 22753 45336
rect 22704 45296 22710 45308
rect 22741 45305 22753 45308
rect 22787 45305 22799 45339
rect 25056 45336 25084 45367
rect 26234 45364 26240 45376
rect 26292 45364 26298 45416
rect 27706 45364 27712 45416
rect 27764 45404 27770 45416
rect 28092 45413 28120 45444
rect 29270 45432 29276 45444
rect 29328 45432 29334 45484
rect 32950 45432 32956 45484
rect 33008 45472 33014 45484
rect 33137 45475 33195 45481
rect 33137 45472 33149 45475
rect 33008 45444 33149 45472
rect 33008 45432 33014 45444
rect 33137 45441 33149 45444
rect 33183 45441 33195 45475
rect 33137 45435 33195 45441
rect 27801 45407 27859 45413
rect 27801 45404 27813 45407
rect 27764 45376 27813 45404
rect 27764 45364 27770 45376
rect 27801 45373 27813 45376
rect 27847 45373 27859 45407
rect 27801 45367 27859 45373
rect 28077 45407 28135 45413
rect 28077 45373 28089 45407
rect 28123 45404 28135 45407
rect 28442 45404 28448 45416
rect 28123 45376 28448 45404
rect 28123 45373 28135 45376
rect 28077 45367 28135 45373
rect 28442 45364 28448 45376
rect 28500 45364 28506 45416
rect 28629 45407 28687 45413
rect 28629 45373 28641 45407
rect 28675 45404 28687 45407
rect 29086 45404 29092 45416
rect 28675 45376 29092 45404
rect 28675 45373 28687 45376
rect 28629 45367 28687 45373
rect 29086 45364 29092 45376
rect 29144 45364 29150 45416
rect 32398 45364 32404 45416
rect 32456 45404 32462 45416
rect 33244 45413 33272 45512
rect 58158 45500 58164 45512
rect 58216 45500 58222 45552
rect 33045 45407 33103 45413
rect 33045 45404 33057 45407
rect 32456 45376 33057 45404
rect 32456 45364 32462 45376
rect 33045 45373 33057 45376
rect 33091 45373 33103 45407
rect 33045 45367 33103 45373
rect 33229 45407 33287 45413
rect 33229 45373 33241 45407
rect 33275 45373 33287 45407
rect 33229 45367 33287 45373
rect 56502 45364 56508 45416
rect 56560 45404 56566 45416
rect 56597 45407 56655 45413
rect 56597 45404 56609 45407
rect 56560 45376 56609 45404
rect 56560 45364 56566 45376
rect 56597 45373 56609 45376
rect 56643 45373 56655 45407
rect 56597 45367 56655 45373
rect 57330 45364 57336 45416
rect 57388 45404 57394 45416
rect 57425 45407 57483 45413
rect 57425 45404 57437 45407
rect 57388 45376 57437 45404
rect 57388 45364 57394 45376
rect 57425 45373 57437 45376
rect 57471 45373 57483 45407
rect 57425 45367 57483 45373
rect 26418 45336 26424 45348
rect 22741 45299 22799 45305
rect 24504 45308 25084 45336
rect 26379 45308 26424 45336
rect 24504 45280 24532 45308
rect 26418 45296 26424 45308
rect 26476 45296 26482 45348
rect 27982 45336 27988 45348
rect 27895 45308 27988 45336
rect 27982 45296 27988 45308
rect 28040 45336 28046 45348
rect 28721 45339 28779 45345
rect 28721 45336 28733 45339
rect 28040 45308 28733 45336
rect 28040 45296 28046 45308
rect 28721 45305 28733 45308
rect 28767 45305 28779 45339
rect 28721 45299 28779 45305
rect 29540 45339 29598 45345
rect 29540 45305 29552 45339
rect 29586 45336 29598 45339
rect 30466 45336 30472 45348
rect 29586 45308 30472 45336
rect 29586 45305 29598 45308
rect 29540 45299 29598 45305
rect 30466 45296 30472 45308
rect 30524 45296 30530 45348
rect 31297 45339 31355 45345
rect 31297 45336 31309 45339
rect 30668 45308 31309 45336
rect 17402 45268 17408 45280
rect 17363 45240 17408 45268
rect 17402 45228 17408 45240
rect 17460 45228 17466 45280
rect 19978 45268 19984 45280
rect 19939 45240 19984 45268
rect 19978 45228 19984 45240
rect 20036 45268 20042 45280
rect 20162 45268 20168 45280
rect 20036 45240 20168 45268
rect 20036 45228 20042 45240
rect 20162 45228 20168 45240
rect 20220 45228 20226 45280
rect 20714 45268 20720 45280
rect 20675 45240 20720 45268
rect 20714 45228 20720 45240
rect 20772 45228 20778 45280
rect 23382 45268 23388 45280
rect 23343 45240 23388 45268
rect 23382 45228 23388 45240
rect 23440 45228 23446 45280
rect 24486 45268 24492 45280
rect 24447 45240 24492 45268
rect 24486 45228 24492 45240
rect 24544 45228 24550 45280
rect 30668 45277 30696 45308
rect 31297 45305 31309 45308
rect 31343 45336 31355 45339
rect 31386 45336 31392 45348
rect 31343 45308 31392 45336
rect 31343 45305 31355 45308
rect 31297 45299 31355 45305
rect 31386 45296 31392 45308
rect 31444 45296 31450 45348
rect 31478 45296 31484 45348
rect 31536 45345 31542 45348
rect 31536 45339 31560 45345
rect 31548 45305 31560 45339
rect 31536 45299 31560 45305
rect 57977 45339 58035 45345
rect 57977 45305 57989 45339
rect 58023 45336 58035 45339
rect 58802 45336 58808 45348
rect 58023 45308 58808 45336
rect 58023 45305 58035 45308
rect 57977 45299 58035 45305
rect 31536 45296 31542 45299
rect 58802 45296 58808 45308
rect 58860 45296 58866 45348
rect 30653 45271 30711 45277
rect 30653 45237 30665 45271
rect 30699 45237 30711 45271
rect 30653 45231 30711 45237
rect 1104 45178 58880 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 50326 45178
rect 50378 45126 50390 45178
rect 50442 45126 50454 45178
rect 50506 45126 50518 45178
rect 50570 45126 58880 45178
rect 1104 45104 58880 45126
rect 18138 45064 18144 45076
rect 18099 45036 18144 45064
rect 18138 45024 18144 45036
rect 18196 45024 18202 45076
rect 18601 45067 18659 45073
rect 18601 45033 18613 45067
rect 18647 45064 18659 45067
rect 18690 45064 18696 45076
rect 18647 45036 18696 45064
rect 18647 45033 18659 45036
rect 18601 45027 18659 45033
rect 18690 45024 18696 45036
rect 18748 45024 18754 45076
rect 21634 45064 21640 45076
rect 21595 45036 21640 45064
rect 21634 45024 21640 45036
rect 21692 45024 21698 45076
rect 25130 45024 25136 45076
rect 25188 45064 25194 45076
rect 27890 45064 27896 45076
rect 25188 45036 27752 45064
rect 27851 45036 27896 45064
rect 25188 45024 25194 45036
rect 17028 44999 17086 45005
rect 17028 44965 17040 44999
rect 17074 44996 17086 44999
rect 17402 44996 17408 45008
rect 17074 44968 17408 44996
rect 17074 44965 17086 44968
rect 17028 44959 17086 44965
rect 17402 44956 17408 44968
rect 17460 44956 17466 45008
rect 20070 44996 20076 45008
rect 18800 44968 20076 44996
rect 1394 44928 1400 44940
rect 1355 44900 1400 44928
rect 1394 44888 1400 44900
rect 1452 44888 1458 44940
rect 16758 44928 16764 44940
rect 16719 44900 16764 44928
rect 16758 44888 16764 44900
rect 16816 44888 16822 44940
rect 18800 44937 18828 44968
rect 20070 44956 20076 44968
rect 20128 44996 20134 45008
rect 20346 44996 20352 45008
rect 20128 44968 20352 44996
rect 20128 44956 20134 44968
rect 20346 44956 20352 44968
rect 20404 44956 20410 45008
rect 20524 44999 20582 45005
rect 20524 44965 20536 44999
rect 20570 44996 20582 44999
rect 20714 44996 20720 45008
rect 20570 44968 20720 44996
rect 20570 44965 20582 44968
rect 20524 44959 20582 44965
rect 20714 44956 20720 44968
rect 20772 44956 20778 45008
rect 25584 44999 25642 45005
rect 25584 44965 25596 44999
rect 25630 44996 25642 44999
rect 26418 44996 26424 45008
rect 25630 44968 26424 44996
rect 25630 44965 25642 44968
rect 25584 44959 25642 44965
rect 26418 44956 26424 44968
rect 26476 44956 26482 45008
rect 27724 44996 27752 45036
rect 27890 45024 27896 45036
rect 27948 45024 27954 45076
rect 30466 45064 30472 45076
rect 30427 45036 30472 45064
rect 30466 45024 30472 45036
rect 30524 45024 30530 45076
rect 30653 45067 30711 45073
rect 30653 45033 30665 45067
rect 30699 45064 30711 45067
rect 31478 45064 31484 45076
rect 30699 45036 31484 45064
rect 30699 45033 30711 45036
rect 30653 45027 30711 45033
rect 31478 45024 31484 45036
rect 31536 45024 31542 45076
rect 27724 44968 28672 44996
rect 18785 44931 18843 44937
rect 18785 44897 18797 44931
rect 18831 44897 18843 44931
rect 18785 44891 18843 44897
rect 19061 44931 19119 44937
rect 19061 44897 19073 44931
rect 19107 44928 19119 44931
rect 19978 44928 19984 44940
rect 19107 44900 19984 44928
rect 19107 44897 19119 44900
rect 19061 44891 19119 44897
rect 19978 44888 19984 44900
rect 20036 44888 20042 44940
rect 22741 44931 22799 44937
rect 22741 44897 22753 44931
rect 22787 44928 22799 44931
rect 23382 44928 23388 44940
rect 22787 44900 23388 44928
rect 22787 44897 22799 44900
rect 22741 44891 22799 44897
rect 23382 44888 23388 44900
rect 23440 44888 23446 44940
rect 24029 44931 24087 44937
rect 24029 44897 24041 44931
rect 24075 44928 24087 44931
rect 24486 44928 24492 44940
rect 24075 44900 24492 44928
rect 24075 44897 24087 44900
rect 24029 44891 24087 44897
rect 24486 44888 24492 44900
rect 24544 44888 24550 44940
rect 24670 44888 24676 44940
rect 24728 44928 24734 44940
rect 25317 44931 25375 44937
rect 25317 44928 25329 44931
rect 24728 44900 25329 44928
rect 24728 44888 24734 44900
rect 25317 44897 25329 44900
rect 25363 44897 25375 44931
rect 27157 44931 27215 44937
rect 27157 44928 27169 44931
rect 25317 44891 25375 44897
rect 26712 44900 27169 44928
rect 19426 44820 19432 44872
rect 19484 44860 19490 44872
rect 20257 44863 20315 44869
rect 20257 44860 20269 44863
rect 19484 44832 20269 44860
rect 19484 44820 19490 44832
rect 20257 44829 20269 44832
rect 20303 44829 20315 44863
rect 22922 44860 22928 44872
rect 22883 44832 22928 44860
rect 20257 44823 20315 44829
rect 22922 44820 22928 44832
rect 22980 44820 22986 44872
rect 23017 44863 23075 44869
rect 23017 44829 23029 44863
rect 23063 44860 23075 44863
rect 23934 44860 23940 44872
rect 23063 44832 23940 44860
rect 23063 44829 23075 44832
rect 23017 44823 23075 44829
rect 23934 44820 23940 44832
rect 23992 44820 23998 44872
rect 24302 44860 24308 44872
rect 24263 44832 24308 44860
rect 24302 44820 24308 44832
rect 24360 44820 24366 44872
rect 18969 44795 19027 44801
rect 18969 44761 18981 44795
rect 19015 44792 19027 44795
rect 19334 44792 19340 44804
rect 19015 44764 19340 44792
rect 19015 44761 19027 44764
rect 18969 44755 19027 44761
rect 19334 44752 19340 44764
rect 19392 44792 19398 44804
rect 19886 44792 19892 44804
rect 19392 44764 19892 44792
rect 19392 44752 19398 44764
rect 19886 44752 19892 44764
rect 19944 44752 19950 44804
rect 26712 44801 26740 44900
rect 27157 44897 27169 44900
rect 27203 44897 27215 44931
rect 27157 44891 27215 44897
rect 27614 44888 27620 44940
rect 27672 44928 27678 44940
rect 28644 44937 28672 44968
rect 31938 44956 31944 45008
rect 31996 44996 32002 45008
rect 32033 44999 32091 45005
rect 32033 44996 32045 44999
rect 31996 44968 32045 44996
rect 31996 44956 32002 44968
rect 32033 44965 32045 44968
rect 32079 44996 32091 44999
rect 33962 44996 33968 45008
rect 32079 44968 33968 44996
rect 32079 44965 32091 44968
rect 32033 44959 32091 44965
rect 33962 44956 33968 44968
rect 34020 44956 34026 45008
rect 27801 44931 27859 44937
rect 27801 44928 27813 44931
rect 27672 44900 27813 44928
rect 27672 44888 27678 44900
rect 27801 44897 27813 44900
rect 27847 44897 27859 44931
rect 27801 44891 27859 44897
rect 28629 44931 28687 44937
rect 28629 44897 28641 44931
rect 28675 44897 28687 44931
rect 28629 44891 28687 44897
rect 28902 44888 28908 44940
rect 28960 44928 28966 44940
rect 29089 44931 29147 44937
rect 29089 44928 29101 44931
rect 28960 44900 29101 44928
rect 28960 44888 28966 44900
rect 29089 44897 29101 44900
rect 29135 44897 29147 44931
rect 29089 44891 29147 44897
rect 29273 44931 29331 44937
rect 29273 44897 29285 44931
rect 29319 44897 29331 44931
rect 29273 44891 29331 44897
rect 30650 44931 30708 44937
rect 30650 44897 30662 44931
rect 30696 44928 30708 44931
rect 31113 44931 31171 44937
rect 31113 44928 31125 44931
rect 30696 44900 31125 44928
rect 30696 44897 30708 44900
rect 30650 44891 30708 44897
rect 31113 44897 31125 44900
rect 31159 44928 31171 44931
rect 31386 44928 31392 44940
rect 31159 44900 31392 44928
rect 31159 44897 31171 44900
rect 31113 44891 31171 44897
rect 28994 44820 29000 44872
rect 29052 44860 29058 44872
rect 29288 44860 29316 44891
rect 31386 44888 31392 44900
rect 31444 44888 31450 44940
rect 32214 44928 32220 44940
rect 32175 44900 32220 44928
rect 32214 44888 32220 44900
rect 32272 44888 32278 44940
rect 32306 44888 32312 44940
rect 32364 44928 32370 44940
rect 32364 44900 32409 44928
rect 32364 44888 32370 44900
rect 56962 44888 56968 44940
rect 57020 44928 57026 44940
rect 57241 44931 57299 44937
rect 57241 44928 57253 44931
rect 57020 44900 57253 44928
rect 57020 44888 57026 44900
rect 57241 44897 57253 44900
rect 57287 44928 57299 44931
rect 57606 44928 57612 44940
rect 57287 44900 57612 44928
rect 57287 44897 57299 44900
rect 57241 44891 57299 44897
rect 57606 44888 57612 44900
rect 57664 44888 57670 44940
rect 57974 44928 57980 44940
rect 57935 44900 57980 44928
rect 57974 44888 57980 44900
rect 58032 44888 58038 44940
rect 58158 44928 58164 44940
rect 58119 44900 58164 44928
rect 58158 44888 58164 44900
rect 58216 44888 58222 44940
rect 29052 44832 29316 44860
rect 29052 44820 29058 44832
rect 26697 44795 26755 44801
rect 26697 44761 26709 44795
rect 26743 44761 26755 44795
rect 26697 44755 26755 44761
rect 28445 44795 28503 44801
rect 28445 44761 28457 44795
rect 28491 44792 28503 44795
rect 30650 44792 30656 44804
rect 28491 44764 30656 44792
rect 28491 44761 28503 44764
rect 28445 44755 28503 44761
rect 30650 44752 30656 44764
rect 30708 44752 30714 44804
rect 31021 44795 31079 44801
rect 31021 44761 31033 44795
rect 31067 44792 31079 44795
rect 31478 44792 31484 44804
rect 31067 44764 31484 44792
rect 31067 44761 31079 44764
rect 31021 44755 31079 44761
rect 31478 44752 31484 44764
rect 31536 44792 31542 44804
rect 32122 44792 32128 44804
rect 31536 44764 32128 44792
rect 31536 44752 31542 44764
rect 32122 44752 32128 44764
rect 32180 44752 32186 44804
rect 22557 44727 22615 44733
rect 22557 44693 22569 44727
rect 22603 44724 22615 44727
rect 22646 44724 22652 44736
rect 22603 44696 22652 44724
rect 22603 44693 22615 44696
rect 22557 44687 22615 44693
rect 22646 44684 22652 44696
rect 22704 44684 22710 44736
rect 23842 44724 23848 44736
rect 23803 44696 23848 44724
rect 23842 44684 23848 44696
rect 23900 44684 23906 44736
rect 24210 44724 24216 44736
rect 24171 44696 24216 44724
rect 24210 44684 24216 44696
rect 24268 44684 24274 44736
rect 27246 44724 27252 44736
rect 27207 44696 27252 44724
rect 27246 44684 27252 44696
rect 27304 44684 27310 44736
rect 29086 44724 29092 44736
rect 29047 44696 29092 44724
rect 29086 44684 29092 44696
rect 29144 44684 29150 44736
rect 32030 44724 32036 44736
rect 31991 44696 32036 44724
rect 32030 44684 32036 44696
rect 32088 44684 32094 44736
rect 57330 44684 57336 44736
rect 57388 44724 57394 44736
rect 57425 44727 57483 44733
rect 57425 44724 57437 44727
rect 57388 44696 57437 44724
rect 57388 44684 57394 44696
rect 57425 44693 57437 44696
rect 57471 44693 57483 44727
rect 57425 44687 57483 44693
rect 1104 44634 58880 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 58880 44634
rect 1104 44560 58880 44582
rect 17586 44480 17592 44532
rect 17644 44520 17650 44532
rect 17773 44523 17831 44529
rect 17773 44520 17785 44523
rect 17644 44492 17785 44520
rect 17644 44480 17650 44492
rect 17773 44489 17785 44492
rect 17819 44489 17831 44523
rect 17773 44483 17831 44489
rect 18601 44523 18659 44529
rect 18601 44489 18613 44523
rect 18647 44520 18659 44523
rect 19334 44520 19340 44532
rect 18647 44492 19340 44520
rect 18647 44489 18659 44492
rect 18601 44483 18659 44489
rect 17788 44384 17816 44483
rect 19334 44480 19340 44492
rect 19392 44480 19398 44532
rect 20898 44480 20904 44532
rect 20956 44520 20962 44532
rect 21085 44523 21143 44529
rect 21085 44520 21097 44523
rect 20956 44492 21097 44520
rect 20956 44480 20962 44492
rect 21085 44489 21097 44492
rect 21131 44489 21143 44523
rect 23934 44520 23940 44532
rect 23895 44492 23940 44520
rect 21085 44483 21143 44489
rect 23934 44480 23940 44492
rect 23992 44480 23998 44532
rect 24302 44480 24308 44532
rect 24360 44520 24366 44532
rect 25777 44523 25835 44529
rect 25777 44520 25789 44523
rect 24360 44492 25789 44520
rect 24360 44480 24366 44492
rect 25777 44489 25789 44492
rect 25823 44489 25835 44523
rect 28442 44520 28448 44532
rect 28403 44492 28448 44520
rect 25777 44483 25835 44489
rect 28442 44480 28448 44492
rect 28500 44480 28506 44532
rect 31938 44520 31944 44532
rect 31899 44492 31944 44520
rect 31938 44480 31944 44492
rect 31996 44480 32002 44532
rect 32122 44520 32128 44532
rect 32083 44492 32128 44520
rect 32122 44480 32128 44492
rect 32180 44480 32186 44532
rect 57974 44520 57980 44532
rect 57935 44492 57980 44520
rect 57974 44480 57980 44492
rect 58032 44480 58038 44532
rect 26881 44455 26939 44461
rect 26881 44421 26893 44455
rect 26927 44452 26939 44455
rect 28123 44455 28181 44461
rect 28123 44452 28135 44455
rect 26927 44424 28135 44452
rect 26927 44421 26939 44424
rect 26881 44415 26939 44421
rect 28123 44421 28135 44424
rect 28169 44421 28181 44455
rect 28123 44415 28181 44421
rect 28258 44412 28264 44464
rect 28316 44452 28322 44464
rect 28316 44424 28361 44452
rect 28316 44412 28322 44424
rect 17788 44356 18552 44384
rect 17681 44319 17739 44325
rect 17681 44285 17693 44319
rect 17727 44285 17739 44319
rect 17681 44279 17739 44285
rect 17865 44319 17923 44325
rect 17865 44285 17877 44319
rect 17911 44316 17923 44319
rect 18138 44316 18144 44328
rect 17911 44288 18144 44316
rect 17911 44285 17923 44288
rect 17865 44279 17923 44285
rect 17696 44248 17724 44279
rect 18138 44276 18144 44288
rect 18196 44276 18202 44328
rect 18524 44325 18552 44356
rect 23842 44344 23848 44396
rect 23900 44384 23906 44396
rect 28353 44387 28411 44393
rect 23900 44356 24532 44384
rect 23900 44344 23906 44356
rect 18509 44319 18567 44325
rect 18509 44285 18521 44319
rect 18555 44285 18567 44319
rect 20346 44316 20352 44328
rect 20307 44288 20352 44316
rect 18509 44279 18567 44285
rect 20346 44276 20352 44288
rect 20404 44276 20410 44328
rect 20441 44319 20499 44325
rect 20441 44285 20453 44319
rect 20487 44316 20499 44319
rect 20990 44316 20996 44328
rect 20487 44288 20996 44316
rect 20487 44285 20499 44288
rect 20441 44279 20499 44285
rect 20990 44276 20996 44288
rect 21048 44276 21054 44328
rect 21177 44319 21235 44325
rect 21177 44285 21189 44319
rect 21223 44316 21235 44319
rect 21634 44316 21640 44328
rect 21223 44288 21640 44316
rect 21223 44285 21235 44288
rect 21177 44279 21235 44285
rect 21634 44276 21640 44288
rect 21692 44276 21698 44328
rect 22554 44316 22560 44328
rect 22515 44288 22560 44316
rect 22554 44276 22560 44288
rect 22612 44276 22618 44328
rect 22646 44276 22652 44328
rect 22704 44316 22710 44328
rect 22813 44319 22871 44325
rect 22813 44316 22825 44319
rect 22704 44288 22825 44316
rect 22704 44276 22710 44288
rect 22813 44285 22825 44288
rect 22859 44285 22871 44319
rect 22813 44279 22871 44285
rect 24397 44319 24455 44325
rect 24397 44285 24409 44319
rect 24443 44285 24455 44319
rect 24504 44316 24532 44356
rect 28353 44353 28365 44387
rect 28399 44384 28411 44387
rect 28994 44384 29000 44396
rect 28399 44356 29000 44384
rect 28399 44353 28411 44356
rect 28353 44347 28411 44353
rect 28994 44344 29000 44356
rect 29052 44344 29058 44396
rect 32140 44384 32168 44480
rect 33042 44452 33048 44464
rect 33003 44424 33048 44452
rect 33042 44412 33048 44424
rect 33100 44412 33106 44464
rect 56873 44455 56931 44461
rect 56873 44421 56885 44455
rect 56919 44452 56931 44455
rect 56919 44424 57744 44452
rect 56919 44421 56931 44424
rect 56873 44415 56931 44421
rect 57716 44393 57744 44424
rect 56413 44387 56471 44393
rect 32140 44356 33272 44384
rect 24653 44319 24711 44325
rect 24653 44316 24665 44319
rect 24504 44288 24665 44316
rect 24397 44279 24455 44285
rect 24653 44285 24665 44288
rect 24699 44285 24711 44319
rect 24653 44279 24711 44285
rect 17954 44248 17960 44260
rect 17696 44220 17960 44248
rect 17954 44208 17960 44220
rect 18012 44208 18018 44260
rect 24412 44248 24440 44279
rect 26326 44276 26332 44328
rect 26384 44316 26390 44328
rect 26513 44319 26571 44325
rect 26513 44316 26525 44319
rect 26384 44288 26525 44316
rect 26384 44276 26390 44288
rect 26513 44285 26525 44288
rect 26559 44316 26571 44319
rect 27246 44316 27252 44328
rect 26559 44288 27252 44316
rect 26559 44285 26571 44288
rect 26513 44279 26571 44285
rect 27246 44276 27252 44288
rect 27304 44276 27310 44328
rect 29273 44319 29331 44325
rect 29273 44285 29285 44319
rect 29319 44316 29331 44319
rect 30558 44316 30564 44328
rect 29319 44288 30564 44316
rect 29319 44285 29331 44288
rect 29273 44279 29331 44285
rect 30558 44276 30564 44288
rect 30616 44276 30622 44328
rect 32030 44276 32036 44328
rect 32088 44316 32094 44328
rect 33244 44325 33272 44356
rect 56413 44353 56425 44387
rect 56459 44384 56471 44387
rect 57517 44387 57575 44393
rect 57517 44384 57529 44387
rect 56459 44356 57529 44384
rect 56459 44353 56471 44356
rect 56413 44347 56471 44353
rect 57517 44353 57529 44356
rect 57563 44353 57575 44387
rect 57517 44347 57575 44353
rect 57701 44387 57759 44393
rect 57701 44353 57713 44387
rect 57747 44353 57759 44387
rect 57701 44347 57759 44353
rect 33045 44319 33103 44325
rect 33045 44316 33057 44319
rect 32088 44288 33057 44316
rect 32088 44276 32094 44288
rect 33045 44285 33057 44288
rect 33091 44285 33103 44319
rect 33045 44279 33103 44285
rect 33229 44319 33287 44325
rect 33229 44285 33241 44319
rect 33275 44285 33287 44319
rect 33229 44279 33287 44285
rect 57057 44319 57115 44325
rect 57057 44285 57069 44319
rect 57103 44316 57115 44319
rect 57330 44316 57336 44328
rect 57103 44288 57336 44316
rect 57103 44285 57115 44288
rect 57057 44279 57115 44285
rect 57330 44276 57336 44288
rect 57388 44276 57394 44328
rect 25222 44248 25228 44260
rect 24412 44220 25228 44248
rect 25222 44208 25228 44220
rect 25280 44208 25286 44260
rect 26694 44248 26700 44260
rect 26655 44220 26700 44248
rect 26694 44208 26700 44220
rect 26752 44208 26758 44260
rect 27985 44251 28043 44257
rect 27985 44217 27997 44251
rect 28031 44248 28043 44251
rect 28074 44248 28080 44260
rect 28031 44220 28080 44248
rect 28031 44217 28043 44220
rect 27985 44211 28043 44217
rect 28074 44208 28080 44220
rect 28132 44208 28138 44260
rect 29362 44208 29368 44260
rect 29420 44248 29426 44260
rect 29518 44251 29576 44257
rect 29518 44248 29530 44251
rect 29420 44220 29530 44248
rect 29420 44208 29426 44220
rect 29518 44217 29530 44220
rect 29564 44217 29576 44251
rect 29518 44211 29576 44217
rect 31757 44251 31815 44257
rect 31757 44217 31769 44251
rect 31803 44248 31815 44251
rect 32214 44248 32220 44260
rect 31803 44220 32220 44248
rect 31803 44217 31815 44220
rect 31757 44211 31815 44217
rect 32214 44208 32220 44220
rect 32272 44208 32278 44260
rect 30466 44140 30472 44192
rect 30524 44180 30530 44192
rect 30653 44183 30711 44189
rect 30653 44180 30665 44183
rect 30524 44152 30665 44180
rect 30524 44140 30530 44152
rect 30653 44149 30665 44152
rect 30699 44149 30711 44183
rect 30653 44143 30711 44149
rect 31938 44140 31944 44192
rect 31996 44189 32002 44192
rect 31996 44183 32020 44189
rect 32008 44180 32020 44183
rect 32306 44180 32312 44192
rect 32008 44152 32312 44180
rect 32008 44149 32020 44152
rect 31996 44143 32020 44149
rect 31996 44140 32002 44143
rect 32306 44140 32312 44152
rect 32364 44140 32370 44192
rect 1104 44090 58880 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 58880 44090
rect 1104 44016 58880 44038
rect 23753 43979 23811 43985
rect 23753 43945 23765 43979
rect 23799 43976 23811 43979
rect 24210 43976 24216 43988
rect 23799 43948 24216 43976
rect 23799 43945 23811 43948
rect 23753 43939 23811 43945
rect 24210 43936 24216 43948
rect 24268 43936 24274 43988
rect 25130 43936 25136 43988
rect 25188 43976 25194 43988
rect 25225 43979 25283 43985
rect 25225 43976 25237 43979
rect 25188 43948 25237 43976
rect 25188 43936 25194 43948
rect 25225 43945 25237 43948
rect 25271 43945 25283 43979
rect 25225 43939 25283 43945
rect 26145 43979 26203 43985
rect 26145 43945 26157 43979
rect 26191 43976 26203 43979
rect 26234 43976 26240 43988
rect 26191 43948 26240 43976
rect 26191 43945 26203 43948
rect 26145 43939 26203 43945
rect 26234 43936 26240 43948
rect 26292 43936 26298 43988
rect 29457 43979 29515 43985
rect 29457 43945 29469 43979
rect 29503 43976 29515 43979
rect 30561 43979 30619 43985
rect 30561 43976 30573 43979
rect 29503 43948 30573 43976
rect 29503 43945 29515 43948
rect 29457 43939 29515 43945
rect 30561 43945 30573 43948
rect 30607 43945 30619 43979
rect 30561 43939 30619 43945
rect 31573 43979 31631 43985
rect 31573 43945 31585 43979
rect 31619 43976 31631 43979
rect 31938 43976 31944 43988
rect 31619 43948 31944 43976
rect 31619 43945 31631 43948
rect 31573 43939 31631 43945
rect 21082 43908 21088 43920
rect 21043 43880 21088 43908
rect 21082 43868 21088 43880
rect 21140 43868 21146 43920
rect 21174 43868 21180 43920
rect 21232 43908 21238 43920
rect 21290 43911 21348 43917
rect 21290 43908 21302 43911
rect 21232 43880 21302 43908
rect 21232 43868 21238 43880
rect 21290 43877 21302 43880
rect 21336 43877 21348 43911
rect 21290 43871 21348 43877
rect 27525 43911 27583 43917
rect 27525 43877 27537 43911
rect 27571 43908 27583 43911
rect 28994 43908 29000 43920
rect 27571 43880 28212 43908
rect 27571 43877 27583 43880
rect 27525 43871 27583 43877
rect 1394 43840 1400 43852
rect 1355 43812 1400 43840
rect 1394 43800 1400 43812
rect 1452 43800 1458 43852
rect 20441 43843 20499 43849
rect 20441 43809 20453 43843
rect 20487 43809 20499 43843
rect 20441 43803 20499 43809
rect 20625 43843 20683 43849
rect 20625 43809 20637 43843
rect 20671 43840 20683 43843
rect 20671 43812 21496 43840
rect 20671 43809 20683 43812
rect 20625 43803 20683 43809
rect 20456 43772 20484 43803
rect 20898 43772 20904 43784
rect 20456 43744 20904 43772
rect 20898 43732 20904 43744
rect 20956 43732 20962 43784
rect 21468 43713 21496 43812
rect 23382 43800 23388 43852
rect 23440 43840 23446 43852
rect 23661 43843 23719 43849
rect 23661 43840 23673 43843
rect 23440 43812 23673 43840
rect 23440 43800 23446 43812
rect 23661 43809 23673 43812
rect 23707 43809 23719 43843
rect 23661 43803 23719 43809
rect 25314 43800 25320 43852
rect 25372 43840 25378 43852
rect 25409 43843 25467 43849
rect 25409 43840 25421 43843
rect 25372 43812 25421 43840
rect 25372 43800 25378 43812
rect 25409 43809 25421 43812
rect 25455 43809 25467 43843
rect 26326 43840 26332 43852
rect 26287 43812 26332 43840
rect 25409 43803 25467 43809
rect 26326 43800 26332 43812
rect 26384 43800 26390 43852
rect 27433 43843 27491 43849
rect 27433 43809 27445 43843
rect 27479 43840 27491 43843
rect 27890 43840 27896 43852
rect 27479 43812 27896 43840
rect 27479 43809 27491 43812
rect 27433 43803 27491 43809
rect 27890 43800 27896 43812
rect 27948 43800 27954 43852
rect 28074 43840 28080 43852
rect 28035 43812 28080 43840
rect 28074 43800 28080 43812
rect 28132 43800 28138 43852
rect 28184 43849 28212 43880
rect 28368 43880 29000 43908
rect 28169 43843 28227 43849
rect 28169 43809 28181 43843
rect 28215 43840 28227 43843
rect 28258 43840 28264 43852
rect 28215 43812 28264 43840
rect 28215 43809 28227 43812
rect 28169 43803 28227 43809
rect 28258 43800 28264 43812
rect 28316 43800 28322 43852
rect 28368 43849 28396 43880
rect 28994 43868 29000 43880
rect 29052 43908 29058 43920
rect 29472 43908 29500 43939
rect 31938 43936 31944 43948
rect 31996 43936 32002 43988
rect 33962 43976 33968 43988
rect 33923 43948 33968 43976
rect 33962 43936 33968 43948
rect 34020 43936 34026 43988
rect 32214 43908 32220 43920
rect 29052 43880 29500 43908
rect 31726 43880 32220 43908
rect 29052 43868 29058 43880
rect 28353 43843 28411 43849
rect 28353 43809 28365 43843
rect 28399 43809 28411 43843
rect 28353 43803 28411 43809
rect 29086 43800 29092 43852
rect 29144 43840 29150 43852
rect 29273 43843 29331 43849
rect 29273 43840 29285 43843
rect 29144 43812 29285 43840
rect 29144 43800 29150 43812
rect 29273 43809 29285 43812
rect 29319 43809 29331 43843
rect 29273 43803 29331 43809
rect 29549 43843 29607 43849
rect 29549 43809 29561 43843
rect 29595 43809 29607 43843
rect 30466 43840 30472 43852
rect 30427 43812 30472 43840
rect 29549 43803 29607 43809
rect 26605 43775 26663 43781
rect 26605 43741 26617 43775
rect 26651 43772 26663 43775
rect 26694 43772 26700 43784
rect 26651 43744 26700 43772
rect 26651 43741 26663 43744
rect 26605 43735 26663 43741
rect 26694 43732 26700 43744
rect 26752 43732 26758 43784
rect 27522 43732 27528 43784
rect 27580 43772 27586 43784
rect 28537 43775 28595 43781
rect 28537 43772 28549 43775
rect 27580 43744 28549 43772
rect 27580 43732 27586 43744
rect 28537 43741 28549 43744
rect 28583 43741 28595 43775
rect 29564 43772 29592 43803
rect 30466 43800 30472 43812
rect 30524 43800 30530 43852
rect 31570 43843 31628 43849
rect 31570 43809 31582 43843
rect 31616 43840 31628 43843
rect 31726 43840 31754 43880
rect 32214 43868 32220 43880
rect 32272 43868 32278 43920
rect 32852 43911 32910 43917
rect 32852 43877 32864 43911
rect 32898 43908 32910 43911
rect 33042 43908 33048 43920
rect 32898 43880 33048 43908
rect 32898 43877 32910 43880
rect 32852 43871 32910 43877
rect 33042 43868 33048 43880
rect 33100 43868 33106 43920
rect 58158 43908 58164 43920
rect 58119 43880 58164 43908
rect 58158 43868 58164 43880
rect 58216 43868 58222 43920
rect 32585 43843 32643 43849
rect 32585 43840 32597 43843
rect 31616 43812 31754 43840
rect 31956 43812 32597 43840
rect 31616 43809 31628 43812
rect 31570 43803 31628 43809
rect 28537 43735 28595 43741
rect 29196 43744 29592 43772
rect 21453 43707 21511 43713
rect 21453 43673 21465 43707
rect 21499 43704 21511 43707
rect 22738 43704 22744 43716
rect 21499 43676 22744 43704
rect 21499 43673 21511 43676
rect 21453 43667 21511 43673
rect 22738 43664 22744 43676
rect 22796 43664 22802 43716
rect 26326 43664 26332 43716
rect 26384 43704 26390 43716
rect 26513 43707 26571 43713
rect 26513 43704 26525 43707
rect 26384 43676 26525 43704
rect 26384 43664 26390 43676
rect 26513 43673 26525 43676
rect 26559 43704 26571 43707
rect 27540 43704 27568 43732
rect 26559 43676 27568 43704
rect 26559 43673 26571 43676
rect 26513 43667 26571 43673
rect 28074 43664 28080 43716
rect 28132 43704 28138 43716
rect 28902 43704 28908 43716
rect 28132 43676 28908 43704
rect 28132 43664 28138 43676
rect 28902 43664 28908 43676
rect 28960 43704 28966 43716
rect 29196 43704 29224 43744
rect 30558 43732 30564 43784
rect 30616 43772 30622 43784
rect 31662 43772 31668 43784
rect 30616 43744 31668 43772
rect 30616 43732 30622 43744
rect 31662 43732 31668 43744
rect 31720 43772 31726 43784
rect 31956 43772 31984 43812
rect 32585 43809 32597 43812
rect 32631 43809 32643 43843
rect 32585 43803 32643 43809
rect 54938 43800 54944 43852
rect 54996 43840 55002 43852
rect 57977 43843 58035 43849
rect 57977 43840 57989 43843
rect 54996 43812 57989 43840
rect 54996 43800 55002 43812
rect 57977 43809 57989 43812
rect 58023 43809 58035 43843
rect 57977 43803 58035 43809
rect 31720 43744 31984 43772
rect 32033 43775 32091 43781
rect 31720 43732 31726 43744
rect 32033 43741 32045 43775
rect 32079 43772 32091 43775
rect 32214 43772 32220 43784
rect 32079 43744 32220 43772
rect 32079 43741 32091 43744
rect 32033 43735 32091 43741
rect 32214 43732 32220 43744
rect 32272 43732 32278 43784
rect 28960 43676 29224 43704
rect 29273 43707 29331 43713
rect 28960 43664 28966 43676
rect 29273 43673 29285 43707
rect 29319 43704 29331 43707
rect 29362 43704 29368 43716
rect 29319 43676 29368 43704
rect 29319 43673 29331 43676
rect 29273 43667 29331 43673
rect 29362 43664 29368 43676
rect 29420 43664 29426 43716
rect 20438 43636 20444 43648
rect 20399 43608 20444 43636
rect 20438 43596 20444 43608
rect 20496 43596 20502 43648
rect 21269 43639 21327 43645
rect 21269 43605 21281 43639
rect 21315 43636 21327 43639
rect 21358 43636 21364 43648
rect 21315 43608 21364 43636
rect 21315 43605 21327 43608
rect 21269 43599 21327 43605
rect 21358 43596 21364 43608
rect 21416 43596 21422 43648
rect 31386 43636 31392 43648
rect 31347 43608 31392 43636
rect 31386 43596 31392 43608
rect 31444 43596 31450 43648
rect 31938 43636 31944 43648
rect 31851 43608 31944 43636
rect 31938 43596 31944 43608
rect 31996 43636 32002 43648
rect 32858 43636 32864 43648
rect 31996 43608 32864 43636
rect 31996 43596 32002 43608
rect 32858 43596 32864 43608
rect 32916 43596 32922 43648
rect 57422 43636 57428 43648
rect 57383 43608 57428 43636
rect 57422 43596 57428 43608
rect 57480 43596 57486 43648
rect 1104 43546 58880 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 58880 43546
rect 1104 43472 58880 43494
rect 26326 43432 26332 43444
rect 26287 43404 26332 43432
rect 26326 43392 26332 43404
rect 26384 43392 26390 43444
rect 32033 43435 32091 43441
rect 32033 43401 32045 43435
rect 32079 43432 32091 43435
rect 32214 43432 32220 43444
rect 32079 43404 32220 43432
rect 32079 43401 32091 43404
rect 32033 43395 32091 43401
rect 32214 43392 32220 43404
rect 32272 43392 32278 43444
rect 22738 43324 22744 43376
rect 22796 43364 22802 43376
rect 23109 43367 23167 43373
rect 23109 43364 23121 43367
rect 22796 43336 23121 43364
rect 22796 43324 22802 43336
rect 23109 43333 23121 43336
rect 23155 43364 23167 43367
rect 23658 43364 23664 43376
rect 23155 43336 23664 43364
rect 23155 43333 23167 43336
rect 23109 43327 23167 43333
rect 23658 43324 23664 43336
rect 23716 43324 23722 43376
rect 30558 43324 30564 43376
rect 30616 43364 30622 43376
rect 58158 43364 58164 43376
rect 30616 43336 30696 43364
rect 58119 43336 58164 43364
rect 30616 43324 30622 43336
rect 30668 43305 30696 43336
rect 58158 43324 58164 43336
rect 58216 43324 58222 43376
rect 30653 43299 30711 43305
rect 23032 43268 23244 43296
rect 20162 43228 20168 43240
rect 20123 43200 20168 43228
rect 20162 43188 20168 43200
rect 20220 43188 20226 43240
rect 20438 43237 20444 43240
rect 20432 43228 20444 43237
rect 20399 43200 20444 43228
rect 20432 43191 20444 43200
rect 20438 43188 20444 43191
rect 20496 43188 20502 43240
rect 22738 43231 22796 43237
rect 22738 43197 22750 43231
rect 22784 43228 22796 43231
rect 23032 43228 23060 43268
rect 23216 43237 23244 43268
rect 30653 43265 30665 43299
rect 30699 43265 30711 43299
rect 30653 43259 30711 43265
rect 22784 43200 23060 43228
rect 23201 43231 23259 43237
rect 22784 43197 22796 43200
rect 22738 43191 22796 43197
rect 23201 43197 23213 43231
rect 23247 43228 23259 43231
rect 23382 43228 23388 43240
rect 23247 43200 23388 43228
rect 23247 43197 23259 43200
rect 23201 43191 23259 43197
rect 23382 43188 23388 43200
rect 23440 43188 23446 43240
rect 23753 43231 23811 43237
rect 23753 43197 23765 43231
rect 23799 43197 23811 43231
rect 23753 43191 23811 43197
rect 26053 43231 26111 43237
rect 26053 43197 26065 43231
rect 26099 43197 26111 43231
rect 26053 43191 26111 43197
rect 26145 43231 26203 43237
rect 26145 43197 26157 43231
rect 26191 43228 26203 43231
rect 26234 43228 26240 43240
rect 26191 43200 26240 43228
rect 26191 43197 26203 43200
rect 26145 43191 26203 43197
rect 22646 43120 22652 43172
rect 22704 43160 22710 43172
rect 23768 43160 23796 43191
rect 22704 43132 23796 43160
rect 24020 43163 24078 43169
rect 22704 43120 22710 43132
rect 24020 43129 24032 43163
rect 24066 43160 24078 43163
rect 24302 43160 24308 43172
rect 24066 43132 24308 43160
rect 24066 43129 24078 43132
rect 24020 43123 24078 43129
rect 24302 43120 24308 43132
rect 24360 43120 24366 43172
rect 26068 43160 26096 43191
rect 26234 43188 26240 43200
rect 26292 43188 26298 43240
rect 26421 43231 26479 43237
rect 26421 43197 26433 43231
rect 26467 43228 26479 43231
rect 26694 43228 26700 43240
rect 26467 43200 26700 43228
rect 26467 43197 26479 43200
rect 26421 43191 26479 43197
rect 26694 43188 26700 43200
rect 26752 43228 26758 43240
rect 27154 43228 27160 43240
rect 26752 43200 27160 43228
rect 26752 43188 26758 43200
rect 27154 43188 27160 43200
rect 27212 43188 27218 43240
rect 27798 43228 27804 43240
rect 27759 43200 27804 43228
rect 27798 43188 27804 43200
rect 27856 43188 27862 43240
rect 28902 43188 28908 43240
rect 28960 43228 28966 43240
rect 29641 43231 29699 43237
rect 29641 43228 29653 43231
rect 28960 43200 29653 43228
rect 28960 43188 28966 43200
rect 29641 43197 29653 43200
rect 29687 43197 29699 43231
rect 29641 43191 29699 43197
rect 29825 43231 29883 43237
rect 29825 43197 29837 43231
rect 29871 43228 29883 43231
rect 30558 43228 30564 43240
rect 29871 43200 30564 43228
rect 29871 43197 29883 43200
rect 29825 43191 29883 43197
rect 30558 43188 30564 43200
rect 30616 43188 30622 43240
rect 30920 43231 30978 43237
rect 30920 43197 30932 43231
rect 30966 43228 30978 43231
rect 31386 43228 31392 43240
rect 30966 43200 31392 43228
rect 30966 43197 30978 43200
rect 30920 43191 30978 43197
rect 31386 43188 31392 43200
rect 31444 43188 31450 43240
rect 56502 43188 56508 43240
rect 56560 43228 56566 43240
rect 56597 43231 56655 43237
rect 56597 43228 56609 43231
rect 56560 43200 56609 43228
rect 56560 43188 56566 43200
rect 56597 43197 56609 43200
rect 56643 43197 56655 43231
rect 56597 43191 56655 43197
rect 57330 43188 57336 43240
rect 57388 43228 57394 43240
rect 57425 43231 57483 43237
rect 57425 43228 57437 43231
rect 57388 43200 57437 43228
rect 57388 43188 57394 43200
rect 57425 43197 57437 43200
rect 57471 43197 57483 43231
rect 57425 43191 57483 43197
rect 26602 43160 26608 43172
rect 26068 43132 26608 43160
rect 26602 43120 26608 43132
rect 26660 43120 26666 43172
rect 27982 43120 27988 43172
rect 28040 43169 28046 43172
rect 28040 43163 28104 43169
rect 28040 43129 28058 43163
rect 28092 43129 28104 43163
rect 28040 43123 28104 43129
rect 28040 43120 28046 43123
rect 29730 43120 29736 43172
rect 29788 43160 29794 43172
rect 30009 43163 30067 43169
rect 30009 43160 30021 43163
rect 29788 43132 30021 43160
rect 29788 43120 29794 43132
rect 30009 43129 30021 43132
rect 30055 43129 30067 43163
rect 57974 43160 57980 43172
rect 57935 43132 57980 43160
rect 30009 43123 30067 43129
rect 57974 43120 57980 43132
rect 58032 43120 58038 43172
rect 21358 43052 21364 43104
rect 21416 43092 21422 43104
rect 21545 43095 21603 43101
rect 21545 43092 21557 43095
rect 21416 43064 21557 43092
rect 21416 43052 21422 43064
rect 21545 43061 21557 43064
rect 21591 43061 21603 43095
rect 22554 43092 22560 43104
rect 22515 43064 22560 43092
rect 21545 43055 21603 43061
rect 22554 43052 22560 43064
rect 22612 43052 22618 43104
rect 22738 43092 22744 43104
rect 22699 43064 22744 43092
rect 22738 43052 22744 43064
rect 22796 43052 22802 43104
rect 25130 43092 25136 43104
rect 25091 43064 25136 43092
rect 25130 43052 25136 43064
rect 25188 43052 25194 43104
rect 25866 43092 25872 43104
rect 25827 43064 25872 43092
rect 25866 43052 25872 43064
rect 25924 43052 25930 43104
rect 27890 43052 27896 43104
rect 27948 43092 27954 43104
rect 29181 43095 29239 43101
rect 29181 43092 29193 43095
rect 27948 43064 29193 43092
rect 27948 43052 27954 43064
rect 29181 43061 29193 43064
rect 29227 43061 29239 43095
rect 29181 43055 29239 43061
rect 57241 43095 57299 43101
rect 57241 43061 57253 43095
rect 57287 43092 57299 43095
rect 57698 43092 57704 43104
rect 57287 43064 57704 43092
rect 57287 43061 57299 43064
rect 57241 43055 57299 43061
rect 57698 43052 57704 43064
rect 57756 43052 57762 43104
rect 1104 43002 58880 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 58880 43002
rect 1104 42928 58880 42950
rect 20441 42891 20499 42897
rect 20441 42857 20453 42891
rect 20487 42888 20499 42891
rect 21174 42888 21180 42900
rect 20487 42860 21180 42888
rect 20487 42857 20499 42860
rect 20441 42851 20499 42857
rect 21174 42848 21180 42860
rect 21232 42848 21238 42900
rect 23293 42891 23351 42897
rect 23293 42857 23305 42891
rect 23339 42857 23351 42891
rect 23293 42851 23351 42857
rect 22180 42823 22238 42829
rect 22180 42789 22192 42823
rect 22226 42820 22238 42823
rect 22554 42820 22560 42832
rect 22226 42792 22560 42820
rect 22226 42789 22238 42792
rect 22180 42783 22238 42789
rect 22554 42780 22560 42792
rect 22612 42780 22618 42832
rect 23308 42820 23336 42851
rect 23658 42848 23664 42900
rect 23716 42888 23722 42900
rect 23842 42888 23848 42900
rect 23716 42860 23848 42888
rect 23716 42848 23722 42860
rect 23842 42848 23848 42860
rect 23900 42888 23906 42900
rect 23958 42891 24016 42897
rect 23958 42888 23970 42891
rect 23900 42860 23970 42888
rect 23900 42848 23906 42860
rect 23958 42857 23970 42860
rect 24004 42857 24016 42891
rect 26602 42888 26608 42900
rect 26563 42860 26608 42888
rect 23958 42851 24016 42857
rect 26602 42848 26608 42860
rect 26660 42848 26666 42900
rect 27154 42888 27160 42900
rect 27115 42860 27160 42888
rect 27154 42848 27160 42860
rect 27212 42848 27218 42900
rect 27982 42888 27988 42900
rect 27943 42860 27988 42888
rect 27982 42848 27988 42860
rect 28040 42848 28046 42900
rect 57974 42848 57980 42900
rect 58032 42888 58038 42900
rect 58161 42891 58219 42897
rect 58161 42888 58173 42891
rect 58032 42860 58173 42888
rect 58032 42848 58038 42860
rect 58161 42857 58173 42860
rect 58207 42857 58219 42891
rect 58161 42851 58219 42857
rect 23382 42820 23388 42832
rect 23308 42792 23388 42820
rect 23382 42780 23388 42792
rect 23440 42820 23446 42832
rect 23753 42823 23811 42829
rect 23753 42820 23765 42823
rect 23440 42792 23765 42820
rect 23440 42780 23446 42792
rect 23753 42789 23765 42792
rect 23799 42789 23811 42823
rect 23753 42783 23811 42789
rect 25492 42823 25550 42829
rect 25492 42789 25504 42823
rect 25538 42820 25550 42823
rect 25866 42820 25872 42832
rect 25538 42792 25872 42820
rect 25538 42789 25550 42792
rect 25492 42783 25550 42789
rect 25866 42780 25872 42792
rect 25924 42780 25930 42832
rect 1394 42752 1400 42764
rect 1355 42724 1400 42752
rect 1394 42712 1400 42724
rect 1452 42712 1458 42764
rect 20438 42755 20496 42761
rect 20438 42721 20450 42755
rect 20484 42752 20496 42755
rect 20901 42755 20959 42761
rect 20901 42752 20913 42755
rect 20484 42724 20913 42752
rect 20484 42721 20496 42724
rect 20438 42715 20496 42721
rect 20901 42721 20913 42724
rect 20947 42752 20959 42755
rect 21082 42752 21088 42764
rect 20947 42724 21088 42752
rect 20947 42721 20959 42724
rect 20901 42715 20959 42721
rect 21082 42712 21088 42724
rect 21140 42712 21146 42764
rect 21913 42755 21971 42761
rect 21913 42721 21925 42755
rect 21959 42752 21971 42755
rect 22646 42752 22652 42764
rect 21959 42724 22652 42752
rect 21959 42721 21971 42724
rect 21913 42715 21971 42721
rect 22646 42712 22652 42724
rect 22704 42712 22710 42764
rect 25222 42752 25228 42764
rect 25183 42724 25228 42752
rect 25222 42712 25228 42724
rect 25280 42712 25286 42764
rect 26620 42752 26648 42848
rect 27065 42755 27123 42761
rect 27065 42752 27077 42755
rect 26620 42724 27077 42752
rect 27065 42721 27077 42724
rect 27111 42721 27123 42755
rect 27065 42715 27123 42721
rect 27522 42712 27528 42764
rect 27580 42752 27586 42764
rect 28169 42755 28227 42761
rect 28169 42752 28181 42755
rect 27580 42724 28181 42752
rect 27580 42712 27586 42724
rect 28169 42721 28181 42724
rect 28215 42721 28227 42755
rect 28169 42715 28227 42721
rect 28353 42755 28411 42761
rect 28353 42721 28365 42755
rect 28399 42752 28411 42755
rect 29086 42752 29092 42764
rect 28399 42724 29092 42752
rect 28399 42721 28411 42724
rect 28353 42715 28411 42721
rect 29086 42712 29092 42724
rect 29144 42712 29150 42764
rect 29181 42755 29239 42761
rect 29181 42721 29193 42755
rect 29227 42721 29239 42755
rect 29181 42715 29239 42721
rect 29365 42755 29423 42761
rect 29365 42721 29377 42755
rect 29411 42752 29423 42755
rect 29546 42752 29552 42764
rect 29411 42724 29552 42752
rect 29411 42721 29423 42724
rect 29365 42715 29423 42721
rect 20809 42687 20867 42693
rect 20809 42653 20821 42687
rect 20855 42684 20867 42687
rect 21174 42684 21180 42696
rect 20855 42656 21180 42684
rect 20855 42653 20867 42656
rect 20809 42647 20867 42653
rect 21174 42644 21180 42656
rect 21232 42644 21238 42696
rect 27890 42644 27896 42696
rect 27948 42684 27954 42696
rect 28445 42687 28503 42693
rect 28445 42684 28457 42687
rect 27948 42656 28457 42684
rect 27948 42644 27954 42656
rect 28445 42653 28457 42656
rect 28491 42653 28503 42687
rect 29196 42684 29224 42715
rect 29546 42712 29552 42724
rect 29604 42712 29610 42764
rect 30466 42752 30472 42764
rect 30427 42724 30472 42752
rect 30466 42712 30472 42724
rect 30524 42712 30530 42764
rect 30650 42712 30656 42764
rect 30708 42752 30714 42764
rect 31297 42755 31355 42761
rect 31297 42752 31309 42755
rect 30708 42724 31309 42752
rect 30708 42712 30714 42724
rect 31297 42721 31309 42724
rect 31343 42721 31355 42755
rect 31941 42755 31999 42761
rect 31941 42752 31953 42755
rect 31297 42715 31355 42721
rect 31726 42724 31953 42752
rect 29196 42656 30604 42684
rect 28445 42647 28503 42653
rect 25130 42616 25136 42628
rect 23952 42588 25136 42616
rect 20254 42548 20260 42560
rect 20215 42520 20260 42548
rect 20254 42508 20260 42520
rect 20312 42508 20318 42560
rect 23566 42508 23572 42560
rect 23624 42548 23630 42560
rect 23952 42557 23980 42588
rect 25130 42576 25136 42588
rect 25188 42576 25194 42628
rect 23937 42551 23995 42557
rect 23937 42548 23949 42551
rect 23624 42520 23949 42548
rect 23624 42508 23630 42520
rect 23937 42517 23949 42520
rect 23983 42517 23995 42551
rect 23937 42511 23995 42517
rect 24121 42551 24179 42557
rect 24121 42517 24133 42551
rect 24167 42548 24179 42551
rect 24486 42548 24492 42560
rect 24167 42520 24492 42548
rect 24167 42517 24179 42520
rect 24121 42511 24179 42517
rect 24486 42508 24492 42520
rect 24544 42508 24550 42560
rect 28442 42508 28448 42560
rect 28500 42548 28506 42560
rect 30576 42557 30604 42656
rect 31726 42616 31754 42724
rect 31941 42721 31953 42724
rect 31987 42721 31999 42755
rect 31941 42715 31999 42721
rect 32493 42755 32551 42761
rect 32493 42721 32505 42755
rect 32539 42721 32551 42755
rect 32493 42715 32551 42721
rect 32677 42755 32735 42761
rect 32677 42721 32689 42755
rect 32723 42752 32735 42755
rect 32858 42752 32864 42764
rect 32723 42724 32864 42752
rect 32723 42721 32735 42724
rect 32677 42715 32735 42721
rect 32508 42684 32536 42715
rect 32858 42712 32864 42724
rect 32916 42712 32922 42764
rect 56870 42752 56876 42764
rect 56831 42724 56876 42752
rect 56870 42712 56876 42724
rect 56928 42712 56934 42764
rect 57054 42752 57060 42764
rect 57015 42724 57060 42752
rect 57054 42712 57060 42724
rect 57112 42712 57118 42764
rect 57422 42712 57428 42764
rect 57480 42752 57486 42764
rect 57517 42755 57575 42761
rect 57517 42752 57529 42755
rect 57480 42724 57529 42752
rect 57480 42712 57486 42724
rect 57517 42721 57529 42724
rect 57563 42721 57575 42755
rect 57698 42752 57704 42764
rect 57659 42724 57704 42752
rect 57517 42715 57575 42721
rect 57698 42712 57704 42724
rect 57756 42712 57762 42764
rect 33226 42684 33232 42696
rect 32508 42656 33232 42684
rect 33226 42644 33232 42656
rect 33284 42644 33290 42696
rect 31128 42588 31754 42616
rect 31128 42560 31156 42588
rect 29549 42551 29607 42557
rect 29549 42548 29561 42551
rect 28500 42520 29561 42548
rect 28500 42508 28506 42520
rect 29549 42517 29561 42520
rect 29595 42517 29607 42551
rect 29549 42511 29607 42517
rect 30561 42551 30619 42557
rect 30561 42517 30573 42551
rect 30607 42548 30619 42551
rect 30834 42548 30840 42560
rect 30607 42520 30840 42548
rect 30607 42517 30619 42520
rect 30561 42511 30619 42517
rect 30834 42508 30840 42520
rect 30892 42508 30898 42560
rect 31110 42548 31116 42560
rect 31071 42520 31116 42548
rect 31110 42508 31116 42520
rect 31168 42508 31174 42560
rect 31662 42508 31668 42560
rect 31720 42548 31726 42560
rect 31757 42551 31815 42557
rect 31757 42548 31769 42551
rect 31720 42520 31769 42548
rect 31720 42508 31726 42520
rect 31757 42517 31769 42520
rect 31803 42517 31815 42551
rect 31757 42511 31815 42517
rect 32493 42551 32551 42557
rect 32493 42517 32505 42551
rect 32539 42548 32551 42551
rect 33134 42548 33140 42560
rect 32539 42520 33140 42548
rect 32539 42517 32551 42520
rect 32493 42511 32551 42517
rect 33134 42508 33140 42520
rect 33192 42508 33198 42560
rect 1104 42458 58880 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 58880 42458
rect 1104 42384 58880 42406
rect 20898 42304 20904 42356
rect 20956 42344 20962 42356
rect 21361 42347 21419 42353
rect 21361 42344 21373 42347
rect 20956 42316 21373 42344
rect 20956 42304 20962 42316
rect 21361 42313 21373 42316
rect 21407 42313 21419 42347
rect 24302 42344 24308 42356
rect 24263 42316 24308 42344
rect 21361 42307 21419 42313
rect 24302 42304 24308 42316
rect 24360 42304 24366 42356
rect 24946 42304 24952 42356
rect 25004 42344 25010 42356
rect 25222 42344 25228 42356
rect 25004 42316 25228 42344
rect 25004 42304 25010 42316
rect 25222 42304 25228 42316
rect 25280 42344 25286 42356
rect 25869 42347 25927 42353
rect 25869 42344 25881 42347
rect 25280 42316 25881 42344
rect 25280 42304 25286 42316
rect 25869 42313 25881 42316
rect 25915 42344 25927 42347
rect 26142 42344 26148 42356
rect 25915 42316 26148 42344
rect 25915 42313 25927 42316
rect 25869 42307 25927 42313
rect 26142 42304 26148 42316
rect 26200 42304 26206 42356
rect 26234 42304 26240 42356
rect 26292 42344 26298 42356
rect 26605 42347 26663 42353
rect 26605 42344 26617 42347
rect 26292 42316 26617 42344
rect 26292 42304 26298 42316
rect 26605 42313 26617 42316
rect 26651 42313 26663 42347
rect 26605 42307 26663 42313
rect 28058 42347 28116 42353
rect 28058 42313 28070 42347
rect 28104 42344 28116 42347
rect 28442 42344 28448 42356
rect 28104 42316 28448 42344
rect 28104 42313 28116 42316
rect 28058 42307 28116 42313
rect 28442 42304 28448 42316
rect 28500 42304 28506 42356
rect 30466 42344 30472 42356
rect 30427 42316 30472 42344
rect 30466 42304 30472 42316
rect 30524 42304 30530 42356
rect 23569 42279 23627 42285
rect 23569 42245 23581 42279
rect 23615 42245 23627 42279
rect 26160 42276 26188 42304
rect 27798 42276 27804 42288
rect 26160 42248 27804 42276
rect 23569 42239 23627 42245
rect 21174 42168 21180 42220
rect 21232 42208 21238 42220
rect 23584 42208 23612 42239
rect 27798 42236 27804 42248
rect 27856 42236 27862 42288
rect 28166 42276 28172 42288
rect 28127 42248 28172 42276
rect 28166 42236 28172 42248
rect 28224 42236 28230 42288
rect 30926 42236 30932 42288
rect 30984 42276 30990 42288
rect 31662 42276 31668 42288
rect 30984 42248 31668 42276
rect 30984 42236 30990 42248
rect 31662 42236 31668 42248
rect 31720 42276 31726 42288
rect 31720 42248 33088 42276
rect 31720 42236 31726 42248
rect 28261 42211 28319 42217
rect 21232 42180 21680 42208
rect 23584 42180 24348 42208
rect 21232 42168 21238 42180
rect 1394 42140 1400 42152
rect 1355 42112 1400 42140
rect 1394 42100 1400 42112
rect 1452 42100 1458 42152
rect 19521 42143 19579 42149
rect 19521 42109 19533 42143
rect 19567 42109 19579 42143
rect 19521 42103 19579 42109
rect 19788 42143 19846 42149
rect 19788 42109 19800 42143
rect 19834 42140 19846 42143
rect 20254 42140 20260 42152
rect 19834 42112 20260 42140
rect 19834 42109 19846 42112
rect 19788 42103 19846 42109
rect 19536 42072 19564 42103
rect 20254 42100 20260 42112
rect 20312 42100 20318 42152
rect 21358 42140 21364 42152
rect 21319 42112 21364 42140
rect 21358 42100 21364 42112
rect 21416 42100 21422 42152
rect 21652 42149 21680 42180
rect 21637 42143 21695 42149
rect 21637 42109 21649 42143
rect 21683 42109 21695 42143
rect 21637 42103 21695 42109
rect 23382 42100 23388 42152
rect 23440 42140 23446 42152
rect 23753 42143 23811 42149
rect 23753 42140 23765 42143
rect 23440 42112 23765 42140
rect 23440 42100 23446 42112
rect 23753 42109 23765 42112
rect 23799 42109 23811 42143
rect 23753 42103 23811 42109
rect 23842 42100 23848 42152
rect 23900 42140 23906 42152
rect 24320 42149 24348 42180
rect 28261 42177 28273 42211
rect 28307 42208 28319 42211
rect 28442 42208 28448 42220
rect 28307 42180 28448 42208
rect 28307 42177 28319 42180
rect 28261 42171 28319 42177
rect 28442 42168 28448 42180
rect 28500 42168 28506 42220
rect 32033 42211 32091 42217
rect 32033 42208 32045 42211
rect 31588 42180 32045 42208
rect 24305 42143 24363 42149
rect 23900 42112 23945 42140
rect 23900 42100 23906 42112
rect 24305 42109 24317 42143
rect 24351 42109 24363 42143
rect 24486 42140 24492 42152
rect 24447 42112 24492 42140
rect 24305 42103 24363 42109
rect 24486 42100 24492 42112
rect 24544 42100 24550 42152
rect 24578 42100 24584 42152
rect 24636 42140 24642 42152
rect 24949 42143 25007 42149
rect 24949 42140 24961 42143
rect 24636 42112 24961 42140
rect 24636 42100 24642 42112
rect 24949 42109 24961 42112
rect 24995 42109 25007 42143
rect 24949 42103 25007 42109
rect 26053 42143 26111 42149
rect 26053 42109 26065 42143
rect 26099 42109 26111 42143
rect 26053 42103 26111 42109
rect 20162 42072 20168 42084
rect 19536 42044 20168 42072
rect 20162 42032 20168 42044
rect 20220 42072 20226 42084
rect 20714 42072 20720 42084
rect 20220 42044 20720 42072
rect 20220 42032 20226 42044
rect 20714 42032 20720 42044
rect 20772 42032 20778 42084
rect 23566 42072 23572 42084
rect 23527 42044 23572 42072
rect 23566 42032 23572 42044
rect 23624 42032 23630 42084
rect 20901 42007 20959 42013
rect 20901 41973 20913 42007
rect 20947 42004 20959 42007
rect 21082 42004 21088 42016
rect 20947 41976 21088 42004
rect 20947 41973 20959 41976
rect 20901 41967 20959 41973
rect 21082 41964 21088 41976
rect 21140 42004 21146 42016
rect 21545 42007 21603 42013
rect 21545 42004 21557 42007
rect 21140 41976 21557 42004
rect 21140 41964 21146 41976
rect 21545 41973 21557 41976
rect 21591 41973 21603 42007
rect 21545 41967 21603 41973
rect 25041 42007 25099 42013
rect 25041 41973 25053 42007
rect 25087 42004 25099 42007
rect 25682 42004 25688 42016
rect 25087 41976 25688 42004
rect 25087 41973 25099 41976
rect 25041 41967 25099 41973
rect 25682 41964 25688 41976
rect 25740 41964 25746 42016
rect 26068 42004 26096 42103
rect 26326 42100 26332 42152
rect 26384 42140 26390 42152
rect 26513 42143 26571 42149
rect 26513 42140 26525 42143
rect 26384 42112 26525 42140
rect 26384 42100 26390 42112
rect 26513 42109 26525 42112
rect 26559 42109 26571 42143
rect 26513 42103 26571 42109
rect 28074 42100 28080 42152
rect 28132 42140 28138 42152
rect 28629 42143 28687 42149
rect 28629 42140 28641 42143
rect 28132 42112 28641 42140
rect 28132 42100 28138 42112
rect 28629 42109 28641 42112
rect 28675 42109 28687 42143
rect 28629 42103 28687 42109
rect 28810 42100 28816 42152
rect 28868 42140 28874 42152
rect 29089 42143 29147 42149
rect 29089 42140 29101 42143
rect 28868 42112 29101 42140
rect 28868 42100 28874 42112
rect 29089 42109 29101 42112
rect 29135 42109 29147 42143
rect 29089 42103 29147 42109
rect 29356 42143 29414 42149
rect 29356 42109 29368 42143
rect 29402 42140 29414 42143
rect 29730 42140 29736 42152
rect 29402 42112 29736 42140
rect 29402 42109 29414 42112
rect 29356 42103 29414 42109
rect 29730 42100 29736 42112
rect 29788 42100 29794 42152
rect 27890 42072 27896 42084
rect 27851 42044 27896 42072
rect 27890 42032 27896 42044
rect 27948 42032 27954 42084
rect 31110 42072 31116 42084
rect 28460 42044 31116 42072
rect 28460 42004 28488 42044
rect 31110 42032 31116 42044
rect 31168 42032 31174 42084
rect 31478 42004 31484 42016
rect 26068 41976 28488 42004
rect 31439 41976 31484 42004
rect 31478 41964 31484 41976
rect 31536 41964 31542 42016
rect 31588 42004 31616 42180
rect 32033 42177 32045 42180
rect 32079 42208 32091 42211
rect 32674 42208 32680 42220
rect 32079 42180 32680 42208
rect 32079 42177 32091 42180
rect 32033 42171 32091 42177
rect 32674 42168 32680 42180
rect 32732 42168 32738 42220
rect 33060 42217 33088 42248
rect 33045 42211 33103 42217
rect 33045 42177 33057 42211
rect 33091 42177 33103 42211
rect 33045 42171 33103 42177
rect 31662 42143 31720 42149
rect 31662 42109 31674 42143
rect 31708 42140 31720 42143
rect 32122 42140 32128 42152
rect 31708 42112 32128 42140
rect 31708 42109 31720 42112
rect 31662 42103 31720 42109
rect 32122 42100 32128 42112
rect 32180 42100 32186 42152
rect 33134 42100 33140 42152
rect 33192 42140 33198 42152
rect 33301 42143 33359 42149
rect 33301 42140 33313 42143
rect 33192 42112 33313 42140
rect 33192 42100 33198 42112
rect 33301 42109 33313 42112
rect 33347 42109 33359 42143
rect 33301 42103 33359 42109
rect 56502 42100 56508 42152
rect 56560 42140 56566 42152
rect 56597 42143 56655 42149
rect 56597 42140 56609 42143
rect 56560 42112 56609 42140
rect 56560 42100 56566 42112
rect 56597 42109 56609 42112
rect 56643 42109 56655 42143
rect 56597 42103 56655 42109
rect 57425 42143 57483 42149
rect 57425 42109 57437 42143
rect 57471 42140 57483 42143
rect 57514 42140 57520 42152
rect 57471 42112 57520 42140
rect 57471 42109 57483 42112
rect 57425 42103 57483 42109
rect 57514 42100 57520 42112
rect 57572 42100 57578 42152
rect 57974 42072 57980 42084
rect 57935 42044 57980 42072
rect 57974 42032 57980 42044
rect 58032 42032 58038 42084
rect 58158 42072 58164 42084
rect 58119 42044 58164 42072
rect 58158 42032 58164 42044
rect 58216 42032 58222 42084
rect 31665 42007 31723 42013
rect 31665 42004 31677 42007
rect 31588 41976 31677 42004
rect 31665 41973 31677 41976
rect 31711 41973 31723 42007
rect 31665 41967 31723 41973
rect 33318 41964 33324 42016
rect 33376 42004 33382 42016
rect 34425 42007 34483 42013
rect 34425 42004 34437 42007
rect 33376 41976 34437 42004
rect 33376 41964 33382 41976
rect 34425 41973 34437 41976
rect 34471 41973 34483 42007
rect 34425 41967 34483 41973
rect 1104 41914 58880 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 58880 41914
rect 1104 41840 58880 41862
rect 20901 41803 20959 41809
rect 20901 41769 20913 41803
rect 20947 41800 20959 41803
rect 21174 41800 21180 41812
rect 20947 41772 21180 41800
rect 20947 41769 20959 41772
rect 20901 41763 20959 41769
rect 21174 41760 21180 41772
rect 21232 41760 21238 41812
rect 27709 41803 27767 41809
rect 27709 41769 27721 41803
rect 27755 41769 27767 41803
rect 27709 41763 27767 41769
rect 24210 41732 24216 41744
rect 23860 41704 24216 41732
rect 20806 41664 20812 41676
rect 20767 41636 20812 41664
rect 20806 41624 20812 41636
rect 20864 41624 20870 41676
rect 21174 41624 21180 41676
rect 21232 41664 21238 41676
rect 23860 41673 23888 41704
rect 24210 41692 24216 41704
rect 24268 41732 24274 41744
rect 24578 41732 24584 41744
rect 24268 41704 24584 41732
rect 24268 41692 24274 41704
rect 24578 41692 24584 41704
rect 24636 41692 24642 41744
rect 27724 41732 27752 41763
rect 27798 41760 27804 41812
rect 27856 41800 27862 41812
rect 28810 41800 28816 41812
rect 27856 41772 28816 41800
rect 27856 41760 27862 41772
rect 28810 41760 28816 41772
rect 28868 41800 28874 41812
rect 32033 41803 32091 41809
rect 28868 41772 30052 41800
rect 28868 41760 28874 41772
rect 27724 41704 29408 41732
rect 21709 41667 21767 41673
rect 21709 41664 21721 41667
rect 21232 41636 21721 41664
rect 21232 41624 21238 41636
rect 21709 41633 21721 41636
rect 21755 41633 21767 41667
rect 21709 41627 21767 41633
rect 23845 41667 23903 41673
rect 23845 41633 23857 41667
rect 23891 41633 23903 41667
rect 24026 41664 24032 41676
rect 23939 41636 24032 41664
rect 23845 41627 23903 41633
rect 24026 41624 24032 41636
rect 24084 41664 24090 41676
rect 24486 41664 24492 41676
rect 24084 41636 24492 41664
rect 24084 41624 24090 41636
rect 24486 41624 24492 41636
rect 24544 41624 24550 41676
rect 25498 41664 25504 41676
rect 25459 41636 25504 41664
rect 25498 41624 25504 41636
rect 25556 41624 25562 41676
rect 25682 41664 25688 41676
rect 25643 41636 25688 41664
rect 25682 41624 25688 41636
rect 25740 41624 25746 41676
rect 26142 41624 26148 41676
rect 26200 41664 26206 41676
rect 26329 41667 26387 41673
rect 26329 41664 26341 41667
rect 26200 41636 26341 41664
rect 26200 41624 26206 41636
rect 26329 41633 26341 41636
rect 26375 41633 26387 41667
rect 26329 41627 26387 41633
rect 26596 41667 26654 41673
rect 26596 41633 26608 41667
rect 26642 41664 26654 41667
rect 27798 41664 27804 41676
rect 26642 41636 27804 41664
rect 26642 41633 26654 41636
rect 26596 41627 26654 41633
rect 27798 41624 27804 41636
rect 27856 41624 27862 41676
rect 27890 41624 27896 41676
rect 27948 41664 27954 41676
rect 28074 41664 28080 41676
rect 27948 41636 28080 41664
rect 27948 41624 27954 41636
rect 28074 41624 28080 41636
rect 28132 41664 28138 41676
rect 28169 41667 28227 41673
rect 28169 41664 28181 41667
rect 28132 41636 28181 41664
rect 28132 41624 28138 41636
rect 28169 41633 28181 41636
rect 28215 41633 28227 41667
rect 28442 41664 28448 41676
rect 28355 41636 28448 41664
rect 28169 41627 28227 41633
rect 28442 41624 28448 41636
rect 28500 41664 28506 41676
rect 29380 41673 29408 41704
rect 29365 41667 29423 41673
rect 28500 41636 29040 41664
rect 28500 41624 28506 41636
rect 20714 41556 20720 41608
rect 20772 41596 20778 41608
rect 21453 41599 21511 41605
rect 21453 41596 21465 41599
rect 20772 41568 21465 41596
rect 20772 41556 20778 41568
rect 21453 41565 21465 41568
rect 21499 41565 21511 41599
rect 24118 41596 24124 41608
rect 24079 41568 24124 41596
rect 21453 41559 21511 41565
rect 24118 41556 24124 41568
rect 24176 41556 24182 41608
rect 25777 41599 25835 41605
rect 25777 41565 25789 41599
rect 25823 41596 25835 41599
rect 25866 41596 25872 41608
rect 25823 41568 25872 41596
rect 25823 41565 25835 41568
rect 25777 41559 25835 41565
rect 25866 41556 25872 41568
rect 25924 41556 25930 41608
rect 28902 41596 28908 41608
rect 28863 41568 28908 41596
rect 28902 41556 28908 41568
rect 28960 41556 28966 41608
rect 29012 41596 29040 41636
rect 29365 41633 29377 41667
rect 29411 41633 29423 41667
rect 30024 41664 30052 41772
rect 32033 41769 32045 41803
rect 32079 41800 32091 41803
rect 32122 41800 32128 41812
rect 32079 41772 32128 41800
rect 32079 41769 32091 41772
rect 32033 41763 32091 41769
rect 32122 41760 32128 41772
rect 32180 41800 32186 41812
rect 33505 41803 33563 41809
rect 33505 41800 33517 41803
rect 32180 41772 33517 41800
rect 32180 41760 32186 41772
rect 30920 41735 30978 41741
rect 30920 41701 30932 41735
rect 30966 41732 30978 41735
rect 31478 41732 31484 41744
rect 30966 41704 31484 41732
rect 30966 41701 30978 41704
rect 30920 41695 30978 41701
rect 31478 41692 31484 41704
rect 31536 41692 31542 41744
rect 32508 41741 32536 41772
rect 33505 41769 33517 41772
rect 33551 41769 33563 41803
rect 33505 41763 33563 41769
rect 57974 41760 57980 41812
rect 58032 41800 58038 41812
rect 58161 41803 58219 41809
rect 58161 41800 58173 41803
rect 58032 41772 58173 41800
rect 58032 41760 58038 41772
rect 58161 41769 58173 41772
rect 58207 41769 58219 41803
rect 58161 41763 58219 41769
rect 32493 41735 32551 41741
rect 32493 41701 32505 41735
rect 32539 41701 32551 41735
rect 32493 41695 32551 41701
rect 32674 41692 32680 41744
rect 32732 41741 32738 41744
rect 32732 41735 32756 41741
rect 32744 41701 32756 41735
rect 33318 41732 33324 41744
rect 33279 41704 33324 41732
rect 32732 41695 32756 41701
rect 32732 41692 32738 41695
rect 33318 41692 33324 41704
rect 33376 41692 33382 41744
rect 30653 41667 30711 41673
rect 30653 41664 30665 41667
rect 30024 41636 30665 41664
rect 29365 41627 29423 41633
rect 30653 41633 30665 41636
rect 30699 41633 30711 41667
rect 33336 41664 33364 41692
rect 30653 41627 30711 41633
rect 32692 41636 33364 41664
rect 33597 41667 33655 41673
rect 29457 41599 29515 41605
rect 29457 41596 29469 41599
rect 29012 41568 29469 41596
rect 29457 41565 29469 41568
rect 29503 41565 29515 41599
rect 29457 41559 29515 41565
rect 28166 41488 28172 41540
rect 28224 41528 28230 41540
rect 28261 41531 28319 41537
rect 28261 41528 28273 41531
rect 28224 41500 28273 41528
rect 28224 41488 28230 41500
rect 28261 41497 28273 41500
rect 28307 41497 28319 41531
rect 28261 41491 28319 41497
rect 22370 41420 22376 41472
rect 22428 41460 22434 41472
rect 22833 41463 22891 41469
rect 22833 41460 22845 41463
rect 22428 41432 22845 41460
rect 22428 41420 22434 41432
rect 22833 41429 22845 41432
rect 22879 41429 22891 41463
rect 23658 41460 23664 41472
rect 23619 41432 23664 41460
rect 22833 41423 22891 41429
rect 23658 41420 23664 41432
rect 23716 41420 23722 41472
rect 25222 41420 25228 41472
rect 25280 41460 25286 41472
rect 32692 41469 32720 41636
rect 33597 41633 33609 41667
rect 33643 41633 33655 41667
rect 57054 41664 57060 41676
rect 57015 41636 57060 41664
rect 33597 41627 33655 41633
rect 33042 41556 33048 41608
rect 33100 41596 33106 41608
rect 33612 41596 33640 41627
rect 57054 41624 57060 41636
rect 57112 41664 57118 41676
rect 57330 41664 57336 41676
rect 57112 41636 57336 41664
rect 57112 41624 57118 41636
rect 57330 41624 57336 41636
rect 57388 41624 57394 41676
rect 57514 41664 57520 41676
rect 57475 41636 57520 41664
rect 57514 41624 57520 41636
rect 57572 41624 57578 41676
rect 57701 41599 57759 41605
rect 57701 41596 57713 41599
rect 33100 41568 33640 41596
rect 56888 41568 57713 41596
rect 33100 41556 33106 41568
rect 32858 41528 32864 41540
rect 32819 41500 32864 41528
rect 32858 41488 32864 41500
rect 32916 41488 32922 41540
rect 33226 41488 33232 41540
rect 33284 41528 33290 41540
rect 56888 41537 56916 41568
rect 57701 41565 57713 41568
rect 57747 41565 57759 41599
rect 57701 41559 57759 41565
rect 33321 41531 33379 41537
rect 33321 41528 33333 41531
rect 33284 41500 33333 41528
rect 33284 41488 33290 41500
rect 33321 41497 33333 41500
rect 33367 41497 33379 41531
rect 33321 41491 33379 41497
rect 56873 41531 56931 41537
rect 56873 41497 56885 41531
rect 56919 41497 56931 41531
rect 56873 41491 56931 41497
rect 25317 41463 25375 41469
rect 25317 41460 25329 41463
rect 25280 41432 25329 41460
rect 25280 41420 25286 41432
rect 25317 41429 25329 41432
rect 25363 41429 25375 41463
rect 25317 41423 25375 41429
rect 32677 41463 32735 41469
rect 32677 41429 32689 41463
rect 32723 41429 32735 41463
rect 32677 41423 32735 41429
rect 1104 41370 58880 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 58880 41370
rect 1104 41296 58880 41318
rect 21174 41256 21180 41268
rect 21135 41228 21180 41256
rect 21174 41216 21180 41228
rect 21232 41216 21238 41268
rect 24118 41216 24124 41268
rect 24176 41256 24182 41268
rect 24489 41259 24547 41265
rect 24489 41256 24501 41259
rect 24176 41228 24501 41256
rect 24176 41216 24182 41228
rect 24489 41225 24501 41228
rect 24535 41225 24547 41259
rect 24489 41219 24547 41225
rect 25866 41216 25872 41268
rect 25924 41256 25930 41268
rect 26329 41259 26387 41265
rect 26329 41256 26341 41259
rect 25924 41228 26341 41256
rect 25924 41216 25930 41228
rect 26329 41225 26341 41228
rect 26375 41225 26387 41259
rect 27798 41256 27804 41268
rect 27759 41228 27804 41256
rect 26329 41219 26387 41225
rect 27798 41216 27804 41228
rect 27856 41216 27862 41268
rect 30558 41216 30564 41268
rect 30616 41256 30622 41268
rect 30653 41259 30711 41265
rect 30653 41256 30665 41259
rect 30616 41228 30665 41256
rect 30616 41216 30622 41228
rect 30653 41225 30665 41228
rect 30699 41225 30711 41259
rect 57330 41256 57336 41268
rect 57291 41228 57336 41256
rect 30653 41219 30711 41225
rect 57330 41216 57336 41228
rect 57388 41216 57394 41268
rect 22646 41080 22652 41132
rect 22704 41120 22710 41132
rect 23109 41123 23167 41129
rect 23109 41120 23121 41123
rect 22704 41092 23121 41120
rect 22704 41080 22710 41092
rect 23109 41089 23121 41092
rect 23155 41089 23167 41123
rect 28810 41120 28816 41132
rect 28771 41092 28816 41120
rect 23109 41083 23167 41089
rect 28810 41080 28816 41092
rect 28868 41080 28874 41132
rect 29822 41080 29828 41132
rect 29880 41120 29886 41132
rect 31021 41123 31079 41129
rect 31021 41120 31033 41123
rect 29880 41092 31033 41120
rect 29880 41080 29886 41092
rect 31021 41089 31033 41092
rect 31067 41089 31079 41123
rect 31021 41083 31079 41089
rect 1394 41052 1400 41064
rect 1355 41024 1400 41052
rect 1394 41012 1400 41024
rect 1452 41012 1458 41064
rect 20806 41012 20812 41064
rect 20864 41052 20870 41064
rect 21361 41055 21419 41061
rect 21361 41052 21373 41055
rect 20864 41024 21373 41052
rect 20864 41012 20870 41024
rect 21361 41021 21373 41024
rect 21407 41021 21419 41055
rect 21542 41052 21548 41064
rect 21503 41024 21548 41052
rect 21361 41015 21419 41021
rect 21376 40984 21404 41015
rect 21542 41012 21548 41024
rect 21600 41012 21606 41064
rect 21637 41055 21695 41061
rect 21637 41021 21649 41055
rect 21683 41052 21695 41055
rect 22370 41052 22376 41064
rect 21683 41024 22376 41052
rect 21683 41021 21695 41024
rect 21637 41015 21695 41021
rect 22370 41012 22376 41024
rect 22428 41012 22434 41064
rect 23376 41055 23434 41061
rect 23376 41021 23388 41055
rect 23422 41052 23434 41055
rect 23658 41052 23664 41064
rect 23422 41024 23664 41052
rect 23422 41021 23434 41024
rect 23376 41015 23434 41021
rect 23658 41012 23664 41024
rect 23716 41012 23722 41064
rect 24946 41052 24952 41064
rect 24859 41024 24952 41052
rect 24946 41012 24952 41024
rect 25004 41012 25010 41064
rect 25222 41061 25228 41064
rect 25216 41015 25228 41061
rect 25280 41052 25286 41064
rect 25280 41024 25316 41052
rect 25222 41012 25228 41015
rect 25280 41012 25286 41024
rect 27614 41012 27620 41064
rect 27672 41052 27678 41064
rect 28074 41052 28080 41064
rect 27672 41024 28080 41052
rect 27672 41012 27678 41024
rect 28074 41012 28080 41024
rect 28132 41012 28138 41064
rect 28902 41012 28908 41064
rect 28960 41052 28966 41064
rect 29840 41052 29868 41080
rect 30834 41052 30840 41064
rect 28960 41024 29868 41052
rect 30795 41024 30840 41052
rect 28960 41012 28966 41024
rect 30834 41012 30840 41024
rect 30892 41012 30898 41064
rect 31113 41055 31171 41061
rect 31113 41021 31125 41055
rect 31159 41021 31171 41055
rect 31113 41015 31171 41021
rect 21726 40984 21732 40996
rect 21376 40956 21732 40984
rect 21726 40944 21732 40956
rect 21784 40944 21790 40996
rect 24964 40984 24992 41012
rect 25406 40984 25412 40996
rect 24964 40956 25412 40984
rect 25406 40944 25412 40956
rect 25464 40944 25470 40996
rect 27798 40984 27804 40996
rect 27759 40956 27804 40984
rect 27798 40944 27804 40956
rect 27856 40944 27862 40996
rect 27982 40944 27988 40996
rect 28040 40984 28046 40996
rect 28442 40984 28448 40996
rect 28040 40956 28448 40984
rect 28040 40944 28046 40956
rect 28442 40944 28448 40956
rect 28500 40944 28506 40996
rect 28994 40944 29000 40996
rect 29052 40993 29058 40996
rect 29052 40987 29116 40993
rect 29052 40953 29070 40987
rect 29104 40953 29116 40987
rect 29052 40947 29116 40953
rect 29052 40944 29058 40947
rect 29546 40944 29552 40996
rect 29604 40984 29610 40996
rect 31128 40984 31156 41015
rect 31754 41012 31760 41064
rect 31812 41052 31818 41064
rect 31849 41055 31907 41061
rect 31849 41052 31861 41055
rect 31812 41024 31861 41052
rect 31812 41012 31818 41024
rect 31849 41021 31861 41024
rect 31895 41021 31907 41055
rect 31849 41015 31907 41021
rect 32582 41012 32588 41064
rect 32640 41052 32646 41064
rect 33045 41055 33103 41061
rect 33045 41052 33057 41055
rect 32640 41024 33057 41052
rect 32640 41012 32646 41024
rect 33045 41021 33057 41024
rect 33091 41021 33103 41055
rect 33045 41015 33103 41021
rect 33134 41012 33140 41064
rect 33192 41052 33198 41064
rect 33229 41055 33287 41061
rect 33229 41052 33241 41055
rect 33192 41024 33241 41052
rect 33192 41012 33198 41024
rect 33229 41021 33241 41024
rect 33275 41021 33287 41055
rect 56502 41052 56508 41064
rect 56463 41024 56508 41052
rect 33229 41015 33287 41021
rect 56502 41012 56508 41024
rect 56560 41012 56566 41064
rect 29604 40956 31156 40984
rect 57241 40987 57299 40993
rect 29604 40944 29610 40956
rect 57241 40953 57253 40987
rect 57287 40984 57299 40987
rect 57514 40984 57520 40996
rect 57287 40956 57520 40984
rect 57287 40953 57299 40956
rect 57241 40947 57299 40953
rect 57514 40944 57520 40956
rect 57572 40944 57578 40996
rect 57974 40984 57980 40996
rect 57935 40956 57980 40984
rect 57974 40944 57980 40956
rect 58032 40944 58038 40996
rect 58158 40984 58164 40996
rect 58119 40956 58164 40984
rect 58158 40944 58164 40956
rect 58216 40944 58222 40996
rect 30190 40916 30196 40928
rect 30151 40888 30196 40916
rect 30190 40876 30196 40888
rect 30248 40876 30254 40928
rect 31846 40876 31852 40928
rect 31904 40916 31910 40928
rect 31941 40919 31999 40925
rect 31941 40916 31953 40919
rect 31904 40888 31953 40916
rect 31904 40876 31910 40888
rect 31941 40885 31953 40888
rect 31987 40885 31999 40919
rect 33134 40916 33140 40928
rect 33095 40888 33140 40916
rect 31941 40879 31999 40885
rect 33134 40876 33140 40888
rect 33192 40876 33198 40928
rect 1104 40826 58880 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 58880 40826
rect 1104 40752 58880 40774
rect 21542 40672 21548 40724
rect 21600 40712 21606 40724
rect 21637 40715 21695 40721
rect 21637 40712 21649 40715
rect 21600 40684 21649 40712
rect 21600 40672 21606 40684
rect 21637 40681 21649 40684
rect 21683 40681 21695 40715
rect 21637 40675 21695 40681
rect 20070 40644 20076 40656
rect 18800 40616 20076 40644
rect 15105 40579 15163 40585
rect 15105 40545 15117 40579
rect 15151 40576 15163 40579
rect 15194 40576 15200 40588
rect 15151 40548 15200 40576
rect 15151 40545 15163 40548
rect 15105 40539 15163 40545
rect 15194 40536 15200 40548
rect 15252 40536 15258 40588
rect 15286 40536 15292 40588
rect 15344 40576 15350 40588
rect 18800 40585 18828 40616
rect 20070 40604 20076 40616
rect 20128 40604 20134 40656
rect 18785 40579 18843 40585
rect 15344 40548 15389 40576
rect 15344 40536 15350 40548
rect 18785 40545 18797 40579
rect 18831 40545 18843 40579
rect 18785 40539 18843 40545
rect 18969 40579 19027 40585
rect 18969 40545 18981 40579
rect 19015 40576 19027 40579
rect 19978 40576 19984 40588
rect 19015 40548 19984 40576
rect 19015 40545 19027 40548
rect 18969 40539 19027 40545
rect 19978 40536 19984 40548
rect 20036 40536 20042 40588
rect 20165 40579 20223 40585
rect 20165 40545 20177 40579
rect 20211 40545 20223 40579
rect 20165 40539 20223 40545
rect 20809 40579 20867 40585
rect 20809 40545 20821 40579
rect 20855 40576 20867 40579
rect 20898 40576 20904 40588
rect 20855 40548 20904 40576
rect 20855 40545 20867 40548
rect 20809 40539 20867 40545
rect 19061 40511 19119 40517
rect 19061 40477 19073 40511
rect 19107 40508 19119 40511
rect 19702 40508 19708 40520
rect 19107 40480 19708 40508
rect 19107 40477 19119 40480
rect 19061 40471 19119 40477
rect 19702 40468 19708 40480
rect 19760 40508 19766 40520
rect 20180 40508 20208 40539
rect 20898 40536 20904 40548
rect 20956 40576 20962 40588
rect 21545 40579 21603 40585
rect 21545 40576 21557 40579
rect 20956 40548 21557 40576
rect 20956 40536 20962 40548
rect 21545 40545 21557 40548
rect 21591 40545 21603 40579
rect 21652 40576 21680 40675
rect 21726 40672 21732 40724
rect 21784 40712 21790 40724
rect 22281 40715 22339 40721
rect 22281 40712 22293 40715
rect 21784 40684 22293 40712
rect 21784 40672 21790 40684
rect 22281 40681 22293 40684
rect 22327 40681 22339 40715
rect 24210 40712 24216 40724
rect 24171 40684 24216 40712
rect 22281 40675 22339 40681
rect 24210 40672 24216 40684
rect 24268 40672 24274 40724
rect 28994 40712 29000 40724
rect 28955 40684 29000 40712
rect 28994 40672 29000 40684
rect 29052 40672 29058 40724
rect 32582 40712 32588 40724
rect 32543 40684 32588 40712
rect 32582 40672 32588 40684
rect 32640 40672 32646 40724
rect 57974 40672 57980 40724
rect 58032 40712 58038 40724
rect 58161 40715 58219 40721
rect 58161 40712 58173 40715
rect 58032 40684 58173 40712
rect 58032 40672 58038 40684
rect 58161 40681 58173 40684
rect 58207 40681 58219 40715
rect 58161 40675 58219 40681
rect 27982 40644 27988 40656
rect 27080 40616 27988 40644
rect 22189 40579 22247 40585
rect 22189 40576 22201 40579
rect 21652 40548 22201 40576
rect 21545 40539 21603 40545
rect 22189 40545 22201 40548
rect 22235 40545 22247 40579
rect 22370 40576 22376 40588
rect 22331 40548 22376 40576
rect 22189 40539 22247 40545
rect 22370 40536 22376 40548
rect 22428 40536 22434 40588
rect 24026 40576 24032 40588
rect 23987 40548 24032 40576
rect 24026 40536 24032 40548
rect 24084 40536 24090 40588
rect 24118 40536 24124 40588
rect 24176 40576 24182 40588
rect 24213 40579 24271 40585
rect 24213 40576 24225 40579
rect 24176 40548 24225 40576
rect 24176 40536 24182 40548
rect 24213 40545 24225 40548
rect 24259 40545 24271 40579
rect 25682 40576 25688 40588
rect 25643 40548 25688 40576
rect 24213 40539 24271 40545
rect 25682 40536 25688 40548
rect 25740 40536 25746 40588
rect 25866 40576 25872 40588
rect 25827 40548 25872 40576
rect 25866 40536 25872 40548
rect 25924 40536 25930 40588
rect 27080 40585 27108 40616
rect 27982 40604 27988 40616
rect 28040 40604 28046 40656
rect 30190 40644 30196 40656
rect 29196 40616 30196 40644
rect 26881 40579 26939 40585
rect 26881 40545 26893 40579
rect 26927 40545 26939 40579
rect 26881 40539 26939 40545
rect 27065 40579 27123 40585
rect 27065 40545 27077 40579
rect 27111 40545 27123 40579
rect 27065 40539 27123 40545
rect 27709 40579 27767 40585
rect 27709 40545 27721 40579
rect 27755 40576 27767 40579
rect 28902 40576 28908 40588
rect 27755 40548 28908 40576
rect 27755 40545 27767 40548
rect 27709 40539 27767 40545
rect 21082 40508 21088 40520
rect 19760 40480 20208 40508
rect 21043 40480 21088 40508
rect 19760 40468 19766 40480
rect 21082 40468 21088 40480
rect 21140 40468 21146 40520
rect 26896 40508 26924 40539
rect 28902 40536 28908 40548
rect 28960 40536 28966 40588
rect 29196 40585 29224 40616
rect 30190 40604 30196 40616
rect 30248 40644 30254 40656
rect 33505 40647 33563 40653
rect 33505 40644 33517 40647
rect 30248 40616 30512 40644
rect 30248 40604 30254 40616
rect 29181 40579 29239 40585
rect 29181 40545 29193 40579
rect 29227 40545 29239 40579
rect 29181 40539 29239 40545
rect 29270 40536 29276 40588
rect 29328 40576 29334 40588
rect 29546 40576 29552 40588
rect 29328 40548 29373 40576
rect 29507 40548 29552 40576
rect 29328 40536 29334 40548
rect 29546 40536 29552 40548
rect 29604 40536 29610 40588
rect 30484 40585 30512 40616
rect 32784 40616 33517 40644
rect 30469 40579 30527 40585
rect 30469 40545 30481 40579
rect 30515 40545 30527 40579
rect 30469 40539 30527 40545
rect 31481 40579 31539 40585
rect 31481 40545 31493 40579
rect 31527 40545 31539 40579
rect 31481 40539 31539 40545
rect 27614 40508 27620 40520
rect 25700 40480 27620 40508
rect 25498 40400 25504 40452
rect 25556 40440 25562 40452
rect 25700 40449 25728 40480
rect 27614 40468 27620 40480
rect 27672 40468 27678 40520
rect 27982 40508 27988 40520
rect 27943 40480 27988 40508
rect 27982 40468 27988 40480
rect 28040 40468 28046 40520
rect 29564 40508 29592 40536
rect 30561 40511 30619 40517
rect 30561 40508 30573 40511
rect 29564 40480 30573 40508
rect 30561 40477 30573 40480
rect 30607 40477 30619 40511
rect 31496 40508 31524 40539
rect 31570 40536 31576 40588
rect 31628 40576 31634 40588
rect 31846 40576 31852 40588
rect 31628 40548 31673 40576
rect 31807 40548 31852 40576
rect 31628 40536 31634 40548
rect 31846 40536 31852 40548
rect 31904 40536 31910 40588
rect 32784 40585 32812 40616
rect 33505 40613 33517 40616
rect 33551 40644 33563 40647
rect 34054 40644 34060 40656
rect 33551 40616 34060 40644
rect 33551 40613 33563 40616
rect 33505 40607 33563 40613
rect 34054 40604 34060 40616
rect 34112 40604 34118 40656
rect 32769 40579 32827 40585
rect 32769 40545 32781 40579
rect 32815 40545 32827 40579
rect 32769 40539 32827 40545
rect 33689 40579 33747 40585
rect 33689 40545 33701 40579
rect 33735 40545 33747 40579
rect 57054 40576 57060 40588
rect 57015 40548 57060 40576
rect 33689 40539 33747 40545
rect 31754 40508 31760 40520
rect 31496 40480 31760 40508
rect 30561 40471 30619 40477
rect 31754 40468 31760 40480
rect 31812 40468 31818 40520
rect 31864 40508 31892 40536
rect 33045 40511 33103 40517
rect 33045 40508 33057 40511
rect 31864 40480 33057 40508
rect 33045 40477 33057 40480
rect 33091 40508 33103 40511
rect 33704 40508 33732 40539
rect 57054 40536 57060 40548
rect 57112 40536 57118 40588
rect 33091 40480 33732 40508
rect 33091 40477 33103 40480
rect 33045 40471 33103 40477
rect 57422 40468 57428 40520
rect 57480 40508 57486 40520
rect 57517 40511 57575 40517
rect 57517 40508 57529 40511
rect 57480 40480 57529 40508
rect 57480 40468 57486 40480
rect 57517 40477 57529 40480
rect 57563 40477 57575 40511
rect 57517 40471 57575 40477
rect 57701 40511 57759 40517
rect 57701 40477 57713 40511
rect 57747 40477 57759 40511
rect 57701 40471 57759 40477
rect 25685 40443 25743 40449
rect 25685 40440 25697 40443
rect 25556 40412 25697 40440
rect 25556 40400 25562 40412
rect 25685 40409 25697 40412
rect 25731 40409 25743 40443
rect 25685 40403 25743 40409
rect 26881 40443 26939 40449
rect 26881 40409 26893 40443
rect 26927 40440 26939 40443
rect 27798 40440 27804 40452
rect 26927 40412 27804 40440
rect 26927 40409 26939 40412
rect 26881 40403 26939 40409
rect 27798 40400 27804 40412
rect 27856 40440 27862 40452
rect 27893 40443 27951 40449
rect 27893 40440 27905 40443
rect 27856 40412 27905 40440
rect 27856 40400 27862 40412
rect 27893 40409 27905 40412
rect 27939 40409 27951 40443
rect 27893 40403 27951 40409
rect 29457 40443 29515 40449
rect 29457 40409 29469 40443
rect 29503 40440 29515 40443
rect 29822 40440 29828 40452
rect 29503 40412 29828 40440
rect 29503 40409 29515 40412
rect 29457 40403 29515 40409
rect 29822 40400 29828 40412
rect 29880 40400 29886 40452
rect 56873 40443 56931 40449
rect 56873 40409 56885 40443
rect 56919 40440 56931 40443
rect 57716 40440 57744 40471
rect 56919 40412 57744 40440
rect 56919 40409 56931 40412
rect 56873 40403 56931 40409
rect 15105 40375 15163 40381
rect 15105 40341 15117 40375
rect 15151 40372 15163 40375
rect 15378 40372 15384 40384
rect 15151 40344 15384 40372
rect 15151 40341 15163 40344
rect 15105 40335 15163 40341
rect 15378 40332 15384 40344
rect 15436 40332 15442 40384
rect 18598 40372 18604 40384
rect 18559 40344 18604 40372
rect 18598 40332 18604 40344
rect 18656 40332 18662 40384
rect 20438 40332 20444 40384
rect 20496 40372 20502 40384
rect 20625 40375 20683 40381
rect 20625 40372 20637 40375
rect 20496 40344 20637 40372
rect 20496 40332 20502 40344
rect 20625 40341 20637 40344
rect 20671 40341 20683 40375
rect 20625 40335 20683 40341
rect 20806 40332 20812 40384
rect 20864 40372 20870 40384
rect 20993 40375 21051 40381
rect 20993 40372 21005 40375
rect 20864 40344 21005 40372
rect 20864 40332 20870 40344
rect 20993 40341 21005 40344
rect 21039 40341 21051 40375
rect 20993 40335 21051 40341
rect 27525 40375 27583 40381
rect 27525 40341 27537 40375
rect 27571 40372 27583 40375
rect 27706 40372 27712 40384
rect 27571 40344 27712 40372
rect 27571 40341 27583 40344
rect 27525 40335 27583 40341
rect 27706 40332 27712 40344
rect 27764 40332 27770 40384
rect 31294 40372 31300 40384
rect 31255 40344 31300 40372
rect 31294 40332 31300 40344
rect 31352 40332 31358 40384
rect 31757 40375 31815 40381
rect 31757 40341 31769 40375
rect 31803 40372 31815 40375
rect 31846 40372 31852 40384
rect 31803 40344 31852 40372
rect 31803 40341 31815 40344
rect 31757 40335 31815 40341
rect 31846 40332 31852 40344
rect 31904 40372 31910 40384
rect 32953 40375 33011 40381
rect 32953 40372 32965 40375
rect 31904 40344 32965 40372
rect 31904 40332 31910 40344
rect 32953 40341 32965 40344
rect 32999 40341 33011 40375
rect 33870 40372 33876 40384
rect 33831 40344 33876 40372
rect 32953 40335 33011 40341
rect 33870 40332 33876 40344
rect 33928 40332 33934 40384
rect 1104 40282 58880 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 58880 40282
rect 1104 40208 58880 40230
rect 19702 40168 19708 40180
rect 19663 40140 19708 40168
rect 19702 40128 19708 40140
rect 19760 40128 19766 40180
rect 21082 40128 21088 40180
rect 21140 40168 21146 40180
rect 21545 40171 21603 40177
rect 21545 40168 21557 40171
rect 21140 40140 21557 40168
rect 21140 40128 21146 40140
rect 21545 40137 21557 40140
rect 21591 40137 21603 40171
rect 21545 40131 21603 40137
rect 29270 40128 29276 40180
rect 29328 40168 29334 40180
rect 29733 40171 29791 40177
rect 29733 40168 29745 40171
rect 29328 40140 29745 40168
rect 29328 40128 29334 40140
rect 29733 40137 29745 40140
rect 29779 40137 29791 40171
rect 29733 40131 29791 40137
rect 31754 40128 31760 40180
rect 31812 40168 31818 40180
rect 31849 40171 31907 40177
rect 31849 40168 31861 40171
rect 31812 40140 31861 40168
rect 31812 40128 31818 40140
rect 31849 40137 31861 40140
rect 31895 40137 31907 40171
rect 57422 40168 57428 40180
rect 57383 40140 57428 40168
rect 31849 40131 31907 40137
rect 57422 40128 57428 40140
rect 57480 40128 57486 40180
rect 14737 40103 14795 40109
rect 14737 40069 14749 40103
rect 14783 40100 14795 40103
rect 15746 40100 15752 40112
rect 14783 40072 15752 40100
rect 14783 40069 14795 40072
rect 14737 40063 14795 40069
rect 1394 39964 1400 39976
rect 1355 39936 1400 39964
rect 1394 39924 1400 39936
rect 1452 39924 1458 39976
rect 12437 39967 12495 39973
rect 12437 39933 12449 39967
rect 12483 39933 12495 39967
rect 12618 39964 12624 39976
rect 12579 39936 12624 39964
rect 12437 39927 12495 39933
rect 12452 39896 12480 39927
rect 12618 39924 12624 39936
rect 12676 39924 12682 39976
rect 12713 39967 12771 39973
rect 12713 39933 12725 39967
rect 12759 39964 12771 39967
rect 13262 39964 13268 39976
rect 12759 39936 13268 39964
rect 12759 39933 12771 39936
rect 12713 39927 12771 39933
rect 13262 39924 13268 39936
rect 13320 39924 13326 39976
rect 15337 39973 15365 40072
rect 15746 40060 15752 40072
rect 15804 40100 15810 40112
rect 15804 40072 15884 40100
rect 15804 40060 15810 40072
rect 15856 40041 15884 40072
rect 15841 40035 15899 40041
rect 15841 40001 15853 40035
rect 15887 40001 15899 40035
rect 15841 39995 15899 40001
rect 34054 39992 34060 40044
rect 34112 40032 34118 40044
rect 34977 40035 35035 40041
rect 34977 40032 34989 40035
rect 34112 40004 34989 40032
rect 34112 39992 34118 40004
rect 34977 40001 34989 40004
rect 35023 40001 35035 40035
rect 34977 39995 35035 40001
rect 13357 39967 13415 39973
rect 13357 39933 13369 39967
rect 13403 39964 13415 39967
rect 15335 39967 15393 39973
rect 13403 39936 13584 39964
rect 13403 39933 13415 39936
rect 13357 39927 13415 39933
rect 13446 39896 13452 39908
rect 12452 39868 13452 39896
rect 13446 39856 13452 39868
rect 13504 39856 13510 39908
rect 12250 39828 12256 39840
rect 12211 39800 12256 39828
rect 12250 39788 12256 39800
rect 12308 39788 12314 39840
rect 13556 39828 13584 39936
rect 15335 39933 15347 39967
rect 15381 39933 15393 39967
rect 15749 39967 15807 39973
rect 15749 39964 15761 39967
rect 15335 39927 15393 39933
rect 15488 39936 15761 39964
rect 13624 39899 13682 39905
rect 13624 39865 13636 39899
rect 13670 39896 13682 39899
rect 13670 39868 15240 39896
rect 13670 39865 13682 39868
rect 13624 39859 13682 39865
rect 13722 39828 13728 39840
rect 13556 39800 13728 39828
rect 13722 39788 13728 39800
rect 13780 39828 13786 39840
rect 13998 39828 14004 39840
rect 13780 39800 14004 39828
rect 13780 39788 13786 39800
rect 13998 39788 14004 39800
rect 14056 39788 14062 39840
rect 15212 39837 15240 39868
rect 15488 39840 15516 39936
rect 15749 39933 15761 39936
rect 15795 39933 15807 39967
rect 15749 39927 15807 39933
rect 16758 39924 16764 39976
rect 16816 39964 16822 39976
rect 17678 39964 17684 39976
rect 16816 39936 17684 39964
rect 16816 39924 16822 39936
rect 17678 39924 17684 39936
rect 17736 39964 17742 39976
rect 18598 39973 18604 39976
rect 18325 39967 18383 39973
rect 18325 39964 18337 39967
rect 17736 39936 18337 39964
rect 17736 39924 17742 39936
rect 18325 39933 18337 39936
rect 18371 39933 18383 39967
rect 18592 39964 18604 39973
rect 18559 39936 18604 39964
rect 18325 39927 18383 39933
rect 18592 39927 18604 39936
rect 18598 39924 18604 39927
rect 18656 39924 18662 39976
rect 20438 39973 20444 39976
rect 20165 39967 20223 39973
rect 20165 39933 20177 39967
rect 20211 39933 20223 39967
rect 20432 39964 20444 39973
rect 20399 39936 20444 39964
rect 20165 39927 20223 39933
rect 20432 39927 20444 39936
rect 20180 39896 20208 39927
rect 20438 39924 20444 39927
rect 20496 39924 20502 39976
rect 25958 39964 25964 39976
rect 25919 39936 25964 39964
rect 25958 39924 25964 39936
rect 26016 39924 26022 39976
rect 27801 39967 27859 39973
rect 27801 39933 27813 39967
rect 27847 39964 27859 39967
rect 29641 39967 29699 39973
rect 27847 39936 29592 39964
rect 27847 39933 27859 39936
rect 27801 39927 27859 39933
rect 20714 39896 20720 39908
rect 20180 39868 20720 39896
rect 20714 39856 20720 39868
rect 20772 39856 20778 39908
rect 27706 39856 27712 39908
rect 27764 39896 27770 39908
rect 28046 39899 28104 39905
rect 28046 39896 28058 39899
rect 27764 39868 28058 39896
rect 27764 39856 27770 39868
rect 28046 39865 28058 39868
rect 28092 39865 28104 39899
rect 29564 39896 29592 39936
rect 29641 39933 29653 39967
rect 29687 39964 29699 39967
rect 29822 39964 29828 39976
rect 29687 39936 29828 39964
rect 29687 39933 29699 39936
rect 29641 39927 29699 39933
rect 29822 39924 29828 39936
rect 29880 39924 29886 39976
rect 30469 39967 30527 39973
rect 30469 39933 30481 39967
rect 30515 39933 30527 39967
rect 30469 39927 30527 39933
rect 30736 39967 30794 39973
rect 30736 39933 30748 39967
rect 30782 39964 30794 39967
rect 31294 39964 31300 39976
rect 30782 39936 31300 39964
rect 30782 39933 30794 39936
rect 30736 39927 30794 39933
rect 30484 39896 30512 39927
rect 31294 39924 31300 39936
rect 31352 39924 31358 39976
rect 33045 39967 33103 39973
rect 33045 39933 33057 39967
rect 33091 39933 33103 39967
rect 33045 39927 33103 39933
rect 30926 39896 30932 39908
rect 29564 39868 30932 39896
rect 28046 39859 28104 39865
rect 30926 39856 30932 39868
rect 30984 39856 30990 39908
rect 33060 39896 33088 39927
rect 33134 39924 33140 39976
rect 33192 39964 33198 39976
rect 33301 39967 33359 39973
rect 33301 39964 33313 39967
rect 33192 39936 33313 39964
rect 33192 39924 33198 39936
rect 33301 39933 33313 39936
rect 33347 39933 33359 39967
rect 34885 39967 34943 39973
rect 34885 39964 34897 39967
rect 33301 39927 33359 39933
rect 34440 39936 34897 39964
rect 33410 39896 33416 39908
rect 33060 39868 33416 39896
rect 33410 39856 33416 39868
rect 33468 39856 33474 39908
rect 15197 39831 15255 39837
rect 15197 39797 15209 39831
rect 15243 39797 15255 39831
rect 15197 39791 15255 39797
rect 15381 39831 15439 39837
rect 15381 39797 15393 39831
rect 15427 39828 15439 39831
rect 15470 39828 15476 39840
rect 15427 39800 15476 39828
rect 15427 39797 15439 39800
rect 15381 39791 15439 39797
rect 15470 39788 15476 39800
rect 15528 39788 15534 39840
rect 26050 39828 26056 39840
rect 26011 39800 26056 39828
rect 26050 39788 26056 39800
rect 26108 39788 26114 39840
rect 27890 39788 27896 39840
rect 27948 39828 27954 39840
rect 34440 39837 34468 39936
rect 34885 39933 34897 39936
rect 34931 39933 34943 39967
rect 34885 39927 34943 39933
rect 57977 39967 58035 39973
rect 57977 39933 57989 39967
rect 58023 39964 58035 39967
rect 58618 39964 58624 39976
rect 58023 39936 58624 39964
rect 58023 39933 58035 39936
rect 57977 39927 58035 39933
rect 58618 39924 58624 39936
rect 58676 39924 58682 39976
rect 58158 39896 58164 39908
rect 58119 39868 58164 39896
rect 58158 39856 58164 39868
rect 58216 39856 58222 39908
rect 29181 39831 29239 39837
rect 29181 39828 29193 39831
rect 27948 39800 29193 39828
rect 27948 39788 27954 39800
rect 29181 39797 29193 39800
rect 29227 39797 29239 39831
rect 29181 39791 29239 39797
rect 34425 39831 34483 39837
rect 34425 39797 34437 39831
rect 34471 39797 34483 39831
rect 34425 39791 34483 39797
rect 1104 39738 58880 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 58880 39738
rect 1104 39664 58880 39686
rect 12618 39584 12624 39636
rect 12676 39624 12682 39636
rect 12897 39627 12955 39633
rect 12897 39624 12909 39627
rect 12676 39596 12909 39624
rect 12676 39584 12682 39596
rect 12897 39593 12909 39596
rect 12943 39593 12955 39627
rect 13446 39624 13452 39636
rect 13407 39596 13452 39624
rect 12897 39587 12955 39593
rect 11784 39559 11842 39565
rect 11784 39525 11796 39559
rect 11830 39556 11842 39559
rect 12250 39556 12256 39568
rect 11830 39528 12256 39556
rect 11830 39525 11842 39528
rect 11784 39519 11842 39525
rect 12250 39516 12256 39528
rect 12308 39516 12314 39568
rect 11517 39491 11575 39497
rect 11517 39457 11529 39491
rect 11563 39488 11575 39491
rect 12912 39488 12940 39587
rect 13446 39584 13452 39596
rect 13504 39584 13510 39636
rect 16758 39584 16764 39636
rect 16816 39624 16822 39636
rect 17313 39627 17371 39633
rect 17313 39624 17325 39627
rect 16816 39596 17325 39624
rect 16816 39584 16822 39596
rect 17313 39593 17325 39596
rect 17359 39593 17371 39627
rect 20898 39624 20904 39636
rect 20859 39596 20904 39624
rect 17313 39587 17371 39593
rect 20898 39584 20904 39596
rect 20956 39584 20962 39636
rect 25958 39584 25964 39636
rect 26016 39624 26022 39636
rect 26881 39627 26939 39633
rect 26881 39624 26893 39627
rect 26016 39596 26893 39624
rect 26016 39584 26022 39596
rect 26881 39593 26893 39596
rect 26927 39593 26939 39627
rect 28166 39624 28172 39636
rect 28127 39596 28172 39624
rect 26881 39587 26939 39593
rect 28166 39584 28172 39596
rect 28224 39584 28230 39636
rect 31297 39627 31355 39633
rect 31297 39593 31309 39627
rect 31343 39624 31355 39627
rect 31570 39624 31576 39636
rect 31343 39596 31576 39624
rect 31343 39593 31355 39596
rect 31297 39587 31355 39593
rect 31570 39584 31576 39596
rect 31628 39584 31634 39636
rect 33042 39624 33048 39636
rect 33003 39596 33048 39624
rect 33042 39584 33048 39596
rect 33100 39584 33106 39636
rect 15378 39516 15384 39568
rect 15436 39565 15442 39568
rect 15436 39559 15500 39565
rect 15436 39525 15454 39559
rect 15488 39525 15500 39559
rect 15436 39519 15500 39525
rect 25768 39559 25826 39565
rect 25768 39525 25780 39559
rect 25814 39556 25826 39559
rect 26050 39556 26056 39568
rect 25814 39528 26056 39556
rect 25814 39525 25826 39528
rect 25768 39519 25826 39525
rect 15436 39516 15442 39519
rect 26050 39516 26056 39528
rect 26108 39516 26114 39568
rect 33870 39556 33876 39568
rect 32600 39528 32996 39556
rect 13357 39491 13415 39497
rect 13357 39488 13369 39491
rect 11563 39460 12848 39488
rect 12912 39460 13369 39488
rect 11563 39457 11575 39460
rect 11517 39451 11575 39457
rect 12820 39352 12848 39460
rect 13357 39457 13369 39460
rect 13403 39457 13415 39491
rect 13357 39451 13415 39457
rect 13541 39491 13599 39497
rect 13541 39457 13553 39491
rect 13587 39457 13599 39491
rect 13541 39451 13599 39457
rect 17497 39491 17555 39497
rect 17497 39457 17509 39491
rect 17543 39488 17555 39491
rect 18046 39488 18052 39500
rect 17543 39460 18052 39488
rect 17543 39457 17555 39460
rect 17497 39451 17555 39457
rect 13262 39380 13268 39432
rect 13320 39420 13326 39432
rect 13556 39420 13584 39451
rect 18046 39448 18052 39460
rect 18104 39448 18110 39500
rect 20070 39448 20076 39500
rect 20128 39488 20134 39500
rect 20165 39491 20223 39497
rect 20165 39488 20177 39491
rect 20128 39460 20177 39488
rect 20128 39448 20134 39460
rect 20165 39457 20177 39460
rect 20211 39457 20223 39491
rect 20165 39451 20223 39457
rect 20257 39491 20315 39497
rect 20257 39457 20269 39491
rect 20303 39488 20315 39491
rect 20806 39488 20812 39500
rect 20303 39460 20812 39488
rect 20303 39457 20315 39460
rect 20257 39451 20315 39457
rect 20806 39448 20812 39460
rect 20864 39448 20870 39500
rect 20993 39491 21051 39497
rect 20993 39457 21005 39491
rect 21039 39488 21051 39491
rect 21082 39488 21088 39500
rect 21039 39460 21088 39488
rect 21039 39457 21051 39460
rect 20993 39451 21051 39457
rect 21082 39448 21088 39460
rect 21140 39448 21146 39500
rect 27338 39488 27344 39500
rect 27299 39460 27344 39488
rect 27338 39448 27344 39460
rect 27396 39448 27402 39500
rect 27982 39448 27988 39500
rect 28040 39488 28046 39500
rect 28077 39491 28135 39497
rect 28077 39488 28089 39491
rect 28040 39460 28089 39488
rect 28040 39448 28046 39460
rect 28077 39457 28089 39460
rect 28123 39457 28135 39491
rect 28077 39451 28135 39457
rect 31205 39491 31263 39497
rect 31205 39457 31217 39491
rect 31251 39488 31263 39491
rect 31754 39488 31760 39500
rect 31251 39460 31760 39488
rect 31251 39457 31263 39460
rect 31205 39451 31263 39457
rect 31754 39448 31760 39460
rect 31812 39448 31818 39500
rect 31849 39491 31907 39497
rect 31849 39457 31861 39491
rect 31895 39488 31907 39491
rect 32122 39488 32128 39500
rect 31895 39460 32128 39488
rect 31895 39457 31907 39460
rect 31849 39451 31907 39457
rect 32122 39448 32128 39460
rect 32180 39448 32186 39500
rect 32600 39497 32628 39528
rect 32585 39491 32643 39497
rect 32585 39457 32597 39491
rect 32631 39457 32643 39491
rect 32585 39451 32643 39457
rect 32769 39491 32827 39497
rect 32769 39457 32781 39491
rect 32815 39457 32827 39491
rect 32769 39451 32827 39457
rect 13320 39392 13584 39420
rect 13320 39380 13326 39392
rect 13722 39380 13728 39432
rect 13780 39420 13786 39432
rect 15197 39423 15255 39429
rect 15197 39420 15209 39423
rect 13780 39392 15209 39420
rect 13780 39380 13786 39392
rect 15197 39389 15209 39392
rect 15243 39389 15255 39423
rect 25498 39420 25504 39432
rect 25459 39392 25504 39420
rect 15197 39383 15255 39389
rect 25498 39380 25504 39392
rect 25556 39380 25562 39432
rect 31941 39423 31999 39429
rect 31941 39389 31953 39423
rect 31987 39420 31999 39423
rect 32784 39420 32812 39451
rect 32858 39420 32864 39432
rect 31987 39392 32864 39420
rect 31987 39389 31999 39392
rect 31941 39383 31999 39389
rect 32858 39380 32864 39392
rect 32916 39380 32922 39432
rect 13740 39352 13768 39380
rect 12820 39324 13768 39352
rect 15562 39244 15568 39296
rect 15620 39284 15626 39296
rect 16577 39287 16635 39293
rect 16577 39284 16589 39287
rect 15620 39256 16589 39284
rect 15620 39244 15626 39256
rect 16577 39253 16589 39256
rect 16623 39253 16635 39287
rect 16577 39247 16635 39253
rect 27433 39287 27491 39293
rect 27433 39253 27445 39287
rect 27479 39284 27491 39287
rect 28534 39284 28540 39296
rect 27479 39256 28540 39284
rect 27479 39253 27491 39256
rect 27433 39247 27491 39253
rect 28534 39244 28540 39256
rect 28592 39244 28598 39296
rect 32968 39284 32996 39528
rect 33060 39528 33876 39556
rect 33060 39497 33088 39528
rect 33870 39516 33876 39528
rect 33928 39516 33934 39568
rect 33045 39491 33103 39497
rect 33045 39457 33057 39491
rect 33091 39457 33103 39491
rect 33045 39451 33103 39457
rect 33137 39491 33195 39497
rect 33137 39457 33149 39491
rect 33183 39457 33195 39491
rect 57974 39488 57980 39500
rect 57935 39460 57980 39488
rect 33137 39451 33195 39457
rect 33152 39420 33180 39451
rect 57974 39448 57980 39460
rect 58032 39448 58038 39500
rect 33060 39392 33180 39420
rect 33060 39364 33088 39392
rect 33042 39312 33048 39364
rect 33100 39312 33106 39364
rect 33226 39284 33232 39296
rect 32968 39256 33232 39284
rect 33226 39244 33232 39256
rect 33284 39244 33290 39296
rect 1104 39194 58880 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 58880 39194
rect 1104 39120 58880 39142
rect 13449 39083 13507 39089
rect 13449 39049 13461 39083
rect 13495 39080 13507 39083
rect 14921 39083 14979 39089
rect 14921 39080 14933 39083
rect 13495 39052 14933 39080
rect 13495 39049 13507 39052
rect 13449 39043 13507 39049
rect 1394 38876 1400 38888
rect 1355 38848 1400 38876
rect 1394 38836 1400 38848
rect 1452 38836 1458 38888
rect 12437 38879 12495 38885
rect 12437 38845 12449 38879
rect 12483 38876 12495 38879
rect 13262 38876 13268 38888
rect 12483 38848 13268 38876
rect 12483 38845 12495 38848
rect 12437 38839 12495 38845
rect 13262 38836 13268 38848
rect 13320 38836 13326 38888
rect 13357 38879 13415 38885
rect 13357 38845 13369 38879
rect 13403 38876 13415 38879
rect 13446 38876 13452 38888
rect 13403 38848 13452 38876
rect 13403 38845 13415 38848
rect 13357 38839 13415 38845
rect 13446 38836 13452 38848
rect 13504 38836 13510 38888
rect 12526 38740 12532 38752
rect 12487 38712 12532 38740
rect 12526 38700 12532 38712
rect 12584 38700 12590 38752
rect 14660 38740 14688 39052
rect 14921 39049 14933 39052
rect 14967 39049 14979 39083
rect 14921 39043 14979 39049
rect 15194 39040 15200 39092
rect 15252 39080 15258 39092
rect 15565 39083 15623 39089
rect 15565 39080 15577 39083
rect 15252 39052 15577 39080
rect 15252 39040 15258 39052
rect 15565 39049 15577 39052
rect 15611 39049 15623 39083
rect 15565 39043 15623 39049
rect 19978 39040 19984 39092
rect 20036 39080 20042 39092
rect 20533 39083 20591 39089
rect 20533 39080 20545 39083
rect 20036 39052 20545 39080
rect 20036 39040 20042 39052
rect 20533 39049 20545 39052
rect 20579 39049 20591 39083
rect 20533 39043 20591 39049
rect 15105 39015 15163 39021
rect 15105 38981 15117 39015
rect 15151 39012 15163 39015
rect 15286 39012 15292 39024
rect 15151 38984 15292 39012
rect 15151 38981 15163 38984
rect 15105 38975 15163 38981
rect 15286 38972 15292 38984
rect 15344 38972 15350 39024
rect 25866 39012 25872 39024
rect 25779 38984 25872 39012
rect 25866 38972 25872 38984
rect 25924 39012 25930 39024
rect 26697 39015 26755 39021
rect 26697 39012 26709 39015
rect 25924 38984 26709 39012
rect 25924 38972 25930 38984
rect 26697 38981 26709 38984
rect 26743 38981 26755 39015
rect 26697 38975 26755 38981
rect 32033 39015 32091 39021
rect 32033 38981 32045 39015
rect 32079 39012 32091 39015
rect 33045 39015 33103 39021
rect 33045 39012 33057 39015
rect 32079 38984 33057 39012
rect 32079 38981 32091 38984
rect 32033 38975 32091 38981
rect 33045 38981 33057 38984
rect 33091 39012 33103 39015
rect 33686 39012 33692 39024
rect 33091 38984 33692 39012
rect 33091 38981 33103 38984
rect 33045 38975 33103 38981
rect 33686 38972 33692 38984
rect 33744 38972 33750 39024
rect 17678 38944 17684 38956
rect 14752 38916 15792 38944
rect 17639 38916 17684 38944
rect 14752 38817 14780 38916
rect 15764 38888 15792 38916
rect 17678 38904 17684 38916
rect 17736 38904 17742 38956
rect 25958 38904 25964 38956
rect 26016 38944 26022 38956
rect 26789 38947 26847 38953
rect 26789 38944 26801 38947
rect 26016 38916 26801 38944
rect 26016 38904 26022 38916
rect 26789 38913 26801 38916
rect 26835 38913 26847 38947
rect 32122 38944 32128 38956
rect 32083 38916 32128 38944
rect 26789 38907 26847 38913
rect 32122 38904 32128 38916
rect 32180 38904 32186 38956
rect 15562 38876 15568 38888
rect 15523 38848 15568 38876
rect 15562 38836 15568 38848
rect 15620 38836 15626 38888
rect 15746 38876 15752 38888
rect 15707 38848 15752 38876
rect 15746 38836 15752 38848
rect 15804 38836 15810 38888
rect 15841 38879 15899 38885
rect 15841 38845 15853 38879
rect 15887 38845 15899 38879
rect 15841 38839 15899 38845
rect 19705 38879 19763 38885
rect 19705 38845 19717 38879
rect 19751 38845 19763 38879
rect 19886 38876 19892 38888
rect 19847 38848 19892 38876
rect 19705 38839 19763 38845
rect 14737 38811 14795 38817
rect 14737 38777 14749 38811
rect 14783 38777 14795 38811
rect 14737 38771 14795 38777
rect 14953 38811 15011 38817
rect 14953 38777 14965 38811
rect 14999 38808 15011 38811
rect 15580 38808 15608 38836
rect 14999 38780 15608 38808
rect 14999 38777 15011 38780
rect 14953 38771 15011 38777
rect 15470 38740 15476 38752
rect 14660 38712 15476 38740
rect 15470 38700 15476 38712
rect 15528 38740 15534 38752
rect 15856 38740 15884 38839
rect 17948 38811 18006 38817
rect 17948 38777 17960 38811
rect 17994 38808 18006 38811
rect 18966 38808 18972 38820
rect 17994 38780 18972 38808
rect 17994 38777 18006 38780
rect 17948 38771 18006 38777
rect 18966 38768 18972 38780
rect 19024 38768 19030 38820
rect 19720 38808 19748 38839
rect 19886 38836 19892 38848
rect 19944 38836 19950 38888
rect 19978 38836 19984 38888
rect 20036 38876 20042 38888
rect 20438 38876 20444 38888
rect 20036 38848 20081 38876
rect 20399 38848 20444 38876
rect 20036 38836 20042 38848
rect 20438 38836 20444 38848
rect 20496 38836 20502 38888
rect 20714 38836 20720 38888
rect 20772 38876 20778 38888
rect 24489 38879 24547 38885
rect 24489 38876 24501 38879
rect 20772 38848 24501 38876
rect 20772 38836 20778 38848
rect 24489 38845 24501 38848
rect 24535 38845 24547 38879
rect 26510 38876 26516 38888
rect 26423 38848 26516 38876
rect 24489 38839 24547 38845
rect 26510 38836 26516 38848
rect 26568 38876 26574 38888
rect 27338 38876 27344 38888
rect 26568 38848 27344 38876
rect 26568 38836 26574 38848
rect 27338 38836 27344 38848
rect 27396 38836 27402 38888
rect 28353 38879 28411 38885
rect 28353 38845 28365 38879
rect 28399 38876 28411 38879
rect 30926 38876 30932 38888
rect 28399 38848 30932 38876
rect 28399 38845 28411 38848
rect 28353 38839 28411 38845
rect 30926 38836 30932 38848
rect 30984 38836 30990 38888
rect 31754 38836 31760 38888
rect 31812 38876 31818 38888
rect 31849 38879 31907 38885
rect 31849 38876 31861 38879
rect 31812 38848 31861 38876
rect 31812 38836 31818 38848
rect 31849 38845 31861 38848
rect 31895 38876 31907 38879
rect 32398 38876 32404 38888
rect 31895 38848 32404 38876
rect 31895 38845 31907 38848
rect 31849 38839 31907 38845
rect 32398 38836 32404 38848
rect 32456 38836 32462 38888
rect 33042 38876 33048 38888
rect 33003 38848 33048 38876
rect 33042 38836 33048 38848
rect 33100 38836 33106 38888
rect 33226 38876 33232 38888
rect 33187 38848 33232 38876
rect 33226 38836 33232 38848
rect 33284 38836 33290 38888
rect 33410 38836 33416 38888
rect 33468 38876 33474 38888
rect 33689 38879 33747 38885
rect 33689 38876 33701 38879
rect 33468 38848 33701 38876
rect 33468 38836 33474 38848
rect 33689 38845 33701 38848
rect 33735 38845 33747 38879
rect 33689 38839 33747 38845
rect 20456 38808 20484 38836
rect 19720 38780 20484 38808
rect 24756 38811 24814 38817
rect 24756 38777 24768 38811
rect 24802 38808 24814 38811
rect 26329 38811 26387 38817
rect 26329 38808 26341 38811
rect 24802 38780 26341 38808
rect 24802 38777 24814 38780
rect 24756 38771 24814 38777
rect 26329 38777 26341 38780
rect 26375 38777 26387 38811
rect 26329 38771 26387 38777
rect 28620 38811 28678 38817
rect 28620 38777 28632 38811
rect 28666 38808 28678 38811
rect 28810 38808 28816 38820
rect 28666 38780 28816 38808
rect 28666 38777 28678 38780
rect 28620 38771 28678 38777
rect 28810 38768 28816 38780
rect 28868 38768 28874 38820
rect 33962 38817 33968 38820
rect 33956 38771 33968 38817
rect 34020 38808 34026 38820
rect 57974 38808 57980 38820
rect 34020 38780 34056 38808
rect 57935 38780 57980 38808
rect 33962 38768 33968 38771
rect 34020 38768 34026 38780
rect 57974 38768 57980 38780
rect 58032 38768 58038 38820
rect 58158 38808 58164 38820
rect 58119 38780 58164 38808
rect 58158 38768 58164 38780
rect 58216 38768 58222 38820
rect 15528 38712 15884 38740
rect 15528 38700 15534 38712
rect 18230 38700 18236 38752
rect 18288 38740 18294 38752
rect 19061 38743 19119 38749
rect 19061 38740 19073 38743
rect 18288 38712 19073 38740
rect 18288 38700 18294 38712
rect 19061 38709 19073 38712
rect 19107 38709 19119 38743
rect 19061 38703 19119 38709
rect 19521 38743 19579 38749
rect 19521 38709 19533 38743
rect 19567 38740 19579 38743
rect 20162 38740 20168 38752
rect 19567 38712 20168 38740
rect 19567 38709 19579 38712
rect 19521 38703 19579 38709
rect 20162 38700 20168 38712
rect 20220 38700 20226 38752
rect 29178 38700 29184 38752
rect 29236 38740 29242 38752
rect 29733 38743 29791 38749
rect 29733 38740 29745 38743
rect 29236 38712 29745 38740
rect 29236 38700 29242 38712
rect 29733 38709 29745 38712
rect 29779 38709 29791 38743
rect 31662 38740 31668 38752
rect 31623 38712 31668 38740
rect 29733 38703 29791 38709
rect 31662 38700 31668 38712
rect 31720 38700 31726 38752
rect 35069 38743 35127 38749
rect 35069 38709 35081 38743
rect 35115 38740 35127 38743
rect 35250 38740 35256 38752
rect 35115 38712 35256 38740
rect 35115 38709 35127 38712
rect 35069 38703 35127 38709
rect 35250 38700 35256 38712
rect 35308 38700 35314 38752
rect 1104 38650 58880 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 58880 38650
rect 1104 38576 58880 38598
rect 13262 38536 13268 38548
rect 13223 38508 13268 38536
rect 13262 38496 13268 38508
rect 13320 38496 13326 38548
rect 17313 38539 17371 38545
rect 17313 38505 17325 38539
rect 17359 38536 17371 38539
rect 18966 38536 18972 38548
rect 17359 38508 18092 38536
rect 18927 38508 18972 38536
rect 17359 38505 17371 38508
rect 17313 38499 17371 38505
rect 12152 38471 12210 38477
rect 12152 38437 12164 38471
rect 12198 38468 12210 38471
rect 12526 38468 12532 38480
rect 12198 38440 12532 38468
rect 12198 38437 12210 38440
rect 12152 38431 12210 38437
rect 12526 38428 12532 38440
rect 12584 38428 12590 38480
rect 16758 38468 16764 38480
rect 15948 38440 16764 38468
rect 1394 38400 1400 38412
rect 1355 38372 1400 38400
rect 1394 38360 1400 38372
rect 1452 38360 1458 38412
rect 11885 38403 11943 38409
rect 11885 38369 11897 38403
rect 11931 38400 11943 38403
rect 13722 38400 13728 38412
rect 11931 38372 13728 38400
rect 11931 38369 11943 38372
rect 11885 38363 11943 38369
rect 13722 38360 13728 38372
rect 13780 38360 13786 38412
rect 14921 38403 14979 38409
rect 14921 38369 14933 38403
rect 14967 38400 14979 38403
rect 15654 38400 15660 38412
rect 14967 38372 15660 38400
rect 14967 38369 14979 38372
rect 14921 38363 14979 38369
rect 15654 38360 15660 38372
rect 15712 38360 15718 38412
rect 15948 38409 15976 38440
rect 16758 38428 16764 38440
rect 16816 38428 16822 38480
rect 17954 38428 17960 38480
rect 18012 38468 18018 38480
rect 18064 38477 18092 38508
rect 18966 38496 18972 38508
rect 19024 38496 19030 38548
rect 19978 38496 19984 38548
rect 20036 38536 20042 38548
rect 21361 38539 21419 38545
rect 21361 38536 21373 38539
rect 20036 38508 21373 38536
rect 20036 38496 20042 38508
rect 21361 38505 21373 38508
rect 21407 38505 21419 38539
rect 21361 38499 21419 38505
rect 26053 38539 26111 38545
rect 26053 38505 26065 38539
rect 26099 38536 26111 38539
rect 26510 38536 26516 38548
rect 26099 38508 26516 38536
rect 26099 38505 26111 38508
rect 26053 38499 26111 38505
rect 26510 38496 26516 38508
rect 26568 38496 26574 38548
rect 27893 38539 27951 38545
rect 27893 38505 27905 38539
rect 27939 38536 27951 38539
rect 29365 38539 29423 38545
rect 29365 38536 29377 38539
rect 27939 38508 29377 38536
rect 27939 38505 27951 38508
rect 27893 38499 27951 38505
rect 18049 38471 18107 38477
rect 18049 38468 18061 38471
rect 18012 38440 18061 38468
rect 18012 38428 18018 38440
rect 18049 38437 18061 38440
rect 18095 38437 18107 38471
rect 18049 38431 18107 38437
rect 18265 38471 18323 38477
rect 18265 38437 18277 38471
rect 18311 38468 18323 38471
rect 18690 38468 18696 38480
rect 18311 38440 18696 38468
rect 18311 38437 18323 38440
rect 18265 38431 18323 38437
rect 18690 38428 18696 38440
rect 18748 38428 18754 38480
rect 20162 38428 20168 38480
rect 20220 38477 20226 38480
rect 28368 38477 28396 38508
rect 29365 38505 29377 38508
rect 29411 38505 29423 38539
rect 29365 38499 29423 38505
rect 32122 38496 32128 38548
rect 32180 38536 32186 38548
rect 32309 38539 32367 38545
rect 32309 38536 32321 38539
rect 32180 38508 32321 38536
rect 32180 38496 32186 38508
rect 32309 38505 32321 38508
rect 32355 38505 32367 38539
rect 32309 38499 32367 38505
rect 32398 38496 32404 38548
rect 32456 38536 32462 38548
rect 33229 38539 33287 38545
rect 33229 38536 33241 38539
rect 32456 38508 33241 38536
rect 32456 38496 32462 38508
rect 33229 38505 33241 38508
rect 33275 38505 33287 38539
rect 33229 38499 33287 38505
rect 57974 38496 57980 38548
rect 58032 38536 58038 38548
rect 58161 38539 58219 38545
rect 58161 38536 58173 38539
rect 58032 38508 58173 38536
rect 58032 38496 58038 38508
rect 58161 38505 58173 38508
rect 58207 38505 58219 38539
rect 58161 38499 58219 38505
rect 20220 38471 20284 38477
rect 20220 38437 20238 38471
rect 20272 38437 20284 38471
rect 20220 38431 20284 38437
rect 28353 38471 28411 38477
rect 28353 38437 28365 38471
rect 28399 38468 28411 38471
rect 28442 38468 28448 38480
rect 28399 38440 28448 38468
rect 28399 38437 28411 38440
rect 28353 38431 28411 38437
rect 20220 38428 20226 38431
rect 28442 38428 28448 38440
rect 28500 38428 28506 38480
rect 28569 38471 28627 38477
rect 28569 38437 28581 38471
rect 28615 38468 28627 38471
rect 29178 38468 29184 38480
rect 28615 38440 29184 38468
rect 28615 38437 28627 38440
rect 28569 38431 28627 38437
rect 29178 38428 29184 38440
rect 29236 38428 29242 38480
rect 31196 38471 31254 38477
rect 31196 38437 31208 38471
rect 31242 38468 31254 38471
rect 31662 38468 31668 38480
rect 31242 38440 31668 38468
rect 31242 38437 31254 38440
rect 31196 38431 31254 38437
rect 31662 38428 31668 38440
rect 31720 38428 31726 38480
rect 33686 38428 33692 38480
rect 33744 38468 33750 38480
rect 33965 38471 34023 38477
rect 33965 38468 33977 38471
rect 33744 38440 33977 38468
rect 33744 38428 33750 38440
rect 33965 38437 33977 38440
rect 34011 38437 34023 38471
rect 33965 38431 34023 38437
rect 15933 38403 15991 38409
rect 15933 38369 15945 38403
rect 15979 38369 15991 38403
rect 15933 38363 15991 38369
rect 16200 38403 16258 38409
rect 16200 38369 16212 38403
rect 16246 38400 16258 38403
rect 17310 38400 17316 38412
rect 16246 38372 17316 38400
rect 16246 38369 16258 38372
rect 16200 38363 16258 38369
rect 17310 38360 17316 38372
rect 17368 38360 17374 38412
rect 18874 38400 18880 38412
rect 18835 38372 18880 38400
rect 18874 38360 18880 38372
rect 18932 38360 18938 38412
rect 19061 38403 19119 38409
rect 19061 38369 19073 38403
rect 19107 38400 19119 38403
rect 19886 38400 19892 38412
rect 19107 38372 19892 38400
rect 19107 38369 19119 38372
rect 19061 38363 19119 38369
rect 15102 38292 15108 38344
rect 15160 38332 15166 38344
rect 15197 38335 15255 38341
rect 15197 38332 15209 38335
rect 15160 38304 15209 38332
rect 15160 38292 15166 38304
rect 15197 38301 15209 38304
rect 15243 38301 15255 38335
rect 15197 38295 15255 38301
rect 18417 38267 18475 38273
rect 18417 38233 18429 38267
rect 18463 38264 18475 38267
rect 19076 38264 19104 38363
rect 19886 38360 19892 38372
rect 19944 38360 19950 38412
rect 19981 38403 20039 38409
rect 19981 38369 19993 38403
rect 20027 38400 20039 38403
rect 20714 38400 20720 38412
rect 20027 38372 20720 38400
rect 20027 38369 20039 38372
rect 19981 38363 20039 38369
rect 20714 38360 20720 38372
rect 20772 38360 20778 38412
rect 25866 38400 25872 38412
rect 25827 38372 25872 38400
rect 25866 38360 25872 38372
rect 25924 38360 25930 38412
rect 25958 38360 25964 38412
rect 26016 38400 26022 38412
rect 26053 38403 26111 38409
rect 26053 38400 26065 38403
rect 26016 38372 26065 38400
rect 26016 38360 26022 38372
rect 26053 38369 26065 38372
rect 26099 38369 26111 38403
rect 26053 38363 26111 38369
rect 26780 38403 26838 38409
rect 26780 38369 26792 38403
rect 26826 38400 26838 38403
rect 27798 38400 27804 38412
rect 26826 38372 27804 38400
rect 26826 38369 26838 38372
rect 26780 38363 26838 38369
rect 27798 38360 27804 38372
rect 27856 38360 27862 38412
rect 29457 38403 29515 38409
rect 29457 38400 29469 38403
rect 28552 38372 29469 38400
rect 28552 38344 28580 38372
rect 29457 38369 29469 38372
rect 29503 38369 29515 38403
rect 30926 38400 30932 38412
rect 30887 38372 30932 38400
rect 29457 38363 29515 38369
rect 30926 38360 30932 38372
rect 30984 38360 30990 38412
rect 32769 38403 32827 38409
rect 32769 38369 32781 38403
rect 32815 38369 32827 38403
rect 32769 38363 32827 38369
rect 25498 38292 25504 38344
rect 25556 38332 25562 38344
rect 26513 38335 26571 38341
rect 26513 38332 26525 38335
rect 25556 38304 26525 38332
rect 25556 38292 25562 38304
rect 26513 38301 26525 38304
rect 26559 38301 26571 38335
rect 26513 38295 26571 38301
rect 28534 38292 28540 38344
rect 28592 38292 28598 38344
rect 32784 38332 32812 38363
rect 32858 38360 32864 38412
rect 32916 38400 32922 38412
rect 33045 38403 33103 38409
rect 32916 38372 32961 38400
rect 32916 38360 32922 38372
rect 33045 38369 33057 38403
rect 33091 38400 33103 38403
rect 33226 38400 33232 38412
rect 33091 38372 33232 38400
rect 33091 38369 33103 38372
rect 33045 38363 33103 38369
rect 33226 38360 33232 38372
rect 33284 38400 33290 38412
rect 34146 38400 34152 38412
rect 33284 38372 34152 38400
rect 33284 38360 33290 38372
rect 34146 38360 34152 38372
rect 34204 38360 34210 38412
rect 34241 38403 34299 38409
rect 34241 38369 34253 38403
rect 34287 38369 34299 38403
rect 34241 38363 34299 38369
rect 34256 38332 34284 38363
rect 32784 38304 34284 38332
rect 57057 38335 57115 38341
rect 33060 38276 33088 38304
rect 57057 38301 57069 38335
rect 57103 38332 57115 38335
rect 57517 38335 57575 38341
rect 57517 38332 57529 38335
rect 57103 38304 57529 38332
rect 57103 38301 57115 38304
rect 57057 38295 57115 38301
rect 57517 38301 57529 38304
rect 57563 38301 57575 38335
rect 57698 38332 57704 38344
rect 57659 38304 57704 38332
rect 57517 38295 57575 38301
rect 57698 38292 57704 38304
rect 57756 38292 57762 38344
rect 18463 38236 19104 38264
rect 18463 38233 18475 38236
rect 18417 38227 18475 38233
rect 33042 38224 33048 38276
rect 33100 38224 33106 38276
rect 33962 38264 33968 38276
rect 33923 38236 33968 38264
rect 33962 38224 33968 38236
rect 34020 38224 34026 38276
rect 14734 38196 14740 38208
rect 14695 38168 14740 38196
rect 14734 38156 14740 38168
rect 14792 38156 14798 38208
rect 15105 38199 15163 38205
rect 15105 38165 15117 38199
rect 15151 38196 15163 38199
rect 15286 38196 15292 38208
rect 15151 38168 15292 38196
rect 15151 38165 15163 38168
rect 15105 38159 15163 38165
rect 15286 38156 15292 38168
rect 15344 38156 15350 38208
rect 18230 38196 18236 38208
rect 18191 38168 18236 38196
rect 18230 38156 18236 38168
rect 18288 38156 18294 38208
rect 28534 38196 28540 38208
rect 28495 38168 28540 38196
rect 28534 38156 28540 38168
rect 28592 38156 28598 38208
rect 28718 38196 28724 38208
rect 28679 38168 28724 38196
rect 28718 38156 28724 38168
rect 28776 38156 28782 38208
rect 28902 38156 28908 38208
rect 28960 38196 28966 38208
rect 29181 38199 29239 38205
rect 29181 38196 29193 38199
rect 28960 38168 29193 38196
rect 28960 38156 28966 38168
rect 29181 38165 29193 38168
rect 29227 38165 29239 38199
rect 29181 38159 29239 38165
rect 1104 38106 58880 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 58880 38106
rect 1104 38032 58880 38054
rect 15102 37992 15108 38004
rect 15063 37964 15108 37992
rect 15102 37952 15108 37964
rect 15160 37952 15166 38004
rect 15654 37992 15660 38004
rect 15615 37964 15660 37992
rect 15654 37952 15660 37964
rect 15712 37952 15718 38004
rect 17310 37992 17316 38004
rect 17271 37964 17316 37992
rect 17310 37952 17316 37964
rect 17368 37952 17374 38004
rect 18417 37995 18475 38001
rect 18417 37961 18429 37995
rect 18463 37992 18475 37995
rect 18874 37992 18880 38004
rect 18463 37964 18880 37992
rect 18463 37961 18475 37964
rect 18417 37955 18475 37961
rect 18874 37952 18880 37964
rect 18932 37952 18938 38004
rect 27798 37992 27804 38004
rect 27759 37964 27804 37992
rect 27798 37952 27804 37964
rect 27856 37952 27862 38004
rect 28353 37995 28411 38001
rect 28353 37961 28365 37995
rect 28399 37992 28411 37995
rect 28534 37992 28540 38004
rect 28399 37964 28540 37992
rect 28399 37961 28411 37964
rect 28353 37955 28411 37961
rect 28534 37952 28540 37964
rect 28592 37952 28598 38004
rect 28810 37952 28816 38004
rect 28868 37992 28874 38004
rect 28905 37995 28963 38001
rect 28905 37992 28917 37995
rect 28868 37964 28917 37992
rect 28868 37952 28874 37964
rect 28905 37961 28917 37964
rect 28951 37961 28963 37995
rect 28905 37955 28963 37961
rect 34146 37952 34152 38004
rect 34204 37992 34210 38004
rect 35161 37995 35219 38001
rect 35161 37992 35173 37995
rect 34204 37964 35173 37992
rect 34204 37952 34210 37964
rect 35161 37961 35173 37964
rect 35207 37961 35219 37995
rect 35161 37955 35219 37961
rect 57241 37995 57299 38001
rect 57241 37961 57253 37995
rect 57287 37992 57299 37995
rect 57698 37992 57704 38004
rect 57287 37964 57704 37992
rect 57287 37961 57299 37964
rect 57241 37955 57299 37961
rect 57698 37952 57704 37964
rect 57756 37952 57762 38004
rect 15120 37856 15148 37952
rect 17865 37927 17923 37933
rect 17865 37893 17877 37927
rect 17911 37924 17923 37927
rect 58158 37924 58164 37936
rect 17911 37896 18736 37924
rect 58119 37896 58164 37924
rect 17911 37893 17923 37896
rect 17865 37887 17923 37893
rect 17954 37856 17960 37868
rect 15120 37828 15792 37856
rect 13722 37788 13728 37800
rect 13683 37760 13728 37788
rect 13722 37748 13728 37760
rect 13780 37748 13786 37800
rect 13992 37791 14050 37797
rect 13992 37757 14004 37791
rect 14038 37788 14050 37791
rect 14734 37788 14740 37800
rect 14038 37760 14740 37788
rect 14038 37757 14050 37760
rect 13992 37751 14050 37757
rect 14734 37748 14740 37760
rect 14792 37748 14798 37800
rect 15286 37748 15292 37800
rect 15344 37788 15350 37800
rect 15764 37797 15792 37828
rect 17788 37828 17960 37856
rect 15565 37791 15623 37797
rect 15565 37788 15577 37791
rect 15344 37760 15577 37788
rect 15344 37748 15350 37760
rect 15565 37757 15577 37760
rect 15611 37757 15623 37791
rect 15565 37751 15623 37757
rect 15749 37791 15807 37797
rect 15749 37757 15761 37791
rect 15795 37757 15807 37791
rect 16390 37788 16396 37800
rect 16351 37760 16396 37788
rect 15749 37751 15807 37757
rect 16390 37748 16396 37760
rect 16448 37748 16454 37800
rect 17494 37791 17552 37797
rect 17494 37757 17506 37791
rect 17540 37788 17552 37791
rect 17788 37788 17816 37828
rect 17954 37816 17960 37828
rect 18012 37856 18018 37868
rect 18012 37828 18644 37856
rect 18012 37816 18018 37828
rect 17540 37760 17816 37788
rect 17540 37757 17552 37760
rect 17494 37751 17552 37757
rect 18230 37748 18236 37800
rect 18288 37788 18294 37800
rect 18616 37797 18644 37828
rect 18708 37800 18736 37896
rect 58158 37884 58164 37896
rect 58216 37884 58222 37936
rect 20990 37816 20996 37868
rect 21048 37856 21054 37868
rect 25314 37856 25320 37868
rect 21048 37828 25320 37856
rect 21048 37816 21054 37828
rect 25314 37816 25320 37828
rect 25372 37816 25378 37868
rect 28442 37856 28448 37868
rect 28276 37828 28448 37856
rect 18417 37791 18475 37797
rect 18417 37788 18429 37791
rect 18288 37760 18429 37788
rect 18288 37748 18294 37760
rect 18417 37757 18429 37760
rect 18463 37757 18475 37791
rect 18417 37751 18475 37757
rect 18601 37791 18659 37797
rect 18601 37757 18613 37791
rect 18647 37757 18659 37791
rect 18601 37751 18659 37757
rect 18690 37748 18696 37800
rect 18748 37788 18754 37800
rect 27982 37791 28040 37797
rect 18748 37760 18793 37788
rect 18748 37748 18754 37760
rect 27982 37757 27994 37791
rect 28028 37788 28040 37791
rect 28276 37788 28304 37828
rect 28442 37816 28448 37828
rect 28500 37816 28506 37868
rect 28718 37816 28724 37868
rect 28776 37856 28782 37868
rect 28776 37828 29132 37856
rect 28776 37816 28782 37828
rect 28902 37788 28908 37800
rect 28028 37760 28304 37788
rect 28863 37760 28908 37788
rect 28028 37757 28040 37760
rect 27982 37751 28040 37757
rect 28902 37748 28908 37760
rect 28960 37748 28966 37800
rect 29104 37797 29132 37828
rect 29089 37791 29147 37797
rect 29089 37757 29101 37791
rect 29135 37757 29147 37791
rect 33318 37788 33324 37800
rect 33279 37760 33324 37788
rect 29089 37751 29147 37757
rect 33318 37748 33324 37760
rect 33376 37748 33382 37800
rect 34425 37791 34483 37797
rect 34425 37757 34437 37791
rect 34471 37788 34483 37791
rect 34790 37788 34796 37800
rect 34471 37760 34796 37788
rect 34471 37757 34483 37760
rect 34425 37751 34483 37757
rect 34790 37748 34796 37760
rect 34848 37748 34854 37800
rect 35069 37791 35127 37797
rect 35069 37757 35081 37791
rect 35115 37788 35127 37791
rect 35250 37788 35256 37800
rect 35115 37760 35256 37788
rect 35115 37757 35127 37760
rect 35069 37751 35127 37757
rect 35250 37748 35256 37760
rect 35308 37748 35314 37800
rect 56502 37748 56508 37800
rect 56560 37788 56566 37800
rect 56597 37791 56655 37797
rect 56597 37788 56609 37791
rect 56560 37760 56609 37788
rect 56560 37748 56566 37760
rect 56597 37757 56609 37760
rect 56643 37757 56655 37791
rect 57422 37788 57428 37800
rect 57383 37760 57428 37788
rect 56597 37751 56655 37757
rect 57422 37748 57428 37760
rect 57480 37748 57486 37800
rect 1302 37680 1308 37732
rect 1360 37720 1366 37732
rect 19705 37723 19763 37729
rect 19705 37720 19717 37723
rect 1360 37692 19717 37720
rect 1360 37680 1366 37692
rect 19705 37689 19717 37692
rect 19751 37689 19763 37723
rect 19705 37683 19763 37689
rect 33042 37680 33048 37732
rect 33100 37720 33106 37732
rect 33137 37723 33195 37729
rect 33137 37720 33149 37723
rect 33100 37692 33149 37720
rect 33100 37680 33106 37692
rect 33137 37689 33149 37692
rect 33183 37689 33195 37723
rect 33502 37720 33508 37732
rect 33463 37692 33508 37720
rect 33137 37683 33195 37689
rect 33502 37680 33508 37692
rect 33560 37680 33566 37732
rect 57977 37723 58035 37729
rect 57977 37689 57989 37723
rect 58023 37720 58035 37723
rect 58710 37720 58716 37732
rect 58023 37692 58716 37720
rect 58023 37689 58035 37692
rect 57977 37683 58035 37689
rect 58710 37680 58716 37692
rect 58768 37680 58774 37732
rect 16206 37652 16212 37664
rect 16167 37624 16212 37652
rect 16206 37612 16212 37624
rect 16264 37612 16270 37664
rect 17497 37655 17555 37661
rect 17497 37621 17509 37655
rect 17543 37652 17555 37655
rect 18690 37652 18696 37664
rect 17543 37624 18696 37652
rect 17543 37621 17555 37624
rect 17497 37615 17555 37621
rect 18690 37612 18696 37624
rect 18748 37612 18754 37664
rect 20990 37652 20996 37664
rect 20951 37624 20996 37652
rect 20990 37612 20996 37624
rect 21048 37612 21054 37664
rect 27985 37655 28043 37661
rect 27985 37621 27997 37655
rect 28031 37652 28043 37655
rect 28534 37652 28540 37664
rect 28031 37624 28540 37652
rect 28031 37621 28043 37624
rect 27985 37615 28043 37621
rect 28534 37612 28540 37624
rect 28592 37612 28598 37664
rect 34514 37652 34520 37664
rect 34475 37624 34520 37652
rect 34514 37612 34520 37624
rect 34572 37612 34578 37664
rect 1104 37562 58880 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 58880 37562
rect 1104 37488 58880 37510
rect 16390 37408 16396 37460
rect 16448 37448 16454 37460
rect 17954 37448 17960 37460
rect 16448 37420 17960 37448
rect 16448 37408 16454 37420
rect 17954 37408 17960 37420
rect 18012 37408 18018 37460
rect 18690 37408 18696 37460
rect 18748 37448 18754 37460
rect 18785 37451 18843 37457
rect 18785 37448 18797 37451
rect 18748 37420 18797 37448
rect 18748 37408 18754 37420
rect 18785 37417 18797 37420
rect 18831 37417 18843 37451
rect 18785 37411 18843 37417
rect 20165 37451 20223 37457
rect 20165 37417 20177 37451
rect 20211 37448 20223 37451
rect 20438 37448 20444 37460
rect 20211 37420 20444 37448
rect 20211 37417 20223 37420
rect 20165 37411 20223 37417
rect 20438 37408 20444 37420
rect 20496 37408 20502 37460
rect 20625 37451 20683 37457
rect 20625 37417 20637 37451
rect 20671 37448 20683 37451
rect 20714 37448 20720 37460
rect 20671 37420 20720 37448
rect 20671 37417 20683 37420
rect 20625 37411 20683 37417
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 34790 37448 34796 37460
rect 34751 37420 34796 37448
rect 34790 37408 34796 37420
rect 34848 37408 34854 37460
rect 57882 37408 57888 37460
rect 57940 37448 57946 37460
rect 58069 37451 58127 37457
rect 58069 37448 58081 37451
rect 57940 37420 58081 37448
rect 57940 37408 57946 37420
rect 58069 37417 58081 37420
rect 58115 37417 58127 37451
rect 58069 37411 58127 37417
rect 15746 37380 15752 37392
rect 15120 37352 15752 37380
rect 1394 37312 1400 37324
rect 1355 37284 1400 37312
rect 1394 37272 1400 37284
rect 1452 37272 1458 37324
rect 15120 37321 15148 37352
rect 15746 37340 15752 37352
rect 15804 37340 15810 37392
rect 18141 37383 18199 37389
rect 18141 37349 18153 37383
rect 18187 37380 18199 37383
rect 18598 37380 18604 37392
rect 18187 37352 18604 37380
rect 18187 37349 18199 37352
rect 18141 37343 18199 37349
rect 18598 37340 18604 37352
rect 18656 37380 18662 37392
rect 18656 37352 18736 37380
rect 18656 37340 18662 37352
rect 14921 37315 14979 37321
rect 14921 37281 14933 37315
rect 14967 37312 14979 37315
rect 15105 37315 15163 37321
rect 14967 37284 15056 37312
rect 14967 37281 14979 37284
rect 14921 37275 14979 37281
rect 15028 37176 15056 37284
rect 15105 37281 15117 37315
rect 15151 37281 15163 37315
rect 15654 37312 15660 37324
rect 15615 37284 15660 37312
rect 15105 37275 15163 37281
rect 15654 37272 15660 37284
rect 15712 37272 15718 37324
rect 16301 37315 16359 37321
rect 16301 37312 16313 37315
rect 15856 37284 16313 37312
rect 15194 37244 15200 37256
rect 15155 37216 15200 37244
rect 15194 37204 15200 37216
rect 15252 37204 15258 37256
rect 15856 37188 15884 37284
rect 16301 37281 16313 37284
rect 16347 37281 16359 37315
rect 16301 37275 16359 37281
rect 16393 37315 16451 37321
rect 16393 37281 16405 37315
rect 16439 37312 16451 37315
rect 16942 37312 16948 37324
rect 16439 37284 16948 37312
rect 16439 37281 16451 37284
rect 16393 37275 16451 37281
rect 16942 37272 16948 37284
rect 17000 37272 17006 37324
rect 17126 37312 17132 37324
rect 17087 37284 17132 37312
rect 17126 37272 17132 37284
rect 17184 37272 17190 37324
rect 18046 37312 18052 37324
rect 18007 37284 18052 37312
rect 18046 37272 18052 37284
rect 18104 37272 18110 37324
rect 18230 37312 18236 37324
rect 18191 37284 18236 37312
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 18708 37321 18736 37352
rect 28074 37340 28080 37392
rect 28132 37380 28138 37392
rect 28445 37383 28503 37389
rect 28445 37380 28457 37383
rect 28132 37352 28457 37380
rect 28132 37340 28138 37352
rect 28445 37349 28457 37352
rect 28491 37380 28503 37383
rect 28491 37352 29040 37380
rect 28491 37349 28503 37352
rect 28445 37343 28503 37349
rect 18693 37315 18751 37321
rect 18693 37281 18705 37315
rect 18739 37281 18751 37315
rect 18693 37275 18751 37281
rect 19886 37272 19892 37324
rect 19944 37312 19950 37324
rect 19981 37315 20039 37321
rect 19981 37312 19993 37315
rect 19944 37284 19993 37312
rect 19944 37272 19950 37284
rect 19981 37281 19993 37284
rect 20027 37281 20039 37315
rect 19981 37275 20039 37281
rect 20070 37272 20076 37324
rect 20128 37312 20134 37324
rect 20165 37315 20223 37321
rect 20165 37312 20177 37315
rect 20128 37284 20177 37312
rect 20128 37272 20134 37284
rect 20165 37281 20177 37284
rect 20211 37281 20223 37315
rect 20165 37275 20223 37281
rect 20714 37272 20720 37324
rect 20772 37312 20778 37324
rect 20809 37315 20867 37321
rect 20809 37312 20821 37315
rect 20772 37284 20821 37312
rect 20772 37272 20778 37284
rect 20809 37281 20821 37284
rect 20855 37281 20867 37315
rect 20809 37275 20867 37281
rect 28353 37315 28411 37321
rect 28353 37281 28365 37315
rect 28399 37281 28411 37315
rect 28353 37275 28411 37281
rect 28537 37315 28595 37321
rect 28537 37281 28549 37315
rect 28583 37312 28595 37315
rect 28626 37312 28632 37324
rect 28583 37284 28632 37312
rect 28583 37281 28595 37284
rect 28537 37275 28595 37281
rect 28258 37204 28264 37256
rect 28316 37244 28322 37256
rect 28368 37244 28396 37275
rect 28626 37272 28632 37284
rect 28684 37272 28690 37324
rect 29012 37321 29040 37352
rect 31128 37352 33180 37380
rect 28997 37315 29055 37321
rect 28997 37281 29009 37315
rect 29043 37281 29055 37315
rect 28997 37275 29055 37281
rect 29089 37315 29147 37321
rect 29089 37281 29101 37315
rect 29135 37312 29147 37315
rect 30466 37312 30472 37324
rect 29135 37284 30472 37312
rect 29135 37281 29147 37284
rect 29089 37275 29147 37281
rect 30466 37272 30472 37284
rect 30524 37272 30530 37324
rect 30650 37312 30656 37324
rect 30611 37284 30656 37312
rect 30650 37272 30656 37284
rect 30708 37272 30714 37324
rect 30926 37272 30932 37324
rect 30984 37312 30990 37324
rect 31128 37321 31156 37352
rect 33152 37324 33180 37352
rect 33502 37340 33508 37392
rect 33560 37380 33566 37392
rect 33658 37383 33716 37389
rect 33658 37380 33670 37383
rect 33560 37352 33670 37380
rect 33560 37340 33566 37352
rect 33658 37349 33670 37352
rect 33704 37349 33716 37383
rect 33658 37343 33716 37349
rect 31113 37315 31171 37321
rect 31113 37312 31125 37315
rect 30984 37284 31125 37312
rect 30984 37272 30990 37284
rect 31113 37281 31125 37284
rect 31159 37281 31171 37315
rect 31113 37275 31171 37281
rect 31380 37315 31438 37321
rect 31380 37281 31392 37315
rect 31426 37312 31438 37315
rect 32214 37312 32220 37324
rect 31426 37284 32220 37312
rect 31426 37281 31438 37284
rect 31380 37275 31438 37281
rect 32214 37272 32220 37284
rect 32272 37272 32278 37324
rect 33134 37272 33140 37324
rect 33192 37312 33198 37324
rect 33410 37312 33416 37324
rect 33192 37284 33416 37312
rect 33192 37272 33198 37284
rect 33410 37272 33416 37284
rect 33468 37272 33474 37324
rect 56778 37272 56784 37324
rect 56836 37312 56842 37324
rect 56962 37312 56968 37324
rect 56836 37284 56968 37312
rect 56836 37272 56842 37284
rect 56962 37272 56968 37284
rect 57020 37312 57026 37324
rect 57241 37315 57299 37321
rect 57241 37312 57253 37315
rect 57020 37284 57253 37312
rect 57020 37272 57026 37284
rect 57241 37281 57253 37284
rect 57287 37281 57299 37315
rect 57974 37312 57980 37324
rect 57935 37284 57980 37312
rect 57241 37275 57299 37281
rect 57974 37272 57980 37284
rect 58032 37272 58038 37324
rect 28718 37244 28724 37256
rect 28316 37216 28724 37244
rect 28316 37204 28322 37216
rect 28718 37204 28724 37216
rect 28776 37204 28782 37256
rect 15838 37176 15844 37188
rect 15028 37148 15844 37176
rect 15838 37136 15844 37148
rect 15896 37136 15902 37188
rect 14734 37108 14740 37120
rect 14695 37080 14740 37108
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 17037 37111 17095 37117
rect 17037 37077 17049 37111
rect 17083 37108 17095 37111
rect 17678 37108 17684 37120
rect 17083 37080 17684 37108
rect 17083 37077 17095 37080
rect 17037 37071 17095 37077
rect 17678 37068 17684 37080
rect 17736 37068 17742 37120
rect 30558 37108 30564 37120
rect 30519 37080 30564 37108
rect 30558 37068 30564 37080
rect 30616 37068 30622 37120
rect 32490 37108 32496 37120
rect 32451 37080 32496 37108
rect 32490 37068 32496 37080
rect 32548 37068 32554 37120
rect 57422 37108 57428 37120
rect 57383 37080 57428 37108
rect 57422 37068 57428 37080
rect 57480 37068 57486 37120
rect 1104 37018 58880 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 58880 37018
rect 1104 36944 58880 36966
rect 15194 36864 15200 36916
rect 15252 36904 15258 36916
rect 15289 36907 15347 36913
rect 15289 36904 15301 36907
rect 15252 36876 15301 36904
rect 15252 36864 15258 36876
rect 15289 36873 15301 36876
rect 15335 36873 15347 36907
rect 15838 36904 15844 36916
rect 15799 36876 15844 36904
rect 15289 36867 15347 36873
rect 15304 36768 15332 36867
rect 15838 36864 15844 36876
rect 15896 36864 15902 36916
rect 18230 36864 18236 36916
rect 18288 36904 18294 36916
rect 18874 36904 18880 36916
rect 18288 36876 18880 36904
rect 18288 36864 18294 36876
rect 18874 36864 18880 36876
rect 18932 36904 18938 36916
rect 18969 36907 19027 36913
rect 18969 36904 18981 36907
rect 18932 36876 18981 36904
rect 18932 36864 18938 36876
rect 18969 36873 18981 36876
rect 19015 36873 19027 36907
rect 28258 36904 28264 36916
rect 28219 36876 28264 36904
rect 18969 36867 19027 36873
rect 28258 36864 28264 36876
rect 28316 36864 28322 36916
rect 30466 36864 30472 36916
rect 30524 36904 30530 36916
rect 31205 36907 31263 36913
rect 31205 36904 31217 36907
rect 30524 36876 31217 36904
rect 30524 36864 30530 36876
rect 31205 36873 31217 36876
rect 31251 36873 31263 36907
rect 57974 36904 57980 36916
rect 57935 36876 57980 36904
rect 31205 36867 31263 36873
rect 57974 36864 57980 36876
rect 58032 36864 58038 36916
rect 30377 36839 30435 36845
rect 30377 36805 30389 36839
rect 30423 36836 30435 36839
rect 30650 36836 30656 36848
rect 30423 36808 30656 36836
rect 30423 36805 30435 36808
rect 30377 36799 30435 36805
rect 30650 36796 30656 36808
rect 30708 36836 30714 36848
rect 33229 36839 33287 36845
rect 30708 36808 31340 36836
rect 30708 36796 30714 36808
rect 17586 36768 17592 36780
rect 15304 36740 15976 36768
rect 17547 36740 17592 36768
rect 13722 36660 13728 36712
rect 13780 36700 13786 36712
rect 13909 36703 13967 36709
rect 13909 36700 13921 36703
rect 13780 36672 13921 36700
rect 13780 36660 13786 36672
rect 13909 36669 13921 36672
rect 13955 36669 13967 36703
rect 13909 36663 13967 36669
rect 14176 36703 14234 36709
rect 14176 36669 14188 36703
rect 14222 36700 14234 36703
rect 14734 36700 14740 36712
rect 14222 36672 14740 36700
rect 14222 36669 14234 36672
rect 14176 36663 14234 36669
rect 13924 36632 13952 36663
rect 14734 36660 14740 36672
rect 14792 36660 14798 36712
rect 15746 36700 15752 36712
rect 15707 36672 15752 36700
rect 15746 36660 15752 36672
rect 15804 36660 15810 36712
rect 15948 36709 15976 36740
rect 17586 36728 17592 36740
rect 17644 36728 17650 36780
rect 30926 36768 30932 36780
rect 30024 36740 30932 36768
rect 15933 36703 15991 36709
rect 15933 36669 15945 36703
rect 15979 36669 15991 36703
rect 28074 36700 28080 36712
rect 28035 36672 28080 36700
rect 15933 36663 15991 36669
rect 28074 36660 28080 36672
rect 28132 36660 28138 36712
rect 28353 36703 28411 36709
rect 28353 36669 28365 36703
rect 28399 36700 28411 36703
rect 28626 36700 28632 36712
rect 28399 36672 28632 36700
rect 28399 36669 28411 36672
rect 28353 36663 28411 36669
rect 28626 36660 28632 36672
rect 28684 36660 28690 36712
rect 28997 36703 29055 36709
rect 28997 36669 29009 36703
rect 29043 36700 29055 36703
rect 30024 36700 30052 36740
rect 30926 36728 30932 36740
rect 30984 36728 30990 36780
rect 31312 36777 31340 36808
rect 33229 36805 33241 36839
rect 33275 36836 33287 36839
rect 34514 36836 34520 36848
rect 33275 36808 34520 36836
rect 33275 36805 33287 36808
rect 33229 36799 33287 36805
rect 34514 36796 34520 36808
rect 34572 36796 34578 36848
rect 31297 36771 31355 36777
rect 31297 36737 31309 36771
rect 31343 36737 31355 36771
rect 33778 36768 33784 36780
rect 31297 36731 31355 36737
rect 33152 36740 33784 36768
rect 29043 36672 30052 36700
rect 29043 36669 29055 36672
rect 28997 36663 29055 36669
rect 30558 36660 30564 36712
rect 30616 36700 30622 36712
rect 31021 36703 31079 36709
rect 31021 36700 31033 36703
rect 30616 36672 31033 36700
rect 30616 36660 30622 36672
rect 31021 36669 31033 36672
rect 31067 36669 31079 36703
rect 31021 36663 31079 36669
rect 31941 36703 31999 36709
rect 31941 36669 31953 36703
rect 31987 36700 31999 36703
rect 32490 36700 32496 36712
rect 31987 36672 32496 36700
rect 31987 36669 31999 36672
rect 31941 36663 31999 36669
rect 32490 36660 32496 36672
rect 32548 36660 32554 36712
rect 33152 36709 33180 36740
rect 33778 36728 33784 36740
rect 33836 36728 33842 36780
rect 33137 36703 33195 36709
rect 33137 36669 33149 36703
rect 33183 36669 33195 36703
rect 33137 36663 33195 36669
rect 33413 36703 33471 36709
rect 33413 36669 33425 36703
rect 33459 36669 33471 36703
rect 33413 36663 33471 36669
rect 56321 36703 56379 36709
rect 56321 36669 56333 36703
rect 56367 36700 56379 36703
rect 57517 36703 57575 36709
rect 57517 36700 57529 36703
rect 56367 36672 57529 36700
rect 56367 36669 56379 36672
rect 56321 36663 56379 36669
rect 57517 36669 57529 36672
rect 57563 36669 57575 36703
rect 57698 36700 57704 36712
rect 57659 36672 57704 36700
rect 57517 36663 57575 36669
rect 16206 36632 16212 36644
rect 13924 36604 16212 36632
rect 16206 36592 16212 36604
rect 16264 36592 16270 36644
rect 17856 36635 17914 36641
rect 17856 36601 17868 36635
rect 17902 36632 17914 36635
rect 18414 36632 18420 36644
rect 17902 36604 18420 36632
rect 17902 36601 17914 36604
rect 17856 36595 17914 36601
rect 18414 36592 18420 36604
rect 18472 36592 18478 36644
rect 29264 36635 29322 36641
rect 29264 36601 29276 36635
rect 29310 36632 29322 36635
rect 30837 36635 30895 36641
rect 30837 36632 30849 36635
rect 29310 36604 30849 36632
rect 29310 36601 29322 36604
rect 29264 36595 29322 36601
rect 30837 36601 30849 36604
rect 30883 36601 30895 36635
rect 33428 36632 33456 36663
rect 57698 36660 57704 36672
rect 57756 36660 57762 36712
rect 30837 36595 30895 36601
rect 32784 36604 33456 36632
rect 56873 36635 56931 36641
rect 32784 36576 32812 36604
rect 56873 36601 56885 36635
rect 56919 36601 56931 36635
rect 57054 36632 57060 36644
rect 57015 36604 57060 36632
rect 56873 36595 56931 36601
rect 27890 36564 27896 36576
rect 27851 36536 27896 36564
rect 27890 36524 27896 36536
rect 27948 36524 27954 36576
rect 32033 36567 32091 36573
rect 32033 36533 32045 36567
rect 32079 36564 32091 36567
rect 32766 36564 32772 36576
rect 32079 36536 32772 36564
rect 32079 36533 32091 36536
rect 32033 36527 32091 36533
rect 32766 36524 32772 36536
rect 32824 36524 32830 36576
rect 33042 36524 33048 36576
rect 33100 36564 33106 36576
rect 33597 36567 33655 36573
rect 33597 36564 33609 36567
rect 33100 36536 33609 36564
rect 33100 36524 33106 36536
rect 33597 36533 33609 36536
rect 33643 36533 33655 36567
rect 56888 36564 56916 36595
rect 57054 36592 57060 36604
rect 57112 36592 57118 36644
rect 56962 36564 56968 36576
rect 56888 36536 56968 36564
rect 33597 36527 33655 36533
rect 56962 36524 56968 36536
rect 57020 36524 57026 36576
rect 1104 36474 58880 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 58880 36474
rect 1104 36400 58880 36422
rect 17037 36363 17095 36369
rect 17037 36329 17049 36363
rect 17083 36360 17095 36363
rect 17126 36360 17132 36372
rect 17083 36332 17132 36360
rect 17083 36329 17095 36332
rect 17037 36323 17095 36329
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 18414 36360 18420 36372
rect 18375 36332 18420 36360
rect 18414 36320 18420 36332
rect 18472 36320 18478 36372
rect 28626 36360 28632 36372
rect 28587 36332 28632 36360
rect 28626 36320 28632 36332
rect 28684 36320 28690 36372
rect 32214 36360 32220 36372
rect 32175 36332 32220 36360
rect 32214 36320 32220 36332
rect 32272 36320 32278 36372
rect 33229 36363 33287 36369
rect 33229 36329 33241 36363
rect 33275 36360 33287 36363
rect 33318 36360 33324 36372
rect 33275 36332 33324 36360
rect 33275 36329 33287 36332
rect 33229 36323 33287 36329
rect 33318 36320 33324 36332
rect 33376 36320 33382 36372
rect 57241 36363 57299 36369
rect 57241 36329 57253 36363
rect 57287 36360 57299 36363
rect 57698 36360 57704 36372
rect 57287 36332 57704 36360
rect 57287 36329 57299 36332
rect 57241 36323 57299 36329
rect 57698 36320 57704 36332
rect 57756 36320 57762 36372
rect 16206 36292 16212 36304
rect 15672 36264 16212 36292
rect 1394 36224 1400 36236
rect 1355 36196 1400 36224
rect 1394 36184 1400 36196
rect 1452 36184 1458 36236
rect 15672 36233 15700 36264
rect 16206 36252 16212 36264
rect 16264 36252 16270 36304
rect 17144 36292 17172 36320
rect 27516 36295 27574 36301
rect 17144 36264 18000 36292
rect 15657 36227 15715 36233
rect 15657 36193 15669 36227
rect 15703 36193 15715 36227
rect 15657 36187 15715 36193
rect 15924 36227 15982 36233
rect 15924 36193 15936 36227
rect 15970 36224 15982 36227
rect 17497 36227 17555 36233
rect 17497 36224 17509 36227
rect 15970 36196 17509 36224
rect 15970 36193 15982 36196
rect 15924 36187 15982 36193
rect 17497 36193 17509 36196
rect 17543 36193 17555 36227
rect 17678 36224 17684 36236
rect 17639 36196 17684 36224
rect 17497 36187 17555 36193
rect 17678 36184 17684 36196
rect 17736 36184 17742 36236
rect 17972 36233 18000 36264
rect 27516 36261 27528 36295
rect 27562 36292 27574 36295
rect 27890 36292 27896 36304
rect 27562 36264 27896 36292
rect 27562 36261 27574 36264
rect 27516 36255 27574 36261
rect 27890 36252 27896 36264
rect 27948 36252 27954 36304
rect 34514 36292 34520 36304
rect 33428 36264 34520 36292
rect 17957 36227 18015 36233
rect 17957 36193 17969 36227
rect 18003 36193 18015 36227
rect 18598 36224 18604 36236
rect 18559 36196 18604 36224
rect 17957 36187 18015 36193
rect 18598 36184 18604 36196
rect 18656 36184 18662 36236
rect 18874 36224 18880 36236
rect 18835 36196 18880 36224
rect 18874 36184 18880 36196
rect 18932 36184 18938 36236
rect 30469 36227 30527 36233
rect 30469 36193 30481 36227
rect 30515 36224 30527 36227
rect 30558 36224 30564 36236
rect 30515 36196 30564 36224
rect 30515 36193 30527 36196
rect 30469 36187 30527 36193
rect 30558 36184 30564 36196
rect 30616 36184 30622 36236
rect 32398 36224 32404 36236
rect 32359 36196 32404 36224
rect 32398 36184 32404 36196
rect 32456 36184 32462 36236
rect 32493 36227 32551 36233
rect 32493 36193 32505 36227
rect 32539 36193 32551 36227
rect 32766 36224 32772 36236
rect 32727 36196 32772 36224
rect 32493 36187 32551 36193
rect 16942 36116 16948 36168
rect 17000 36156 17006 36168
rect 17865 36159 17923 36165
rect 17865 36156 17877 36159
rect 17000 36128 17877 36156
rect 17000 36116 17006 36128
rect 17865 36125 17877 36128
rect 17911 36125 17923 36159
rect 27246 36156 27252 36168
rect 27207 36128 27252 36156
rect 17865 36119 17923 36125
rect 27246 36116 27252 36128
rect 27304 36116 27310 36168
rect 32508 36088 32536 36187
rect 32766 36184 32772 36196
rect 32824 36184 32830 36236
rect 33428 36233 33456 36264
rect 34514 36252 34520 36264
rect 34572 36252 34578 36304
rect 33413 36227 33471 36233
rect 33413 36193 33425 36227
rect 33459 36193 33471 36227
rect 33413 36187 33471 36193
rect 33778 36184 33784 36236
rect 33836 36224 33842 36236
rect 34149 36227 34207 36233
rect 34149 36224 34161 36227
rect 33836 36196 34161 36224
rect 33836 36184 33842 36196
rect 34149 36193 34161 36196
rect 34195 36193 34207 36227
rect 57422 36224 57428 36236
rect 57383 36196 57428 36224
rect 34149 36187 34207 36193
rect 57422 36184 57428 36196
rect 57480 36184 57486 36236
rect 57974 36224 57980 36236
rect 57935 36196 57980 36224
rect 57974 36184 57980 36196
rect 58032 36184 58038 36236
rect 32784 36156 32812 36184
rect 33689 36159 33747 36165
rect 33689 36156 33701 36159
rect 32784 36128 33701 36156
rect 33689 36125 33701 36128
rect 33735 36125 33747 36159
rect 33689 36119 33747 36125
rect 34238 36088 34244 36100
rect 32508 36060 34244 36088
rect 34238 36048 34244 36060
rect 34296 36048 34302 36100
rect 18782 36020 18788 36032
rect 18743 35992 18788 36020
rect 18782 35980 18788 35992
rect 18840 35980 18846 36032
rect 30561 36023 30619 36029
rect 30561 35989 30573 36023
rect 30607 36020 30619 36023
rect 31110 36020 31116 36032
rect 30607 35992 31116 36020
rect 30607 35989 30619 35992
rect 30561 35983 30619 35989
rect 31110 35980 31116 35992
rect 31168 35980 31174 36032
rect 32677 36023 32735 36029
rect 32677 35989 32689 36023
rect 32723 36020 32735 36023
rect 33597 36023 33655 36029
rect 33597 36020 33609 36023
rect 32723 35992 33609 36020
rect 32723 35989 32735 35992
rect 32677 35983 32735 35989
rect 33597 35989 33609 35992
rect 33643 36020 33655 36023
rect 33686 36020 33692 36032
rect 33643 35992 33692 36020
rect 33643 35989 33655 35992
rect 33597 35983 33655 35989
rect 33686 35980 33692 35992
rect 33744 35980 33750 36032
rect 57882 35980 57888 36032
rect 57940 36020 57946 36032
rect 58069 36023 58127 36029
rect 58069 36020 58081 36023
rect 57940 35992 58081 36020
rect 57940 35980 57946 35992
rect 58069 35989 58081 35992
rect 58115 35989 58127 36023
rect 58069 35983 58127 35989
rect 1104 35930 58880 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 58880 35930
rect 1104 35856 58880 35878
rect 17589 35819 17647 35825
rect 17589 35785 17601 35819
rect 17635 35816 17647 35819
rect 18046 35816 18052 35828
rect 17635 35788 18052 35816
rect 17635 35785 17647 35788
rect 17589 35779 17647 35785
rect 18046 35776 18052 35788
rect 18104 35816 18110 35828
rect 18782 35816 18788 35828
rect 18104 35788 18788 35816
rect 18104 35776 18110 35788
rect 18782 35776 18788 35788
rect 18840 35776 18846 35828
rect 31110 35816 31116 35828
rect 31071 35788 31116 35816
rect 31110 35776 31116 35788
rect 31168 35776 31174 35828
rect 57974 35816 57980 35828
rect 57935 35788 57980 35816
rect 57974 35776 57980 35788
rect 58032 35776 58038 35828
rect 17954 35708 17960 35760
rect 18012 35748 18018 35760
rect 18141 35751 18199 35757
rect 18141 35748 18153 35751
rect 18012 35720 18153 35748
rect 18012 35708 18018 35720
rect 18141 35717 18153 35720
rect 18187 35717 18199 35751
rect 18141 35711 18199 35717
rect 31128 35680 31156 35776
rect 33134 35680 33140 35692
rect 31128 35652 31708 35680
rect 33095 35652 33140 35680
rect 1394 35612 1400 35624
rect 1355 35584 1400 35612
rect 1394 35572 1400 35584
rect 1452 35572 1458 35624
rect 17497 35615 17555 35621
rect 17497 35581 17509 35615
rect 17543 35612 17555 35615
rect 17678 35612 17684 35624
rect 17543 35584 17684 35612
rect 17543 35581 17555 35584
rect 17497 35575 17555 35581
rect 17678 35572 17684 35584
rect 17736 35572 17742 35624
rect 18322 35612 18328 35624
rect 18283 35584 18328 35612
rect 18322 35572 18328 35584
rect 18380 35572 18386 35624
rect 31680 35621 31708 35652
rect 33134 35640 33140 35652
rect 33192 35640 33198 35692
rect 34238 35640 34244 35692
rect 34296 35680 34302 35692
rect 34296 35652 35204 35680
rect 34296 35640 34302 35652
rect 30929 35615 30987 35621
rect 30929 35581 30941 35615
rect 30975 35581 30987 35615
rect 30929 35575 30987 35581
rect 31205 35615 31263 35621
rect 31205 35581 31217 35615
rect 31251 35581 31263 35615
rect 31205 35575 31263 35581
rect 31665 35615 31723 35621
rect 31665 35581 31677 35615
rect 31711 35581 31723 35615
rect 31846 35612 31852 35624
rect 31807 35584 31852 35612
rect 31665 35575 31723 35581
rect 30742 35476 30748 35488
rect 30703 35448 30748 35476
rect 30742 35436 30748 35448
rect 30800 35436 30806 35488
rect 30944 35476 30972 35575
rect 31220 35544 31248 35575
rect 31846 35572 31852 35584
rect 31904 35572 31910 35624
rect 34974 35612 34980 35624
rect 34935 35584 34980 35612
rect 34974 35572 34980 35584
rect 35032 35572 35038 35624
rect 35176 35621 35204 35652
rect 35161 35615 35219 35621
rect 35161 35581 35173 35615
rect 35207 35581 35219 35615
rect 56226 35612 56232 35624
rect 56187 35584 56232 35612
rect 35161 35575 35219 35581
rect 56226 35572 56232 35584
rect 56284 35572 56290 35624
rect 57057 35615 57115 35621
rect 57057 35581 57069 35615
rect 57103 35612 57115 35615
rect 57517 35615 57575 35621
rect 57517 35612 57529 35615
rect 57103 35584 57529 35612
rect 57103 35581 57115 35584
rect 57057 35575 57115 35581
rect 57517 35581 57529 35584
rect 57563 35581 57575 35615
rect 57698 35612 57704 35624
rect 57659 35584 57704 35612
rect 57517 35575 57575 35581
rect 57698 35572 57704 35584
rect 57756 35572 57762 35624
rect 31864 35544 31892 35572
rect 31220 35516 31892 35544
rect 33404 35547 33462 35553
rect 33404 35513 33416 35547
rect 33450 35544 33462 35547
rect 35069 35547 35127 35553
rect 35069 35544 35081 35547
rect 33450 35516 35081 35544
rect 33450 35513 33462 35516
rect 33404 35507 33462 35513
rect 35069 35513 35081 35516
rect 35115 35513 35127 35547
rect 35069 35507 35127 35513
rect 31754 35476 31760 35488
rect 30944 35448 31760 35476
rect 31754 35436 31760 35448
rect 31812 35476 31818 35488
rect 31812 35448 31857 35476
rect 31812 35436 31818 35448
rect 34422 35436 34428 35488
rect 34480 35476 34486 35488
rect 34517 35479 34575 35485
rect 34517 35476 34529 35479
rect 34480 35448 34529 35476
rect 34480 35436 34486 35448
rect 34517 35445 34529 35448
rect 34563 35445 34575 35479
rect 34517 35439 34575 35445
rect 1104 35386 58880 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 58880 35386
rect 1104 35312 58880 35334
rect 31846 35272 31852 35284
rect 31807 35244 31852 35272
rect 31846 35232 31852 35244
rect 31904 35232 31910 35284
rect 32309 35275 32367 35281
rect 32309 35241 32321 35275
rect 32355 35272 32367 35275
rect 34974 35272 34980 35284
rect 32355 35244 34980 35272
rect 32355 35241 32367 35244
rect 32309 35235 32367 35241
rect 34974 35232 34980 35244
rect 35032 35232 35038 35284
rect 57241 35275 57299 35281
rect 57241 35241 57253 35275
rect 57287 35272 57299 35275
rect 57698 35272 57704 35284
rect 57287 35244 57704 35272
rect 57287 35241 57299 35244
rect 57241 35235 57299 35241
rect 57698 35232 57704 35244
rect 57756 35232 57762 35284
rect 30742 35213 30748 35216
rect 30736 35204 30748 35213
rect 30703 35176 30748 35204
rect 30736 35167 30748 35176
rect 30742 35164 30748 35167
rect 30800 35164 30806 35216
rect 18322 35096 18328 35148
rect 18380 35136 18386 35148
rect 20165 35139 20223 35145
rect 20165 35136 20177 35139
rect 18380 35108 20177 35136
rect 18380 35096 18386 35108
rect 20165 35105 20177 35108
rect 20211 35105 20223 35139
rect 20165 35099 20223 35105
rect 32493 35139 32551 35145
rect 32493 35105 32505 35139
rect 32539 35105 32551 35139
rect 32493 35099 32551 35105
rect 32677 35139 32735 35145
rect 32677 35105 32689 35139
rect 32723 35136 32735 35139
rect 33226 35136 33232 35148
rect 32723 35108 33232 35136
rect 32723 35105 32735 35108
rect 32677 35099 32735 35105
rect 27246 35028 27252 35080
rect 27304 35068 27310 35080
rect 30466 35068 30472 35080
rect 27304 35040 30472 35068
rect 27304 35028 27310 35040
rect 30466 35028 30472 35040
rect 30524 35028 30530 35080
rect 32508 35000 32536 35099
rect 33226 35096 33232 35108
rect 33284 35096 33290 35148
rect 33505 35139 33563 35145
rect 33505 35105 33517 35139
rect 33551 35136 33563 35139
rect 33778 35136 33784 35148
rect 33551 35108 33784 35136
rect 33551 35105 33563 35108
rect 33505 35099 33563 35105
rect 32769 35071 32827 35077
rect 32769 35037 32781 35071
rect 32815 35068 32827 35071
rect 33520 35068 33548 35099
rect 33778 35096 33784 35108
rect 33836 35096 33842 35148
rect 34422 35136 34428 35148
rect 34383 35108 34428 35136
rect 34422 35096 34428 35108
rect 34480 35096 34486 35148
rect 57422 35136 57428 35148
rect 57383 35108 57428 35136
rect 57422 35096 57428 35108
rect 57480 35096 57486 35148
rect 57514 35096 57520 35148
rect 57572 35136 57578 35148
rect 57698 35136 57704 35148
rect 57572 35108 57704 35136
rect 57572 35096 57578 35108
rect 57698 35096 57704 35108
rect 57756 35096 57762 35148
rect 57977 35139 58035 35145
rect 57977 35105 57989 35139
rect 58023 35136 58035 35139
rect 58066 35136 58072 35148
rect 58023 35108 58072 35136
rect 58023 35105 58035 35108
rect 57977 35099 58035 35105
rect 58066 35096 58072 35108
rect 58124 35096 58130 35148
rect 33686 35068 33692 35080
rect 32815 35040 33548 35068
rect 33647 35040 33692 35068
rect 32815 35037 32827 35040
rect 32769 35031 32827 35037
rect 33686 35028 33692 35040
rect 33744 35028 33750 35080
rect 33321 35003 33379 35009
rect 33321 35000 33333 35003
rect 32508 34972 33333 35000
rect 33321 34969 33333 34972
rect 33367 35000 33379 35003
rect 34517 35003 34575 35009
rect 34517 35000 34529 35003
rect 33367 34972 34529 35000
rect 33367 34969 33379 34972
rect 33321 34963 33379 34969
rect 34517 34969 34529 34972
rect 34563 34969 34575 35003
rect 58158 35000 58164 35012
rect 58119 34972 58164 35000
rect 34517 34963 34575 34969
rect 58158 34960 58164 34972
rect 58216 34960 58222 35012
rect 19981 34935 20039 34941
rect 19981 34901 19993 34935
rect 20027 34932 20039 34935
rect 20714 34932 20720 34944
rect 20027 34904 20720 34932
rect 20027 34901 20039 34904
rect 19981 34895 20039 34901
rect 20714 34892 20720 34904
rect 20772 34892 20778 34944
rect 1104 34842 58880 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 58880 34842
rect 1104 34768 58880 34790
rect 17681 34731 17739 34737
rect 17681 34697 17693 34731
rect 17727 34728 17739 34731
rect 18322 34728 18328 34740
rect 17727 34700 18328 34728
rect 17727 34697 17739 34700
rect 17681 34691 17739 34697
rect 18322 34688 18328 34700
rect 18380 34688 18386 34740
rect 22557 34731 22615 34737
rect 22557 34697 22569 34731
rect 22603 34728 22615 34731
rect 27246 34728 27252 34740
rect 22603 34700 27252 34728
rect 22603 34697 22615 34700
rect 22557 34691 22615 34697
rect 27246 34688 27252 34700
rect 27304 34688 27310 34740
rect 33226 34688 33232 34740
rect 33284 34728 33290 34740
rect 33505 34731 33563 34737
rect 33505 34728 33517 34731
rect 33284 34700 33517 34728
rect 33284 34688 33290 34700
rect 33505 34697 33517 34700
rect 33551 34728 33563 34731
rect 34146 34728 34152 34740
rect 33551 34700 34152 34728
rect 33551 34697 33563 34700
rect 33505 34691 33563 34697
rect 34146 34688 34152 34700
rect 34204 34688 34210 34740
rect 33778 34620 33784 34672
rect 33836 34660 33842 34672
rect 34793 34663 34851 34669
rect 34793 34660 34805 34663
rect 33836 34632 34805 34660
rect 33836 34620 33842 34632
rect 34793 34629 34805 34632
rect 34839 34629 34851 34663
rect 34793 34623 34851 34629
rect 31849 34595 31907 34601
rect 31849 34592 31861 34595
rect 31220 34564 31861 34592
rect 31220 34536 31248 34564
rect 31849 34561 31861 34564
rect 31895 34561 31907 34595
rect 31849 34555 31907 34561
rect 1394 34524 1400 34536
rect 1355 34496 1400 34524
rect 1394 34484 1400 34496
rect 1452 34484 1458 34536
rect 17862 34524 17868 34536
rect 17823 34496 17868 34524
rect 17862 34484 17868 34496
rect 17920 34484 17926 34536
rect 20714 34484 20720 34536
rect 20772 34524 20778 34536
rect 22741 34527 22799 34533
rect 22741 34524 22753 34527
rect 20772 34496 22753 34524
rect 20772 34484 20778 34496
rect 22741 34493 22753 34496
rect 22787 34493 22799 34527
rect 31018 34524 31024 34536
rect 30979 34496 31024 34524
rect 22741 34487 22799 34493
rect 31018 34484 31024 34496
rect 31076 34484 31082 34536
rect 31202 34524 31208 34536
rect 31163 34496 31208 34524
rect 31202 34484 31208 34496
rect 31260 34484 31266 34536
rect 31294 34484 31300 34536
rect 31352 34524 31358 34536
rect 31352 34496 31397 34524
rect 31352 34484 31358 34496
rect 31754 34484 31760 34536
rect 31812 34524 31818 34536
rect 33229 34527 33287 34533
rect 31812 34496 31857 34524
rect 31812 34484 31818 34496
rect 33229 34493 33241 34527
rect 33275 34493 33287 34527
rect 33229 34487 33287 34493
rect 30834 34388 30840 34400
rect 30795 34360 30840 34388
rect 30834 34348 30840 34360
rect 30892 34348 30898 34400
rect 33042 34388 33048 34400
rect 33003 34360 33048 34388
rect 33042 34348 33048 34360
rect 33100 34348 33106 34400
rect 33244 34388 33272 34487
rect 33318 34484 33324 34536
rect 33376 34524 33382 34536
rect 33597 34527 33655 34533
rect 33376 34496 33421 34524
rect 33376 34484 33382 34496
rect 33597 34493 33609 34527
rect 33643 34524 33655 34527
rect 33796 34524 33824 34620
rect 33870 34552 33876 34604
rect 33928 34592 33934 34604
rect 56137 34595 56195 34601
rect 33928 34564 34744 34592
rect 33928 34552 33934 34564
rect 34054 34524 34060 34536
rect 33643 34496 33824 34524
rect 34015 34496 34060 34524
rect 33643 34493 33655 34496
rect 33597 34487 33655 34493
rect 34054 34484 34060 34496
rect 34112 34484 34118 34536
rect 34716 34533 34744 34564
rect 56137 34561 56149 34595
rect 56183 34592 56195 34595
rect 57514 34592 57520 34604
rect 56183 34564 57520 34592
rect 56183 34561 56195 34564
rect 56137 34555 56195 34561
rect 57514 34552 57520 34564
rect 57572 34552 57578 34604
rect 34241 34527 34299 34533
rect 34241 34493 34253 34527
rect 34287 34493 34299 34527
rect 34241 34487 34299 34493
rect 34701 34527 34759 34533
rect 34701 34493 34713 34527
rect 34747 34493 34759 34527
rect 55306 34524 55312 34536
rect 55267 34496 55312 34524
rect 34701 34487 34759 34493
rect 33336 34456 33364 34484
rect 34250 34456 34278 34487
rect 55306 34484 55312 34496
rect 55364 34484 55370 34536
rect 56781 34527 56839 34533
rect 56781 34493 56793 34527
rect 56827 34524 56839 34527
rect 57330 34524 57336 34536
rect 56827 34496 57336 34524
rect 56827 34493 56839 34496
rect 56781 34487 56839 34493
rect 57330 34484 57336 34496
rect 57388 34484 57394 34536
rect 57422 34484 57428 34536
rect 57480 34524 57486 34536
rect 57480 34496 57573 34524
rect 57480 34484 57486 34496
rect 57882 34484 57888 34536
rect 57940 34524 57946 34536
rect 58161 34527 58219 34533
rect 58161 34524 58173 34527
rect 57940 34496 58173 34524
rect 57940 34484 57946 34496
rect 58161 34493 58173 34496
rect 58207 34493 58219 34527
rect 58161 34487 58219 34493
rect 33336 34428 34278 34456
rect 57054 34416 57060 34468
rect 57112 34456 57118 34468
rect 57440 34456 57468 34484
rect 57974 34456 57980 34468
rect 57112 34428 57468 34456
rect 57935 34428 57980 34456
rect 57112 34416 57118 34428
rect 57974 34416 57980 34428
rect 58032 34416 58038 34468
rect 33870 34388 33876 34400
rect 33244 34360 33876 34388
rect 33870 34348 33876 34360
rect 33928 34348 33934 34400
rect 34149 34391 34207 34397
rect 34149 34357 34161 34391
rect 34195 34388 34207 34391
rect 34238 34388 34244 34400
rect 34195 34360 34244 34388
rect 34195 34357 34207 34360
rect 34149 34351 34207 34357
rect 34238 34348 34244 34360
rect 34296 34348 34302 34400
rect 57238 34388 57244 34400
rect 57199 34360 57244 34388
rect 57238 34348 57244 34360
rect 57296 34348 57302 34400
rect 1104 34298 58880 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 58880 34298
rect 1104 34224 58880 34246
rect 22373 34187 22431 34193
rect 22373 34153 22385 34187
rect 22419 34153 22431 34187
rect 22373 34147 22431 34153
rect 20622 34008 20628 34060
rect 20680 34048 20686 34060
rect 21249 34051 21307 34057
rect 21249 34048 21261 34051
rect 20680 34020 21261 34048
rect 20680 34008 20686 34020
rect 21249 34017 21261 34020
rect 21295 34017 21307 34051
rect 22388 34048 22416 34147
rect 31294 34144 31300 34196
rect 31352 34184 31358 34196
rect 31849 34187 31907 34193
rect 31849 34184 31861 34187
rect 31352 34156 31861 34184
rect 31352 34144 31358 34156
rect 31849 34153 31861 34156
rect 31895 34153 31907 34187
rect 31849 34147 31907 34153
rect 33689 34187 33747 34193
rect 33689 34153 33701 34187
rect 33735 34184 33747 34187
rect 33870 34184 33876 34196
rect 33735 34156 33876 34184
rect 33735 34153 33747 34156
rect 33689 34147 33747 34153
rect 33870 34144 33876 34156
rect 33928 34144 33934 34196
rect 57974 34144 57980 34196
rect 58032 34184 58038 34196
rect 58161 34187 58219 34193
rect 58161 34184 58173 34187
rect 58032 34156 58173 34184
rect 58032 34144 58038 34156
rect 58161 34153 58173 34156
rect 58207 34153 58219 34187
rect 58161 34147 58219 34153
rect 30736 34119 30794 34125
rect 30736 34085 30748 34119
rect 30782 34116 30794 34119
rect 30834 34116 30840 34128
rect 30782 34088 30840 34116
rect 30782 34085 30794 34088
rect 30736 34079 30794 34085
rect 30834 34076 30840 34088
rect 30892 34076 30898 34128
rect 32576 34119 32634 34125
rect 32576 34085 32588 34119
rect 32622 34116 32634 34119
rect 33042 34116 33048 34128
rect 32622 34088 33048 34116
rect 32622 34085 32634 34088
rect 32576 34079 32634 34085
rect 33042 34076 33048 34088
rect 33100 34076 33106 34128
rect 33318 34076 33324 34128
rect 33376 34116 33382 34128
rect 34241 34119 34299 34125
rect 34241 34116 34253 34119
rect 33376 34088 34253 34116
rect 33376 34076 33382 34088
rect 34241 34085 34253 34088
rect 34287 34085 34299 34119
rect 34241 34079 34299 34085
rect 22646 34048 22652 34060
rect 22388 34020 22652 34048
rect 21249 34011 21307 34017
rect 22646 34008 22652 34020
rect 22704 34048 22710 34060
rect 23017 34051 23075 34057
rect 23017 34048 23029 34051
rect 22704 34020 23029 34048
rect 22704 34008 22710 34020
rect 23017 34017 23029 34020
rect 23063 34017 23075 34051
rect 23382 34048 23388 34060
rect 23343 34020 23388 34048
rect 23017 34011 23075 34017
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 25682 34008 25688 34060
rect 25740 34048 25746 34060
rect 25740 34020 34100 34048
rect 25740 34008 25746 34020
rect 19886 33940 19892 33992
rect 19944 33980 19950 33992
rect 20993 33983 21051 33989
rect 20993 33980 21005 33983
rect 19944 33952 21005 33980
rect 19944 33940 19950 33952
rect 20993 33949 21005 33952
rect 21039 33949 21051 33983
rect 23106 33980 23112 33992
rect 23067 33952 23112 33980
rect 20993 33943 21051 33949
rect 21008 33844 21036 33943
rect 23106 33940 23112 33952
rect 23164 33940 23170 33992
rect 30466 33980 30472 33992
rect 30427 33952 30472 33980
rect 30466 33940 30472 33952
rect 30524 33940 30530 33992
rect 32309 33983 32367 33989
rect 32309 33980 32321 33983
rect 31726 33952 32321 33980
rect 22922 33872 22928 33924
rect 22980 33912 22986 33924
rect 23017 33915 23075 33921
rect 23017 33912 23029 33915
rect 22980 33884 23029 33912
rect 22980 33872 22986 33884
rect 23017 33881 23029 33884
rect 23063 33881 23075 33915
rect 23017 33875 23075 33881
rect 23658 33844 23664 33856
rect 21008 33816 23664 33844
rect 23658 33804 23664 33816
rect 23716 33804 23722 33856
rect 30484 33844 30512 33940
rect 31726 33844 31754 33952
rect 32309 33949 32321 33952
rect 32355 33949 32367 33983
rect 34072 33980 34100 34020
rect 34146 34008 34152 34060
rect 34204 34048 34210 34060
rect 34204 34020 34249 34048
rect 34204 34008 34210 34020
rect 35342 34008 35348 34060
rect 35400 34048 35406 34060
rect 35713 34051 35771 34057
rect 35713 34048 35725 34051
rect 35400 34020 35725 34048
rect 35400 34008 35406 34020
rect 35713 34017 35725 34020
rect 35759 34017 35771 34051
rect 54110 34048 54116 34060
rect 35713 34011 35771 34017
rect 41386 34020 54116 34048
rect 41386 33980 41414 34020
rect 54110 34008 54116 34020
rect 54168 34008 54174 34060
rect 54941 34051 54999 34057
rect 54941 34017 54953 34051
rect 54987 34048 54999 34051
rect 55214 34048 55220 34060
rect 54987 34020 55220 34048
rect 54987 34017 54999 34020
rect 54941 34011 54999 34017
rect 55214 34008 55220 34020
rect 55272 34008 55278 34060
rect 55769 34051 55827 34057
rect 55769 34017 55781 34051
rect 55815 34048 55827 34051
rect 55858 34048 55864 34060
rect 55815 34020 55864 34048
rect 55815 34017 55827 34020
rect 55769 34011 55827 34017
rect 55858 34008 55864 34020
rect 55916 34008 55922 34060
rect 57054 34048 57060 34060
rect 57015 34020 57060 34048
rect 57054 34008 57060 34020
rect 57112 34008 57118 34060
rect 57514 34048 57520 34060
rect 57475 34020 57520 34048
rect 57514 34008 57520 34020
rect 57572 34008 57578 34060
rect 34072 33952 41414 33980
rect 57701 33983 57759 33989
rect 32309 33943 32367 33949
rect 57701 33949 57713 33983
rect 57747 33949 57759 33983
rect 57701 33943 57759 33949
rect 56873 33915 56931 33921
rect 56873 33881 56885 33915
rect 56919 33912 56931 33915
rect 57716 33912 57744 33943
rect 56919 33884 57744 33912
rect 56919 33881 56931 33884
rect 56873 33875 56931 33881
rect 30484 33816 31754 33844
rect 35805 33847 35863 33853
rect 35805 33813 35817 33847
rect 35851 33844 35863 33847
rect 35894 33844 35900 33856
rect 35851 33816 35900 33844
rect 35851 33813 35863 33816
rect 35805 33807 35863 33813
rect 35894 33804 35900 33816
rect 35952 33804 35958 33856
rect 55585 33847 55643 33853
rect 55585 33813 55597 33847
rect 55631 33844 55643 33847
rect 55766 33844 55772 33856
rect 55631 33816 55772 33844
rect 55631 33813 55643 33816
rect 55585 33807 55643 33813
rect 55766 33804 55772 33816
rect 55824 33804 55830 33856
rect 1104 33754 58880 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 58880 33754
rect 1104 33680 58880 33702
rect 20622 33640 20628 33652
rect 20583 33612 20628 33640
rect 20622 33600 20628 33612
rect 20680 33600 20686 33652
rect 22186 33600 22192 33652
rect 22244 33640 22250 33652
rect 22741 33643 22799 33649
rect 22741 33640 22753 33643
rect 22244 33612 22753 33640
rect 22244 33600 22250 33612
rect 22741 33609 22753 33612
rect 22787 33640 22799 33643
rect 54110 33640 54116 33652
rect 22787 33612 25820 33640
rect 22787 33609 22799 33612
rect 22741 33603 22799 33609
rect 1394 33436 1400 33448
rect 1355 33408 1400 33436
rect 1394 33396 1400 33408
rect 1452 33396 1458 33448
rect 20622 33436 20628 33448
rect 20583 33408 20628 33436
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 20809 33439 20867 33445
rect 20809 33405 20821 33439
rect 20855 33405 20867 33439
rect 20809 33399 20867 33405
rect 21269 33439 21327 33445
rect 21269 33405 21281 33439
rect 21315 33436 21327 33439
rect 22094 33436 22100 33448
rect 21315 33408 22100 33436
rect 21315 33405 21327 33408
rect 21269 33399 21327 33405
rect 20824 33368 20852 33399
rect 22094 33396 22100 33408
rect 22152 33396 22158 33448
rect 22646 33436 22652 33448
rect 22607 33408 22652 33436
rect 22646 33396 22652 33408
rect 22704 33396 22710 33448
rect 23477 33439 23535 33445
rect 23477 33405 23489 33439
rect 23523 33436 23535 33439
rect 23523 33408 23704 33436
rect 23523 33405 23535 33408
rect 23477 33399 23535 33405
rect 20824 33340 21404 33368
rect 21376 33312 21404 33340
rect 23676 33312 23704 33408
rect 24946 33396 24952 33448
rect 25004 33436 25010 33448
rect 25792 33445 25820 33612
rect 26068 33612 45554 33640
rect 54071 33612 54116 33640
rect 26068 33513 26096 33612
rect 31018 33532 31024 33584
rect 31076 33572 31082 33584
rect 31297 33575 31355 33581
rect 31297 33572 31309 33575
rect 31076 33544 31309 33572
rect 31076 33532 31082 33544
rect 31297 33541 31309 33544
rect 31343 33572 31355 33575
rect 31846 33572 31852 33584
rect 31343 33544 31852 33572
rect 31343 33541 31355 33544
rect 31297 33535 31355 33541
rect 31846 33532 31852 33544
rect 31904 33532 31910 33584
rect 32950 33532 32956 33584
rect 33008 33572 33014 33584
rect 33045 33575 33103 33581
rect 33045 33572 33057 33575
rect 33008 33544 33057 33572
rect 33008 33532 33014 33544
rect 33045 33541 33057 33544
rect 33091 33541 33103 33575
rect 35342 33572 35348 33584
rect 35303 33544 35348 33572
rect 33045 33535 33103 33541
rect 35342 33532 35348 33544
rect 35400 33532 35406 33584
rect 26053 33507 26111 33513
rect 26053 33473 26065 33507
rect 26099 33473 26111 33507
rect 26053 33467 26111 33473
rect 25317 33439 25375 33445
rect 25317 33436 25329 33439
rect 25004 33408 25329 33436
rect 25004 33396 25010 33408
rect 25317 33405 25329 33408
rect 25363 33405 25375 33439
rect 25317 33399 25375 33405
rect 25777 33439 25835 33445
rect 25777 33405 25789 33439
rect 25823 33405 25835 33439
rect 31202 33436 31208 33448
rect 31163 33408 31208 33436
rect 25777 33399 25835 33405
rect 31202 33396 31208 33408
rect 31260 33396 31266 33448
rect 31294 33396 31300 33448
rect 31352 33436 31358 33448
rect 31389 33439 31447 33445
rect 31389 33436 31401 33439
rect 31352 33408 31401 33436
rect 31352 33396 31358 33408
rect 31389 33405 31401 33408
rect 31435 33405 31447 33439
rect 31389 33399 31447 33405
rect 32858 33396 32864 33448
rect 32916 33436 32922 33448
rect 33045 33439 33103 33445
rect 33045 33436 33057 33439
rect 32916 33408 33057 33436
rect 32916 33396 32922 33408
rect 33045 33405 33057 33408
rect 33091 33405 33103 33439
rect 33226 33436 33232 33448
rect 33187 33408 33232 33436
rect 33045 33399 33103 33405
rect 33226 33396 33232 33408
rect 33284 33396 33290 33448
rect 33870 33396 33876 33448
rect 33928 33436 33934 33448
rect 34238 33445 34244 33448
rect 33965 33439 34023 33445
rect 33965 33436 33977 33439
rect 33928 33408 33977 33436
rect 33928 33396 33934 33408
rect 33965 33405 33977 33408
rect 34011 33405 34023 33439
rect 34232 33436 34244 33445
rect 34199 33408 34244 33436
rect 33965 33399 34023 33405
rect 34232 33399 34244 33408
rect 34238 33396 34244 33399
rect 34296 33396 34302 33448
rect 35805 33439 35863 33445
rect 35805 33405 35817 33439
rect 35851 33436 35863 33439
rect 35894 33436 35900 33448
rect 35851 33408 35900 33436
rect 35851 33405 35863 33408
rect 35805 33399 35863 33405
rect 35894 33396 35900 33408
rect 35952 33396 35958 33448
rect 35989 33439 36047 33445
rect 35989 33405 36001 33439
rect 36035 33436 36047 33439
rect 36170 33436 36176 33448
rect 36035 33408 36176 33436
rect 36035 33405 36047 33408
rect 35989 33399 36047 33405
rect 36170 33396 36176 33408
rect 36228 33396 36234 33448
rect 23744 33371 23802 33377
rect 23744 33337 23756 33371
rect 23790 33368 23802 33371
rect 23934 33368 23940 33380
rect 23790 33340 23940 33368
rect 23790 33337 23802 33340
rect 23744 33331 23802 33337
rect 23934 33328 23940 33340
rect 23992 33328 23998 33380
rect 34054 33328 34060 33380
rect 34112 33368 34118 33380
rect 35710 33368 35716 33380
rect 34112 33340 35716 33368
rect 34112 33328 34118 33340
rect 35710 33328 35716 33340
rect 35768 33328 35774 33380
rect 21358 33300 21364 33312
rect 21319 33272 21364 33300
rect 21358 33260 21364 33272
rect 21416 33260 21422 33312
rect 23658 33260 23664 33312
rect 23716 33260 23722 33312
rect 24854 33300 24860 33312
rect 24767 33272 24860 33300
rect 24854 33260 24860 33272
rect 24912 33300 24918 33312
rect 26142 33300 26148 33312
rect 24912 33272 26148 33300
rect 24912 33260 24918 33272
rect 26142 33260 26148 33272
rect 26200 33260 26206 33312
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 36173 33303 36231 33309
rect 36173 33300 36185 33303
rect 34572 33272 36185 33300
rect 34572 33260 34578 33272
rect 36173 33269 36185 33272
rect 36219 33269 36231 33303
rect 45526 33300 45554 33612
rect 54110 33600 54116 33612
rect 54168 33600 54174 33652
rect 56962 33600 56968 33652
rect 57020 33640 57026 33652
rect 57698 33640 57704 33652
rect 57020 33612 57704 33640
rect 57020 33600 57026 33612
rect 57698 33600 57704 33612
rect 57756 33600 57762 33652
rect 54128 33504 54156 33600
rect 56778 33532 56784 33584
rect 56836 33572 56842 33584
rect 57606 33572 57612 33584
rect 56836 33544 57612 33572
rect 56836 33532 56842 33544
rect 57606 33532 57612 33544
rect 57664 33532 57670 33584
rect 54389 33507 54447 33513
rect 54389 33504 54401 33507
rect 54128 33476 54401 33504
rect 54389 33473 54401 33476
rect 54435 33473 54447 33507
rect 55030 33504 55036 33516
rect 54991 33476 55036 33504
rect 54389 33467 54447 33473
rect 55030 33464 55036 33476
rect 55088 33464 55094 33516
rect 57054 33504 57060 33516
rect 57015 33476 57060 33504
rect 57054 33464 57060 33476
rect 57112 33464 57118 33516
rect 57238 33464 57244 33516
rect 57296 33504 57302 33516
rect 57701 33507 57759 33513
rect 57701 33504 57713 33507
rect 57296 33476 57713 33504
rect 57296 33464 57302 33476
rect 57701 33473 57713 33476
rect 57747 33473 57759 33507
rect 57701 33467 57759 33473
rect 56321 33439 56379 33445
rect 56321 33405 56333 33439
rect 56367 33436 56379 33439
rect 56367 33408 57284 33436
rect 56367 33405 56379 33408
rect 56321 33399 56379 33405
rect 54478 33368 54484 33380
rect 54439 33340 54484 33368
rect 54478 33328 54484 33340
rect 54536 33328 54542 33380
rect 55677 33371 55735 33377
rect 55677 33337 55689 33371
rect 55723 33337 55735 33371
rect 55677 33331 55735 33337
rect 55692 33300 55720 33331
rect 55766 33328 55772 33380
rect 55824 33368 55830 33380
rect 55824 33340 55869 33368
rect 55824 33328 55830 33340
rect 56778 33328 56784 33380
rect 56836 33368 56842 33380
rect 56873 33371 56931 33377
rect 56873 33368 56885 33371
rect 56836 33340 56885 33368
rect 56836 33328 56842 33340
rect 56873 33337 56885 33340
rect 56919 33337 56931 33371
rect 57256 33368 57284 33408
rect 57330 33396 57336 33448
rect 57388 33436 57394 33448
rect 57517 33439 57575 33445
rect 57517 33436 57529 33439
rect 57388 33408 57529 33436
rect 57388 33396 57394 33408
rect 57517 33405 57529 33408
rect 57563 33405 57575 33439
rect 57517 33399 57575 33405
rect 58802 33368 58808 33380
rect 57256 33340 58808 33368
rect 56873 33331 56931 33337
rect 58802 33328 58808 33340
rect 58860 33328 58866 33380
rect 58158 33300 58164 33312
rect 45526 33272 55720 33300
rect 58119 33272 58164 33300
rect 36173 33263 36231 33269
rect 58158 33260 58164 33272
rect 58216 33260 58222 33312
rect 1104 33210 58880 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 50326 33210
rect 50378 33158 50390 33210
rect 50442 33158 50454 33210
rect 50506 33158 50518 33210
rect 50570 33158 58880 33210
rect 1104 33136 58880 33158
rect 21361 33099 21419 33105
rect 21361 33065 21373 33099
rect 21407 33096 21419 33099
rect 22094 33096 22100 33108
rect 21407 33068 22100 33096
rect 21407 33065 21419 33068
rect 21361 33059 21419 33065
rect 22094 33056 22100 33068
rect 22152 33096 22158 33108
rect 23382 33096 23388 33108
rect 22152 33068 22416 33096
rect 23343 33068 23388 33096
rect 22152 33056 22158 33068
rect 13722 32988 13728 33040
rect 13780 33028 13786 33040
rect 22388 33028 22416 33068
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 23934 33096 23940 33108
rect 23895 33068 23940 33096
rect 23934 33056 23940 33068
rect 23992 33056 23998 33108
rect 32950 33096 32956 33108
rect 31726 33068 32956 33096
rect 23017 33031 23075 33037
rect 13780 33000 22324 33028
rect 13780 32988 13786 33000
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 20248 32963 20306 32969
rect 20248 32929 20260 32963
rect 20294 32960 20306 32963
rect 21082 32960 21088 32972
rect 20294 32932 21088 32960
rect 20294 32929 20306 32932
rect 20248 32923 20306 32929
rect 21082 32920 21088 32932
rect 21140 32920 21146 32972
rect 21358 32920 21364 32972
rect 21416 32960 21422 32972
rect 22005 32963 22063 32969
rect 22005 32960 22017 32963
rect 21416 32932 22017 32960
rect 21416 32920 21422 32932
rect 22005 32929 22017 32932
rect 22051 32929 22063 32963
rect 22005 32923 22063 32929
rect 22097 32963 22155 32969
rect 22097 32929 22109 32963
rect 22143 32960 22155 32963
rect 22186 32960 22192 32972
rect 22143 32932 22192 32960
rect 22143 32929 22155 32932
rect 22097 32923 22155 32929
rect 22186 32920 22192 32932
rect 22244 32920 22250 32972
rect 19886 32852 19892 32904
rect 19944 32892 19950 32904
rect 19981 32895 20039 32901
rect 19981 32892 19993 32895
rect 19944 32864 19993 32892
rect 19944 32852 19950 32864
rect 19981 32861 19993 32864
rect 20027 32861 20039 32895
rect 19981 32855 20039 32861
rect 22296 32824 22324 33000
rect 22388 33000 22968 33028
rect 22388 32969 22416 33000
rect 22373 32963 22431 32969
rect 22373 32929 22385 32963
rect 22419 32929 22431 32963
rect 22830 32960 22836 32972
rect 22791 32932 22836 32960
rect 22373 32923 22431 32929
rect 22830 32920 22836 32932
rect 22888 32920 22894 32972
rect 22940 32960 22968 33000
rect 23017 32997 23029 33031
rect 23063 33028 23075 33031
rect 23566 33028 23572 33040
rect 23063 33000 23572 33028
rect 23063 32997 23075 33000
rect 23017 32991 23075 32997
rect 23566 32988 23572 33000
rect 23624 32988 23630 33040
rect 31573 33031 31631 33037
rect 31573 32997 31585 33031
rect 31619 33028 31631 33031
rect 31726 33028 31754 33068
rect 32950 33056 32956 33068
rect 33008 33056 33014 33108
rect 33321 33099 33379 33105
rect 33321 33065 33333 33099
rect 33367 33096 33379 33099
rect 35710 33096 35716 33108
rect 33367 33068 34560 33096
rect 35671 33068 35716 33096
rect 33367 33065 33379 33068
rect 33321 33059 33379 33065
rect 34057 33031 34115 33037
rect 34057 33028 34069 33031
rect 31619 33000 31754 33028
rect 32876 33000 34069 33028
rect 31619 32997 31631 33000
rect 31573 32991 31631 32997
rect 32876 32972 32904 33000
rect 34057 32997 34069 33000
rect 34103 32997 34115 33031
rect 34532 33028 34560 33068
rect 35710 33056 35716 33068
rect 35768 33056 35774 33108
rect 53653 33099 53711 33105
rect 53653 33065 53665 33099
rect 53699 33096 53711 33099
rect 55769 33099 55827 33105
rect 53699 33068 54524 33096
rect 53699 33065 53711 33068
rect 53653 33059 53711 33065
rect 34698 33028 34704 33040
rect 34532 33000 34704 33028
rect 34057 32991 34115 32997
rect 34698 32988 34704 33000
rect 34756 33028 34762 33040
rect 54496 33037 54524 33068
rect 55769 33065 55781 33099
rect 55815 33096 55827 33099
rect 55858 33096 55864 33108
rect 55815 33068 55864 33096
rect 55815 33065 55827 33068
rect 55769 33059 55827 33065
rect 55858 33056 55864 33068
rect 55916 33056 55922 33108
rect 54481 33031 54539 33037
rect 34756 33000 36124 33028
rect 34756 32988 34762 33000
rect 23106 32960 23112 32972
rect 22940 32932 23112 32960
rect 23106 32920 23112 32932
rect 23164 32920 23170 32972
rect 23201 32963 23259 32969
rect 23201 32929 23213 32963
rect 23247 32929 23259 32963
rect 23842 32960 23848 32972
rect 23803 32932 23848 32960
rect 23201 32923 23259 32929
rect 22646 32852 22652 32904
rect 22704 32892 22710 32904
rect 23216 32892 23244 32923
rect 23842 32920 23848 32932
rect 23900 32920 23906 32972
rect 24026 32960 24032 32972
rect 23987 32932 24032 32960
rect 24026 32920 24032 32932
rect 24084 32920 24090 32972
rect 24946 32920 24952 32972
rect 25004 32960 25010 32972
rect 25225 32963 25283 32969
rect 25225 32960 25237 32963
rect 25004 32932 25237 32960
rect 25004 32920 25010 32932
rect 25225 32929 25237 32932
rect 25271 32929 25283 32963
rect 25774 32960 25780 32972
rect 25735 32932 25780 32960
rect 25225 32923 25283 32929
rect 25774 32920 25780 32932
rect 25832 32920 25838 32972
rect 31754 32960 31760 32972
rect 31715 32932 31760 32960
rect 31754 32920 31760 32932
rect 31812 32920 31818 32972
rect 31846 32920 31852 32972
rect 31904 32960 31910 32972
rect 32858 32960 32864 32972
rect 31904 32932 32864 32960
rect 31904 32920 31910 32932
rect 32858 32920 32864 32932
rect 32916 32920 32922 32972
rect 33107 32963 33165 32969
rect 33107 32929 33119 32963
rect 33153 32960 33165 32963
rect 34204 32963 34262 32969
rect 33153 32932 33272 32960
rect 33153 32929 33165 32932
rect 33107 32923 33165 32929
rect 33244 32904 33272 32932
rect 34204 32929 34216 32963
rect 34250 32960 34262 32963
rect 34514 32960 34520 32972
rect 34250 32932 34520 32960
rect 34250 32929 34262 32932
rect 34204 32923 34262 32929
rect 34514 32920 34520 32932
rect 34572 32920 34578 32972
rect 35894 32960 35900 32972
rect 35855 32932 35900 32960
rect 35894 32920 35900 32932
rect 35952 32920 35958 32972
rect 36096 32969 36124 33000
rect 54481 32997 54493 33031
rect 54527 32997 54539 33031
rect 54481 32991 54539 32997
rect 54570 32988 54576 33040
rect 54628 33028 54634 33040
rect 57333 33031 57391 33037
rect 57333 33028 57345 33031
rect 54628 33000 57345 33028
rect 54628 32988 54634 33000
rect 57333 32997 57345 33000
rect 57379 32997 57391 33031
rect 57333 32991 57391 32997
rect 57885 33031 57943 33037
rect 57885 32997 57897 33031
rect 57931 33028 57943 33031
rect 58250 33028 58256 33040
rect 57931 33000 58256 33028
rect 57931 32997 57943 33000
rect 57885 32991 57943 32997
rect 58250 32988 58256 33000
rect 58308 32988 58314 33040
rect 36081 32963 36139 32969
rect 36081 32929 36093 32963
rect 36127 32929 36139 32963
rect 53834 32960 53840 32972
rect 53795 32932 53840 32960
rect 36081 32923 36139 32929
rect 53834 32920 53840 32932
rect 53892 32920 53898 32972
rect 55585 32963 55643 32969
rect 55585 32929 55597 32963
rect 55631 32960 55643 32963
rect 56226 32960 56232 32972
rect 55631 32932 56232 32960
rect 55631 32929 55643 32932
rect 55585 32923 55643 32929
rect 56226 32920 56232 32932
rect 56284 32920 56290 32972
rect 22704 32864 23244 32892
rect 25961 32895 26019 32901
rect 22704 32852 22710 32864
rect 25961 32861 25973 32895
rect 26007 32892 26019 32895
rect 31662 32892 31668 32904
rect 26007 32864 31668 32892
rect 26007 32861 26019 32864
rect 25961 32855 26019 32861
rect 31662 32852 31668 32864
rect 31720 32852 31726 32904
rect 33226 32852 33232 32904
rect 33284 32892 33290 32904
rect 34425 32895 34483 32901
rect 34425 32892 34437 32895
rect 33284 32864 34437 32892
rect 33284 32852 33290 32864
rect 34425 32861 34437 32864
rect 34471 32861 34483 32895
rect 36170 32892 36176 32904
rect 36131 32864 36176 32892
rect 34425 32855 34483 32861
rect 36170 32852 36176 32864
rect 36228 32852 36234 32904
rect 49970 32852 49976 32904
rect 50028 32892 50034 32904
rect 54389 32895 54447 32901
rect 54389 32892 54401 32895
rect 50028 32864 54401 32892
rect 50028 32852 50034 32864
rect 54389 32861 54401 32864
rect 54435 32861 54447 32895
rect 57241 32895 57299 32901
rect 57241 32892 57253 32895
rect 54389 32855 54447 32861
rect 54496 32864 57253 32892
rect 30926 32824 30932 32836
rect 22296 32796 30932 32824
rect 30926 32784 30932 32796
rect 30984 32784 30990 32836
rect 32953 32827 33011 32833
rect 32953 32793 32965 32827
rect 32999 32824 33011 32827
rect 34054 32824 34060 32836
rect 32999 32796 34060 32824
rect 32999 32793 33011 32796
rect 32953 32787 33011 32793
rect 34054 32784 34060 32796
rect 34112 32824 34118 32836
rect 34333 32827 34391 32833
rect 34333 32824 34345 32827
rect 34112 32796 34345 32824
rect 34112 32784 34118 32796
rect 34333 32793 34345 32796
rect 34379 32793 34391 32827
rect 34333 32787 34391 32793
rect 50338 32784 50344 32836
rect 50396 32824 50402 32836
rect 54496 32824 54524 32864
rect 57241 32861 57253 32864
rect 57287 32861 57299 32895
rect 57241 32855 57299 32861
rect 54938 32824 54944 32836
rect 50396 32796 54524 32824
rect 54899 32796 54944 32824
rect 50396 32784 50402 32796
rect 54938 32784 54944 32796
rect 54996 32784 55002 32836
rect 21634 32716 21640 32768
rect 21692 32756 21698 32768
rect 21821 32759 21879 32765
rect 21821 32756 21833 32759
rect 21692 32728 21833 32756
rect 21692 32716 21698 32728
rect 21821 32725 21833 32728
rect 21867 32725 21879 32759
rect 21821 32719 21879 32725
rect 22281 32759 22339 32765
rect 22281 32725 22293 32759
rect 22327 32756 22339 32759
rect 22646 32756 22652 32768
rect 22327 32728 22652 32756
rect 22327 32725 22339 32728
rect 22281 32719 22339 32725
rect 22646 32716 22652 32728
rect 22704 32716 22710 32768
rect 22830 32716 22836 32768
rect 22888 32756 22894 32768
rect 23290 32756 23296 32768
rect 22888 32728 23296 32756
rect 22888 32716 22894 32728
rect 23290 32716 23296 32728
rect 23348 32756 23354 32768
rect 24854 32756 24860 32768
rect 23348 32728 24860 32756
rect 23348 32716 23354 32728
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 31570 32756 31576 32768
rect 31531 32728 31576 32756
rect 31570 32716 31576 32728
rect 31628 32716 31634 32768
rect 34146 32716 34152 32768
rect 34204 32756 34210 32768
rect 34517 32759 34575 32765
rect 34517 32756 34529 32759
rect 34204 32728 34529 32756
rect 34204 32716 34210 32728
rect 34517 32725 34529 32728
rect 34563 32725 34575 32759
rect 34517 32719 34575 32725
rect 1104 32666 58880 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 58880 32666
rect 1104 32592 58880 32614
rect 20714 32512 20720 32564
rect 20772 32552 20778 32564
rect 50338 32552 50344 32564
rect 20772 32524 50344 32552
rect 20772 32512 20778 32524
rect 50338 32512 50344 32524
rect 50396 32512 50402 32564
rect 54389 32555 54447 32561
rect 54389 32521 54401 32555
rect 54435 32552 54447 32555
rect 54478 32552 54484 32564
rect 54435 32524 54484 32552
rect 54435 32521 54447 32524
rect 54389 32515 54447 32521
rect 54478 32512 54484 32524
rect 54536 32512 54542 32564
rect 17034 32444 17040 32496
rect 17092 32484 17098 32496
rect 20990 32484 20996 32496
rect 17092 32456 20996 32484
rect 17092 32444 17098 32456
rect 20990 32444 20996 32456
rect 21048 32444 21054 32496
rect 23290 32444 23296 32496
rect 23348 32444 23354 32496
rect 23477 32487 23535 32493
rect 23477 32453 23489 32487
rect 23523 32453 23535 32487
rect 23477 32447 23535 32453
rect 13722 32416 13728 32428
rect 13683 32388 13728 32416
rect 13722 32376 13728 32388
rect 13780 32376 13786 32428
rect 14918 32416 14924 32428
rect 14660 32388 14924 32416
rect 13354 32348 13360 32360
rect 13315 32320 13360 32348
rect 13354 32308 13360 32320
rect 13412 32348 13418 32360
rect 13814 32348 13820 32360
rect 13412 32320 13820 32348
rect 13412 32308 13418 32320
rect 13814 32308 13820 32320
rect 13872 32308 13878 32360
rect 14660 32357 14688 32388
rect 14918 32376 14924 32388
rect 14976 32416 14982 32428
rect 14976 32388 15608 32416
rect 14976 32376 14982 32388
rect 15580 32360 15608 32388
rect 14645 32351 14703 32357
rect 14645 32317 14657 32351
rect 14691 32317 14703 32351
rect 14645 32311 14703 32317
rect 14829 32351 14887 32357
rect 14829 32317 14841 32351
rect 14875 32348 14887 32351
rect 15378 32348 15384 32360
rect 14875 32320 15384 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 15378 32308 15384 32320
rect 15436 32308 15442 32360
rect 15473 32351 15531 32357
rect 15473 32317 15485 32351
rect 15519 32317 15531 32351
rect 15473 32311 15531 32317
rect 13170 32280 13176 32292
rect 13131 32252 13176 32280
rect 13170 32240 13176 32252
rect 13228 32240 13234 32292
rect 13906 32240 13912 32292
rect 13964 32280 13970 32292
rect 15488 32280 15516 32311
rect 15562 32308 15568 32360
rect 15620 32348 15626 32360
rect 17957 32351 18015 32357
rect 17957 32348 17969 32351
rect 15620 32320 17969 32348
rect 15620 32308 15626 32320
rect 17957 32317 17969 32320
rect 18003 32317 18015 32351
rect 17957 32311 18015 32317
rect 18141 32351 18199 32357
rect 18141 32317 18153 32351
rect 18187 32348 18199 32351
rect 18874 32348 18880 32360
rect 18187 32320 18880 32348
rect 18187 32317 18199 32320
rect 18141 32311 18199 32317
rect 18874 32308 18880 32320
rect 18932 32308 18938 32360
rect 19426 32348 19432 32360
rect 19387 32320 19432 32348
rect 19426 32308 19432 32320
rect 19484 32308 19490 32360
rect 20622 32308 20628 32360
rect 20680 32348 20686 32360
rect 20797 32351 20855 32357
rect 20797 32348 20809 32351
rect 20680 32320 20809 32348
rect 20680 32308 20686 32320
rect 13964 32252 15516 32280
rect 20732 32280 20760 32320
rect 20797 32317 20809 32320
rect 20843 32317 20855 32351
rect 20990 32348 20996 32360
rect 20951 32320 20996 32348
rect 20797 32311 20855 32317
rect 20990 32308 20996 32320
rect 21048 32308 21054 32360
rect 21450 32348 21456 32360
rect 21411 32320 21456 32348
rect 21450 32308 21456 32320
rect 21508 32308 21514 32360
rect 22830 32308 22836 32360
rect 22888 32348 22894 32360
rect 23308 32357 23336 32444
rect 23492 32360 23520 32447
rect 31754 32444 31760 32496
rect 31812 32484 31818 32496
rect 33137 32487 33195 32493
rect 33137 32484 33149 32487
rect 31812 32456 33149 32484
rect 31812 32444 31818 32456
rect 33137 32453 33149 32456
rect 33183 32484 33195 32487
rect 33226 32484 33232 32496
rect 33183 32456 33232 32484
rect 33183 32453 33195 32456
rect 33137 32447 33195 32453
rect 33226 32444 33232 32456
rect 33284 32444 33290 32496
rect 55490 32444 55496 32496
rect 55548 32484 55554 32496
rect 55953 32487 56011 32493
rect 55953 32484 55965 32487
rect 55548 32456 55965 32484
rect 55548 32444 55554 32456
rect 55953 32453 55965 32456
rect 55999 32484 56011 32487
rect 58161 32487 58219 32493
rect 55999 32456 56272 32484
rect 55999 32453 56011 32456
rect 55953 32447 56011 32453
rect 25682 32416 25688 32428
rect 25643 32388 25688 32416
rect 25682 32376 25688 32388
rect 25740 32376 25746 32428
rect 30466 32376 30472 32428
rect 30524 32416 30530 32428
rect 30561 32419 30619 32425
rect 30561 32416 30573 32419
rect 30524 32388 30573 32416
rect 30524 32376 30530 32388
rect 30561 32385 30573 32388
rect 30607 32385 30619 32419
rect 30561 32379 30619 32385
rect 31662 32376 31668 32428
rect 31720 32416 31726 32428
rect 31720 32388 34008 32416
rect 31720 32376 31726 32388
rect 22925 32351 22983 32357
rect 22925 32348 22937 32351
rect 22888 32320 22937 32348
rect 22888 32308 22894 32320
rect 22925 32317 22937 32320
rect 22971 32317 22983 32351
rect 22925 32311 22983 32317
rect 23293 32351 23351 32357
rect 23293 32317 23305 32351
rect 23339 32317 23351 32351
rect 23293 32311 23351 32317
rect 22554 32280 22560 32292
rect 20732 32252 22560 32280
rect 13964 32240 13970 32252
rect 22554 32240 22560 32252
rect 22612 32240 22618 32292
rect 14734 32212 14740 32224
rect 14695 32184 14740 32212
rect 14734 32172 14740 32184
rect 14792 32172 14798 32224
rect 15289 32215 15347 32221
rect 15289 32181 15301 32215
rect 15335 32212 15347 32215
rect 16022 32212 16028 32224
rect 15335 32184 16028 32212
rect 15335 32181 15347 32184
rect 15289 32175 15347 32181
rect 16022 32172 16028 32184
rect 16080 32172 16086 32224
rect 17954 32172 17960 32224
rect 18012 32212 18018 32224
rect 18049 32215 18107 32221
rect 18049 32212 18061 32215
rect 18012 32184 18061 32212
rect 18012 32172 18018 32184
rect 18049 32181 18061 32184
rect 18095 32181 18107 32215
rect 18049 32175 18107 32181
rect 19334 32172 19340 32224
rect 19392 32212 19398 32224
rect 19521 32215 19579 32221
rect 19521 32212 19533 32215
rect 19392 32184 19533 32212
rect 19392 32172 19398 32184
rect 19521 32181 19533 32184
rect 19567 32212 19579 32215
rect 20438 32212 20444 32224
rect 19567 32184 20444 32212
rect 19567 32181 19579 32184
rect 19521 32175 19579 32181
rect 20438 32172 20444 32184
rect 20496 32172 20502 32224
rect 20898 32212 20904 32224
rect 20859 32184 20904 32212
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21174 32172 21180 32224
rect 21232 32212 21238 32224
rect 21545 32215 21603 32221
rect 21545 32212 21557 32215
rect 21232 32184 21557 32212
rect 21232 32172 21238 32184
rect 21545 32181 21557 32184
rect 21591 32181 21603 32215
rect 22940 32212 22968 32311
rect 23474 32308 23480 32360
rect 23532 32308 23538 32360
rect 23934 32348 23940 32360
rect 23895 32320 23940 32348
rect 23934 32308 23940 32320
rect 23992 32308 23998 32360
rect 24946 32348 24952 32360
rect 24907 32320 24952 32348
rect 24946 32308 24952 32320
rect 25004 32308 25010 32360
rect 25406 32348 25412 32360
rect 25367 32320 25412 32348
rect 25406 32308 25412 32320
rect 25464 32308 25470 32360
rect 26142 32348 26148 32360
rect 26103 32320 26148 32348
rect 26142 32308 26148 32320
rect 26200 32308 26206 32360
rect 30828 32351 30886 32357
rect 30828 32317 30840 32351
rect 30874 32348 30886 32351
rect 31570 32348 31576 32360
rect 30874 32320 31576 32348
rect 30874 32317 30886 32320
rect 30828 32311 30886 32317
rect 31570 32308 31576 32320
rect 31628 32308 31634 32360
rect 33045 32351 33103 32357
rect 33045 32348 33057 32351
rect 31956 32320 33057 32348
rect 23106 32280 23112 32292
rect 23067 32252 23112 32280
rect 23106 32240 23112 32252
rect 23164 32240 23170 32292
rect 23201 32283 23259 32289
rect 23201 32249 23213 32283
rect 23247 32280 23259 32283
rect 23566 32280 23572 32292
rect 23247 32252 23572 32280
rect 23247 32249 23259 32252
rect 23201 32243 23259 32249
rect 23566 32240 23572 32252
rect 23624 32280 23630 32292
rect 23952 32280 23980 32308
rect 23624 32252 23980 32280
rect 23624 32240 23630 32252
rect 24026 32240 24032 32292
rect 24084 32280 24090 32292
rect 24084 32252 24129 32280
rect 24084 32240 24090 32252
rect 25774 32212 25780 32224
rect 22940 32184 25780 32212
rect 21545 32175 21603 32181
rect 25774 32172 25780 32184
rect 25832 32212 25838 32224
rect 31956 32221 31984 32320
rect 33045 32317 33057 32320
rect 33091 32317 33103 32351
rect 33870 32348 33876 32360
rect 33831 32320 33876 32348
rect 33045 32311 33103 32317
rect 33870 32308 33876 32320
rect 33928 32308 33934 32360
rect 33980 32348 34008 32388
rect 53834 32376 53840 32428
rect 53892 32416 53898 32428
rect 55858 32416 55864 32428
rect 53892 32388 55864 32416
rect 53892 32376 53898 32388
rect 54588 32357 54616 32388
rect 55858 32376 55864 32388
rect 55916 32376 55922 32428
rect 56244 32425 56272 32456
rect 58161 32453 58173 32487
rect 58207 32484 58219 32487
rect 58526 32484 58532 32496
rect 58207 32456 58532 32484
rect 58207 32453 58219 32456
rect 58161 32447 58219 32453
rect 58526 32444 58532 32456
rect 58584 32444 58590 32496
rect 56229 32419 56287 32425
rect 56229 32385 56241 32419
rect 56275 32385 56287 32419
rect 57146 32416 57152 32428
rect 57107 32388 57152 32416
rect 56229 32379 56287 32385
rect 57146 32376 57152 32388
rect 57204 32376 57210 32428
rect 54573 32351 54631 32357
rect 33980 32320 41414 32348
rect 34140 32283 34198 32289
rect 34140 32249 34152 32283
rect 34186 32280 34198 32283
rect 34238 32280 34244 32292
rect 34186 32252 34244 32280
rect 34186 32249 34198 32252
rect 34140 32243 34198 32249
rect 34238 32240 34244 32252
rect 34296 32240 34302 32292
rect 41386 32280 41414 32320
rect 54573 32317 54585 32351
rect 54619 32317 54631 32351
rect 54573 32311 54631 32317
rect 54662 32308 54668 32360
rect 54720 32348 54726 32360
rect 55030 32348 55036 32360
rect 54720 32320 55036 32348
rect 54720 32308 54726 32320
rect 55030 32308 55036 32320
rect 55088 32348 55094 32360
rect 55493 32351 55551 32357
rect 55493 32348 55505 32351
rect 55088 32320 55505 32348
rect 55088 32308 55094 32320
rect 55493 32317 55505 32320
rect 55539 32317 55551 32351
rect 55493 32311 55551 32317
rect 57977 32351 58035 32357
rect 57977 32317 57989 32351
rect 58023 32348 58035 32351
rect 58158 32348 58164 32360
rect 58023 32320 58164 32348
rect 58023 32317 58035 32320
rect 57977 32311 58035 32317
rect 58158 32308 58164 32320
rect 58216 32308 58222 32360
rect 49970 32280 49976 32292
rect 41386 32252 49976 32280
rect 49970 32240 49976 32252
rect 50028 32240 50034 32292
rect 56321 32283 56379 32289
rect 55692 32252 56180 32280
rect 26237 32215 26295 32221
rect 26237 32212 26249 32215
rect 25832 32184 26249 32212
rect 25832 32172 25838 32184
rect 26237 32181 26249 32184
rect 26283 32181 26295 32215
rect 26237 32175 26295 32181
rect 31941 32215 31999 32221
rect 31941 32181 31953 32215
rect 31987 32181 31999 32215
rect 31941 32175 31999 32181
rect 34422 32172 34428 32224
rect 34480 32212 34486 32224
rect 35253 32215 35311 32221
rect 35253 32212 35265 32215
rect 34480 32184 35265 32212
rect 34480 32172 34486 32184
rect 35253 32181 35265 32184
rect 35299 32212 35311 32215
rect 35710 32212 35716 32224
rect 35299 32184 35716 32212
rect 35299 32181 35311 32184
rect 35253 32175 35311 32181
rect 35710 32172 35716 32184
rect 35768 32172 35774 32224
rect 55692 32221 55720 32252
rect 55677 32215 55735 32221
rect 55677 32181 55689 32215
rect 55723 32181 55735 32215
rect 56152 32212 56180 32252
rect 56321 32249 56333 32283
rect 56367 32249 56379 32283
rect 56321 32243 56379 32249
rect 56336 32212 56364 32243
rect 56152 32184 56364 32212
rect 55677 32175 55735 32181
rect 1104 32122 58880 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 50326 32122
rect 50378 32070 50390 32122
rect 50442 32070 50454 32122
rect 50506 32070 50518 32122
rect 50570 32070 58880 32122
rect 1104 32048 58880 32070
rect 16850 32008 16856 32020
rect 16763 31980 16856 32008
rect 16850 31968 16856 31980
rect 16908 32008 16914 32020
rect 17862 32008 17868 32020
rect 16908 31980 17868 32008
rect 16908 31968 16914 31980
rect 17862 31968 17868 31980
rect 17920 31968 17926 32020
rect 19061 32011 19119 32017
rect 19061 31977 19073 32011
rect 19107 32008 19119 32011
rect 19426 32008 19432 32020
rect 19107 31980 19432 32008
rect 19107 31977 19119 31980
rect 19061 31971 19119 31977
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 21082 31968 21088 32020
rect 21140 32008 21146 32020
rect 21177 32011 21235 32017
rect 21177 32008 21189 32011
rect 21140 31980 21189 32008
rect 21140 31968 21146 31980
rect 21177 31977 21189 31980
rect 21223 31977 21235 32011
rect 24946 32008 24952 32020
rect 21177 31971 21235 31977
rect 21284 31980 24952 32008
rect 12434 31900 12440 31952
rect 12492 31940 12498 31952
rect 12492 31912 12537 31940
rect 12912 31912 13768 31940
rect 12492 31900 12498 31912
rect 1394 31872 1400 31884
rect 1355 31844 1400 31872
rect 1394 31832 1400 31844
rect 1452 31832 1458 31884
rect 12066 31832 12072 31884
rect 12124 31872 12130 31884
rect 12124 31844 12434 31872
rect 12124 31832 12130 31844
rect 12406 31804 12434 31844
rect 12912 31816 12940 31912
rect 13262 31832 13268 31884
rect 13320 31872 13326 31884
rect 13633 31875 13691 31881
rect 13633 31872 13645 31875
rect 13320 31844 13645 31872
rect 13320 31832 13326 31844
rect 13633 31841 13645 31844
rect 13679 31841 13691 31875
rect 13633 31835 13691 31841
rect 12584 31807 12642 31813
rect 12584 31804 12596 31807
rect 12406 31776 12596 31804
rect 12584 31773 12596 31776
rect 12630 31773 12642 31807
rect 12584 31767 12642 31773
rect 12805 31807 12863 31813
rect 12805 31773 12817 31807
rect 12851 31804 12863 31807
rect 12894 31804 12900 31816
rect 12851 31776 12900 31804
rect 12851 31773 12863 31776
rect 12805 31767 12863 31773
rect 12894 31764 12900 31776
rect 12952 31764 12958 31816
rect 13740 31804 13768 31912
rect 14550 31900 14556 31952
rect 14608 31940 14614 31952
rect 14608 31912 15056 31940
rect 14608 31900 14614 31912
rect 14918 31872 14924 31884
rect 14879 31844 14924 31872
rect 14918 31832 14924 31844
rect 14976 31832 14982 31884
rect 15028 31872 15056 31912
rect 15470 31900 15476 31952
rect 15528 31940 15534 31952
rect 17678 31940 17684 31952
rect 15528 31912 15792 31940
rect 15528 31900 15534 31912
rect 15105 31875 15163 31881
rect 15105 31872 15117 31875
rect 15028 31844 15117 31872
rect 15105 31841 15117 31844
rect 15151 31841 15163 31875
rect 15562 31872 15568 31884
rect 15523 31844 15568 31872
rect 15105 31835 15163 31841
rect 15562 31832 15568 31844
rect 15620 31832 15626 31884
rect 15764 31881 15792 31912
rect 16230 31912 17684 31940
rect 16230 31881 16258 31912
rect 17678 31900 17684 31912
rect 17736 31900 17742 31952
rect 17954 31949 17960 31952
rect 17948 31903 17960 31949
rect 18012 31940 18018 31952
rect 20714 31940 20720 31952
rect 18012 31912 18048 31940
rect 20675 31912 20720 31940
rect 17954 31900 17960 31903
rect 18012 31900 18018 31912
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 21284 31940 21312 31980
rect 24946 31968 24952 31980
rect 25004 31968 25010 32020
rect 32033 32011 32091 32017
rect 32033 31977 32045 32011
rect 32079 32008 32091 32011
rect 33870 32008 33876 32020
rect 32079 31980 33876 32008
rect 32079 31977 32091 31980
rect 32033 31971 32091 31977
rect 33870 31968 33876 31980
rect 33928 31968 33934 32020
rect 34238 32008 34244 32020
rect 34199 31980 34244 32008
rect 34238 31968 34244 31980
rect 34296 31968 34302 32020
rect 41386 31980 55168 32008
rect 22094 31940 22100 31952
rect 20824 31912 21312 31940
rect 21560 31912 22100 31940
rect 15749 31875 15807 31881
rect 15749 31841 15761 31875
rect 15795 31841 15807 31875
rect 15749 31835 15807 31841
rect 16209 31875 16267 31881
rect 16209 31841 16221 31875
rect 16255 31841 16267 31875
rect 16209 31835 16267 31841
rect 16393 31875 16451 31881
rect 16393 31841 16405 31875
rect 16439 31841 16451 31875
rect 17034 31872 17040 31884
rect 16995 31844 17040 31872
rect 16393 31835 16451 31841
rect 13740 31776 13860 31804
rect 13832 31745 13860 31776
rect 15010 31764 15016 31816
rect 15068 31804 15074 31816
rect 15657 31807 15715 31813
rect 15657 31804 15669 31807
rect 15068 31776 15669 31804
rect 15068 31764 15074 31776
rect 15657 31773 15669 31776
rect 15703 31773 15715 31807
rect 16298 31804 16304 31816
rect 16259 31776 16304 31804
rect 15657 31767 15715 31773
rect 16298 31764 16304 31776
rect 16356 31764 16362 31816
rect 13817 31739 13875 31745
rect 13817 31705 13829 31739
rect 13863 31736 13875 31739
rect 13863 31708 13897 31736
rect 13863 31705 13875 31708
rect 13817 31699 13875 31705
rect 13998 31696 14004 31748
rect 14056 31736 14062 31748
rect 16408 31736 16436 31835
rect 17034 31832 17040 31844
rect 17092 31832 17098 31884
rect 19978 31872 19984 31884
rect 17696 31844 19840 31872
rect 19939 31844 19984 31872
rect 17696 31813 17724 31844
rect 17681 31807 17739 31813
rect 17681 31804 17693 31807
rect 16592 31776 17693 31804
rect 16592 31736 16620 31776
rect 17681 31773 17693 31776
rect 17727 31773 17739 31807
rect 19812 31804 19840 31844
rect 19978 31832 19984 31844
rect 20036 31832 20042 31884
rect 20438 31872 20444 31884
rect 20399 31844 20444 31872
rect 20438 31832 20444 31844
rect 20496 31832 20502 31884
rect 19886 31804 19892 31816
rect 19799 31776 19892 31804
rect 17681 31767 17739 31773
rect 19886 31764 19892 31776
rect 19944 31804 19950 31816
rect 20530 31804 20536 31816
rect 19944 31776 20536 31804
rect 19944 31764 19950 31776
rect 20530 31764 20536 31776
rect 20588 31764 20594 31816
rect 20824 31804 20852 31912
rect 21082 31832 21088 31884
rect 21140 31872 21146 31884
rect 21560 31881 21588 31912
rect 22094 31900 22100 31912
rect 22152 31900 22158 31952
rect 22281 31943 22339 31949
rect 22281 31909 22293 31943
rect 22327 31940 22339 31943
rect 22738 31940 22744 31952
rect 22327 31912 22744 31940
rect 22327 31909 22339 31912
rect 22281 31903 22339 31909
rect 22738 31900 22744 31912
rect 22796 31900 22802 31952
rect 21453 31875 21511 31881
rect 21453 31872 21465 31875
rect 21140 31844 21465 31872
rect 21140 31832 21146 31844
rect 21453 31841 21465 31844
rect 21499 31841 21511 31875
rect 21453 31835 21511 31841
rect 21545 31875 21603 31881
rect 21545 31841 21557 31875
rect 21591 31841 21603 31875
rect 21545 31835 21603 31841
rect 21637 31875 21695 31881
rect 21637 31841 21649 31875
rect 21683 31841 21695 31875
rect 21818 31872 21824 31884
rect 21779 31844 21824 31872
rect 21637 31835 21695 31841
rect 20640 31776 20852 31804
rect 14056 31708 16436 31736
rect 16500 31708 16620 31736
rect 14056 31696 14062 31708
rect 12618 31628 12624 31680
rect 12676 31668 12682 31680
rect 12713 31671 12771 31677
rect 12713 31668 12725 31671
rect 12676 31640 12725 31668
rect 12676 31628 12682 31640
rect 12713 31637 12725 31640
rect 12759 31637 12771 31671
rect 12713 31631 12771 31637
rect 13081 31671 13139 31677
rect 13081 31637 13093 31671
rect 13127 31668 13139 31671
rect 13446 31668 13452 31680
rect 13127 31640 13452 31668
rect 13127 31637 13139 31640
rect 13081 31631 13139 31637
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 14918 31668 14924 31680
rect 14879 31640 14924 31668
rect 14918 31628 14924 31640
rect 14976 31628 14982 31680
rect 15102 31628 15108 31680
rect 15160 31668 15166 31680
rect 16500 31668 16528 31708
rect 19978 31696 19984 31748
rect 20036 31736 20042 31748
rect 20640 31736 20668 31776
rect 20036 31708 20668 31736
rect 20036 31696 20042 31708
rect 15160 31640 16528 31668
rect 15160 31628 15166 31640
rect 18046 31628 18052 31680
rect 18104 31668 18110 31680
rect 20806 31668 20812 31680
rect 18104 31640 20812 31668
rect 18104 31628 18110 31640
rect 20806 31628 20812 31640
rect 20864 31668 20870 31680
rect 21652 31668 21680 31835
rect 21818 31832 21824 31844
rect 21876 31832 21882 31884
rect 22462 31872 22468 31884
rect 22423 31844 22468 31872
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 22554 31832 22560 31884
rect 22612 31872 22618 31884
rect 23109 31875 23167 31881
rect 23109 31872 23121 31875
rect 22612 31844 23121 31872
rect 22612 31832 22618 31844
rect 23109 31841 23121 31844
rect 23155 31841 23167 31875
rect 23109 31835 23167 31841
rect 23293 31875 23351 31881
rect 23293 31841 23305 31875
rect 23339 31872 23351 31875
rect 23382 31872 23388 31884
rect 23339 31844 23388 31872
rect 23339 31841 23351 31844
rect 23293 31835 23351 31841
rect 22646 31804 22652 31816
rect 22607 31776 22652 31804
rect 22646 31764 22652 31776
rect 22704 31764 22710 31816
rect 23124 31804 23152 31835
rect 23382 31832 23388 31844
rect 23440 31832 23446 31884
rect 24964 31872 24992 31968
rect 25774 31900 25780 31952
rect 25832 31940 25838 31952
rect 26513 31943 26571 31949
rect 26513 31940 26525 31943
rect 25832 31912 26525 31940
rect 25832 31900 25838 31912
rect 26513 31909 26525 31912
rect 26559 31909 26571 31943
rect 41386 31940 41414 31980
rect 55140 31949 55168 31980
rect 55674 31968 55680 32020
rect 55732 31968 55738 32020
rect 56410 31968 56416 32020
rect 56468 32008 56474 32020
rect 56468 31980 57468 32008
rect 56468 31968 56474 31980
rect 26513 31903 26571 31909
rect 26896 31912 41414 31940
rect 55125 31943 55183 31949
rect 25225 31875 25283 31881
rect 25225 31872 25237 31875
rect 24964 31844 25237 31872
rect 25225 31841 25237 31844
rect 25271 31841 25283 31875
rect 25225 31835 25283 31841
rect 25685 31875 25743 31881
rect 25685 31841 25697 31875
rect 25731 31841 25743 31875
rect 25685 31835 25743 31841
rect 23842 31804 23848 31816
rect 23124 31776 23848 31804
rect 23842 31764 23848 31776
rect 23900 31764 23906 31816
rect 24762 31764 24768 31816
rect 24820 31804 24826 31816
rect 25700 31804 25728 31835
rect 26326 31832 26332 31884
rect 26384 31872 26390 31884
rect 26421 31875 26479 31881
rect 26421 31872 26433 31875
rect 26384 31844 26433 31872
rect 26384 31832 26390 31844
rect 26421 31841 26433 31844
rect 26467 31841 26479 31875
rect 26421 31835 26479 31841
rect 24820 31776 25728 31804
rect 25961 31807 26019 31813
rect 24820 31764 24826 31776
rect 25961 31773 25973 31807
rect 26007 31804 26019 31807
rect 26896 31804 26924 31912
rect 55125 31909 55137 31943
rect 55171 31909 55183 31943
rect 55125 31903 55183 31909
rect 55214 31900 55220 31952
rect 55272 31940 55278 31952
rect 55692 31940 55720 31968
rect 55769 31943 55827 31949
rect 55769 31940 55781 31943
rect 55272 31912 55317 31940
rect 55692 31912 55781 31940
rect 55272 31900 55278 31912
rect 55769 31909 55781 31912
rect 55815 31909 55827 31943
rect 57440 31940 57468 31980
rect 57609 31943 57667 31949
rect 57609 31940 57621 31943
rect 57440 31912 57621 31940
rect 55769 31903 55827 31909
rect 57609 31909 57621 31912
rect 57655 31909 57667 31943
rect 57609 31903 57667 31909
rect 58161 31943 58219 31949
rect 58161 31909 58173 31943
rect 58207 31940 58219 31943
rect 58342 31940 58348 31952
rect 58207 31912 58348 31940
rect 58207 31909 58219 31912
rect 58161 31903 58219 31909
rect 58342 31900 58348 31912
rect 58400 31900 58406 31952
rect 27332 31875 27390 31881
rect 27332 31841 27344 31875
rect 27378 31872 27390 31875
rect 27798 31872 27804 31884
rect 27378 31844 27804 31872
rect 27378 31841 27390 31844
rect 27332 31835 27390 31841
rect 27798 31832 27804 31844
rect 27856 31832 27862 31884
rect 30466 31832 30472 31884
rect 30524 31872 30530 31884
rect 32033 31875 32091 31881
rect 32033 31872 32045 31875
rect 30524 31844 32045 31872
rect 30524 31832 30530 31844
rect 32033 31841 32045 31844
rect 32079 31872 32091 31875
rect 32125 31875 32183 31881
rect 32125 31872 32137 31875
rect 32079 31844 32137 31872
rect 32079 31841 32091 31844
rect 32033 31835 32091 31841
rect 32125 31841 32137 31844
rect 32171 31841 32183 31875
rect 32125 31835 32183 31841
rect 32392 31875 32450 31881
rect 32392 31841 32404 31875
rect 32438 31872 32450 31875
rect 32950 31872 32956 31884
rect 32438 31844 32956 31872
rect 32438 31841 32450 31844
rect 32392 31835 32450 31841
rect 32950 31832 32956 31844
rect 33008 31832 33014 31884
rect 34422 31872 34428 31884
rect 34383 31844 34428 31872
rect 34422 31832 34428 31844
rect 34480 31832 34486 31884
rect 34514 31832 34520 31884
rect 34572 31872 34578 31884
rect 34793 31875 34851 31881
rect 34572 31844 34617 31872
rect 34572 31832 34578 31844
rect 34793 31841 34805 31875
rect 34839 31841 34851 31875
rect 35710 31872 35716 31884
rect 35671 31844 35716 31872
rect 34793 31835 34851 31841
rect 27062 31804 27068 31816
rect 26007 31776 26924 31804
rect 27023 31776 27068 31804
rect 26007 31773 26019 31776
rect 25961 31767 26019 31773
rect 27062 31764 27068 31776
rect 27120 31764 27126 31816
rect 34698 31804 34704 31816
rect 34659 31776 34704 31804
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34808 31804 34836 31835
rect 35710 31832 35716 31844
rect 35768 31832 35774 31884
rect 53834 31832 53840 31884
rect 53892 31872 53898 31884
rect 53929 31875 53987 31881
rect 53929 31872 53941 31875
rect 53892 31844 53941 31872
rect 53892 31832 53898 31844
rect 53929 31841 53941 31844
rect 53975 31841 53987 31875
rect 53929 31835 53987 31841
rect 54573 31875 54631 31881
rect 54573 31841 54585 31875
rect 54619 31872 54631 31875
rect 54662 31872 54668 31884
rect 54619 31844 54668 31872
rect 54619 31841 54631 31844
rect 54573 31835 54631 31841
rect 54662 31832 54668 31844
rect 54720 31832 54726 31884
rect 56686 31832 56692 31884
rect 56744 31872 56750 31884
rect 56781 31875 56839 31881
rect 56781 31872 56793 31875
rect 56744 31844 56793 31872
rect 56744 31832 56750 31844
rect 56781 31841 56793 31844
rect 56827 31841 56839 31875
rect 56962 31872 56968 31884
rect 56923 31844 56968 31872
rect 56781 31835 56839 31841
rect 56962 31832 56968 31844
rect 57020 31832 57026 31884
rect 35805 31807 35863 31813
rect 35805 31804 35817 31807
rect 34808 31776 35817 31804
rect 35805 31773 35817 31776
rect 35851 31804 35863 31807
rect 36170 31804 36176 31816
rect 35851 31776 36176 31804
rect 35851 31773 35863 31776
rect 35805 31767 35863 31773
rect 36170 31764 36176 31776
rect 36228 31764 36234 31816
rect 55214 31804 55220 31816
rect 53760 31776 55220 31804
rect 22738 31696 22744 31748
rect 22796 31736 22802 31748
rect 23474 31736 23480 31748
rect 22796 31708 23480 31736
rect 22796 31696 22802 31708
rect 23474 31696 23480 31708
rect 23532 31696 23538 31748
rect 53760 31745 53788 31776
rect 55214 31764 55220 31776
rect 55272 31764 55278 31816
rect 57333 31807 57391 31813
rect 57333 31773 57345 31807
rect 57379 31804 57391 31807
rect 57517 31807 57575 31813
rect 57517 31804 57529 31807
rect 57379 31776 57529 31804
rect 57379 31773 57391 31776
rect 57333 31767 57391 31773
rect 57517 31773 57529 31776
rect 57563 31804 57575 31807
rect 57882 31804 57888 31816
rect 57563 31776 57888 31804
rect 57563 31773 57575 31776
rect 57517 31767 57575 31773
rect 57882 31764 57888 31776
rect 57940 31764 57946 31816
rect 53745 31739 53803 31745
rect 53745 31705 53757 31739
rect 53791 31705 53803 31739
rect 53745 31699 53803 31705
rect 54389 31739 54447 31745
rect 54389 31705 54401 31739
rect 54435 31736 54447 31739
rect 54570 31736 54576 31748
rect 54435 31708 54576 31736
rect 54435 31705 54447 31708
rect 54389 31699 54447 31705
rect 54570 31696 54576 31708
rect 54628 31696 54634 31748
rect 20864 31640 21680 31668
rect 20864 31628 20870 31640
rect 23014 31628 23020 31680
rect 23072 31668 23078 31680
rect 23109 31671 23167 31677
rect 23109 31668 23121 31671
rect 23072 31640 23121 31668
rect 23072 31628 23078 31640
rect 23109 31637 23121 31640
rect 23155 31637 23167 31671
rect 28442 31668 28448 31680
rect 28403 31640 28448 31668
rect 23109 31631 23167 31637
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 33502 31668 33508 31680
rect 33463 31640 33508 31668
rect 33502 31628 33508 31640
rect 33560 31628 33566 31680
rect 1104 31578 58880 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 58880 31578
rect 1104 31504 58880 31526
rect 12066 31424 12072 31476
rect 12124 31464 12130 31476
rect 12250 31464 12256 31476
rect 12124 31436 12256 31464
rect 12124 31424 12130 31436
rect 12250 31424 12256 31436
rect 12308 31464 12314 31476
rect 12713 31467 12771 31473
rect 12713 31464 12725 31467
rect 12308 31436 12725 31464
rect 12308 31424 12314 31436
rect 12713 31433 12725 31436
rect 12759 31433 12771 31467
rect 12713 31427 12771 31433
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19521 31467 19579 31473
rect 19521 31464 19533 31467
rect 19392 31436 19533 31464
rect 19392 31424 19398 31436
rect 19521 31433 19533 31436
rect 19567 31433 19579 31467
rect 19521 31427 19579 31433
rect 21637 31467 21695 31473
rect 21637 31433 21649 31467
rect 21683 31464 21695 31467
rect 21818 31464 21824 31476
rect 21683 31436 21824 31464
rect 21683 31433 21695 31436
rect 21637 31427 21695 31433
rect 21818 31424 21824 31436
rect 21876 31424 21882 31476
rect 23658 31424 23664 31476
rect 23716 31464 23722 31476
rect 27062 31464 27068 31476
rect 23716 31436 27068 31464
rect 23716 31424 23722 31436
rect 12618 31405 12624 31408
rect 12602 31399 12624 31405
rect 12602 31396 12614 31399
rect 12531 31368 12614 31396
rect 12602 31365 12614 31368
rect 12676 31396 12682 31408
rect 13725 31399 13783 31405
rect 13725 31396 13737 31399
rect 12676 31368 13737 31396
rect 12602 31359 12624 31365
rect 12618 31356 12624 31359
rect 12676 31356 12682 31368
rect 13725 31365 13737 31368
rect 13771 31365 13783 31399
rect 19978 31396 19984 31408
rect 13725 31359 13783 31365
rect 15764 31368 19984 31396
rect 12805 31331 12863 31337
rect 12805 31297 12817 31331
rect 12851 31328 12863 31331
rect 13262 31328 13268 31340
rect 12851 31300 13268 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 13262 31288 13268 31300
rect 13320 31288 13326 31340
rect 15764 31337 15792 31368
rect 19978 31356 19984 31368
rect 20036 31356 20042 31408
rect 22830 31356 22836 31408
rect 22888 31356 22894 31408
rect 15749 31331 15807 31337
rect 15749 31297 15761 31331
rect 15795 31297 15807 31331
rect 18506 31328 18512 31340
rect 15749 31291 15807 31297
rect 17880 31300 18512 31328
rect 12342 31220 12348 31272
rect 12400 31260 12406 31272
rect 12437 31263 12495 31269
rect 12437 31260 12449 31263
rect 12400 31232 12449 31260
rect 12400 31220 12406 31232
rect 12437 31229 12449 31232
rect 12483 31229 12495 31263
rect 13630 31260 13636 31272
rect 13591 31232 13636 31260
rect 12437 31223 12495 31229
rect 13630 31220 13636 31232
rect 13688 31220 13694 31272
rect 14461 31263 14519 31269
rect 14461 31229 14473 31263
rect 14507 31260 14519 31263
rect 15194 31260 15200 31272
rect 14507 31232 15200 31260
rect 14507 31229 14519 31232
rect 14461 31223 14519 31229
rect 15194 31220 15200 31232
rect 15252 31220 15258 31272
rect 15473 31263 15531 31269
rect 15473 31229 15485 31263
rect 15519 31260 15531 31263
rect 15654 31260 15660 31272
rect 15519 31232 15660 31260
rect 15519 31229 15531 31232
rect 15473 31223 15531 31229
rect 15654 31220 15660 31232
rect 15712 31220 15718 31272
rect 17880 31269 17908 31300
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18874 31288 18880 31340
rect 18932 31328 18938 31340
rect 20165 31331 20223 31337
rect 20165 31328 20177 31331
rect 18932 31300 20177 31328
rect 18932 31288 18938 31300
rect 17865 31263 17923 31269
rect 17865 31229 17877 31263
rect 17911 31229 17923 31263
rect 17865 31223 17923 31229
rect 17957 31263 18015 31269
rect 17957 31229 17969 31263
rect 18003 31229 18015 31263
rect 17957 31223 18015 31229
rect 13170 31192 13176 31204
rect 13131 31164 13176 31192
rect 13170 31152 13176 31164
rect 13228 31152 13234 31204
rect 17494 31152 17500 31204
rect 17552 31192 17558 31204
rect 17972 31192 18000 31223
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 18233 31263 18291 31269
rect 18104 31232 18149 31260
rect 18104 31220 18110 31232
rect 18233 31229 18245 31263
rect 18279 31260 18291 31263
rect 18414 31260 18420 31272
rect 18279 31232 18420 31260
rect 18279 31229 18291 31232
rect 18233 31223 18291 31229
rect 18414 31220 18420 31232
rect 18472 31220 18478 31272
rect 19245 31263 19303 31269
rect 19245 31229 19257 31263
rect 19291 31229 19303 31263
rect 19245 31223 19303 31229
rect 19337 31263 19395 31269
rect 19337 31229 19349 31263
rect 19383 31260 19395 31263
rect 19426 31260 19432 31272
rect 19383 31232 19432 31260
rect 19383 31229 19395 31232
rect 19337 31223 19395 31229
rect 17552 31164 18000 31192
rect 19260 31192 19288 31223
rect 19426 31220 19432 31232
rect 19484 31220 19490 31272
rect 19628 31269 19656 31300
rect 20165 31297 20177 31300
rect 20211 31297 20223 31331
rect 21634 31328 21640 31340
rect 20165 31291 20223 31297
rect 21376 31300 21640 31328
rect 19613 31263 19671 31269
rect 19613 31229 19625 31263
rect 19659 31229 19671 31263
rect 20070 31260 20076 31272
rect 20031 31232 20076 31260
rect 19613 31223 19671 31229
rect 20070 31220 20076 31232
rect 20128 31220 20134 31272
rect 21174 31269 21180 31272
rect 20993 31263 21051 31269
rect 20993 31229 21005 31263
rect 21039 31229 21051 31263
rect 20993 31223 21051 31229
rect 21141 31263 21180 31269
rect 21141 31229 21153 31263
rect 21141 31223 21180 31229
rect 20088 31192 20116 31220
rect 19260 31164 20116 31192
rect 17552 31152 17558 31164
rect 14550 31124 14556 31136
rect 14511 31096 14556 31124
rect 14550 31084 14556 31096
rect 14608 31084 14614 31136
rect 17586 31124 17592 31136
rect 17547 31096 17592 31124
rect 17586 31084 17592 31096
rect 17644 31084 17650 31136
rect 19061 31127 19119 31133
rect 19061 31093 19073 31127
rect 19107 31124 19119 31127
rect 19150 31124 19156 31136
rect 19107 31096 19156 31124
rect 19107 31093 19119 31096
rect 19061 31087 19119 31093
rect 19150 31084 19156 31096
rect 19208 31084 19214 31136
rect 19426 31084 19432 31136
rect 19484 31124 19490 31136
rect 20622 31124 20628 31136
rect 19484 31096 20628 31124
rect 19484 31084 19490 31096
rect 20622 31084 20628 31096
rect 20680 31124 20686 31136
rect 21008 31124 21036 31223
rect 21174 31220 21180 31223
rect 21232 31220 21238 31272
rect 21376 31269 21404 31300
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 22094 31288 22100 31340
rect 22152 31328 22158 31340
rect 22848 31328 22876 31356
rect 23017 31331 23075 31337
rect 23017 31328 23029 31331
rect 22152 31300 23029 31328
rect 22152 31288 22158 31300
rect 23017 31297 23029 31300
rect 23063 31297 23075 31331
rect 23017 31291 23075 31297
rect 23474 31288 23480 31340
rect 23532 31328 23538 31340
rect 25148 31337 25176 31436
rect 27062 31424 27068 31436
rect 27120 31464 27126 31476
rect 27246 31464 27252 31476
rect 27120 31436 27252 31464
rect 27120 31424 27126 31436
rect 27246 31424 27252 31436
rect 27304 31424 27310 31476
rect 27798 31464 27804 31476
rect 27759 31436 27804 31464
rect 27798 31424 27804 31436
rect 27856 31424 27862 31476
rect 32950 31424 32956 31476
rect 33008 31464 33014 31476
rect 33045 31467 33103 31473
rect 33045 31464 33057 31467
rect 33008 31436 33057 31464
rect 33008 31424 33014 31436
rect 33045 31433 33057 31436
rect 33091 31433 33103 31467
rect 33045 31427 33103 31433
rect 33134 31424 33140 31476
rect 33192 31464 33198 31476
rect 33413 31467 33471 31473
rect 33413 31464 33425 31467
rect 33192 31436 33425 31464
rect 33192 31424 33198 31436
rect 33413 31433 33425 31436
rect 33459 31433 33471 31467
rect 34054 31464 34060 31476
rect 34015 31436 34060 31464
rect 33413 31427 33471 31433
rect 34054 31424 34060 31436
rect 34112 31424 34118 31476
rect 34514 31424 34520 31476
rect 34572 31464 34578 31476
rect 34701 31467 34759 31473
rect 34701 31464 34713 31467
rect 34572 31436 34713 31464
rect 34572 31424 34578 31436
rect 34701 31433 34713 31436
rect 34747 31433 34759 31467
rect 34701 31427 34759 31433
rect 56502 31396 56508 31408
rect 52932 31368 56508 31396
rect 23569 31331 23627 31337
rect 23569 31328 23581 31331
rect 23532 31300 23581 31328
rect 23532 31288 23538 31300
rect 23569 31297 23581 31300
rect 23615 31328 23627 31331
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 23615 31300 24133 31328
rect 23615 31297 23627 31300
rect 23569 31291 23627 31297
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 33502 31328 33508 31340
rect 33463 31300 33508 31328
rect 25133 31291 25191 31297
rect 33502 31288 33508 31300
rect 33560 31328 33566 31340
rect 33560 31300 34008 31328
rect 33560 31288 33566 31300
rect 21361 31263 21419 31269
rect 21361 31229 21373 31263
rect 21407 31229 21419 31263
rect 21361 31223 21419 31229
rect 21450 31220 21456 31272
rect 21508 31269 21514 31272
rect 21508 31260 21516 31269
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 21508 31232 22569 31260
rect 21508 31223 21516 31232
rect 22557 31229 22569 31232
rect 22603 31229 22615 31263
rect 22738 31260 22744 31272
rect 22699 31232 22744 31260
rect 22557 31223 22615 31229
rect 21508 31220 21514 31223
rect 22738 31220 22744 31232
rect 22796 31220 22802 31272
rect 22833 31263 22891 31269
rect 22833 31229 22845 31263
rect 22879 31229 22891 31263
rect 23106 31260 23112 31272
rect 23067 31232 23112 31260
rect 22833 31223 22891 31229
rect 21269 31195 21327 31201
rect 21269 31161 21281 31195
rect 21315 31161 21327 31195
rect 22462 31192 22468 31204
rect 21269 31155 21327 31161
rect 21560 31164 22468 31192
rect 20680 31096 21036 31124
rect 21284 31124 21312 31155
rect 21560 31124 21588 31164
rect 22462 31152 22468 31164
rect 22520 31152 22526 31204
rect 22848 31192 22876 31223
rect 23106 31220 23112 31232
rect 23164 31220 23170 31272
rect 23753 31263 23811 31269
rect 23753 31229 23765 31263
rect 23799 31229 23811 31263
rect 23753 31223 23811 31229
rect 23474 31192 23480 31204
rect 22848 31164 23480 31192
rect 23474 31152 23480 31164
rect 23532 31192 23538 31204
rect 23768 31192 23796 31223
rect 23842 31220 23848 31272
rect 23900 31260 23906 31272
rect 24670 31260 24676 31272
rect 23900 31232 24676 31260
rect 23900 31220 23906 31232
rect 24670 31220 24676 31232
rect 24728 31260 24734 31272
rect 27801 31263 27859 31269
rect 27801 31260 27813 31263
rect 24728 31232 27813 31260
rect 24728 31220 24734 31232
rect 27801 31229 27813 31232
rect 27847 31229 27859 31263
rect 27801 31223 27859 31229
rect 27985 31263 28043 31269
rect 27985 31229 27997 31263
rect 28031 31260 28043 31263
rect 28166 31260 28172 31272
rect 28031 31232 28172 31260
rect 28031 31229 28043 31232
rect 27985 31223 28043 31229
rect 28166 31220 28172 31232
rect 28224 31220 28230 31272
rect 33980 31269 34008 31300
rect 33229 31263 33287 31269
rect 33229 31229 33241 31263
rect 33275 31229 33287 31263
rect 33229 31223 33287 31229
rect 33965 31263 34023 31269
rect 33965 31229 33977 31263
rect 34011 31229 34023 31263
rect 33965 31223 34023 31229
rect 34609 31263 34667 31269
rect 34609 31229 34621 31263
rect 34655 31260 34667 31263
rect 34698 31260 34704 31272
rect 34655 31232 34704 31260
rect 34655 31229 34667 31232
rect 34609 31223 34667 31229
rect 24029 31195 24087 31201
rect 24029 31192 24041 31195
rect 23532 31164 24041 31192
rect 23532 31152 23538 31164
rect 24029 31161 24041 31164
rect 24075 31161 24087 31195
rect 24029 31155 24087 31161
rect 25400 31195 25458 31201
rect 25400 31161 25412 31195
rect 25446 31192 25458 31195
rect 25958 31192 25964 31204
rect 25446 31164 25964 31192
rect 25446 31161 25458 31164
rect 25400 31155 25458 31161
rect 25958 31152 25964 31164
rect 26016 31152 26022 31204
rect 33244 31192 33272 31223
rect 34624 31192 34652 31223
rect 34698 31220 34704 31232
rect 34756 31220 34762 31272
rect 52932 31269 52960 31368
rect 56502 31356 56508 31368
rect 56560 31356 56566 31408
rect 56870 31328 56876 31340
rect 55324 31300 56876 31328
rect 52917 31263 52975 31269
rect 52917 31229 52929 31263
rect 52963 31229 52975 31263
rect 52917 31223 52975 31229
rect 33244 31164 34652 31192
rect 36538 31152 36544 31204
rect 36596 31192 36602 31204
rect 54481 31195 54539 31201
rect 54481 31192 54493 31195
rect 36596 31164 54493 31192
rect 36596 31152 36602 31164
rect 54481 31161 54493 31164
rect 54527 31161 54539 31195
rect 54481 31155 54539 31161
rect 54570 31152 54576 31204
rect 54628 31192 54634 31204
rect 55125 31195 55183 31201
rect 54628 31164 54673 31192
rect 54628 31152 54634 31164
rect 55125 31161 55137 31195
rect 55171 31192 55183 31195
rect 55324 31192 55352 31300
rect 56870 31288 56876 31300
rect 56928 31288 56934 31340
rect 58161 31331 58219 31337
rect 58161 31297 58173 31331
rect 58207 31328 58219 31331
rect 58434 31328 58440 31340
rect 58207 31300 58440 31328
rect 58207 31297 58219 31300
rect 58161 31291 58219 31297
rect 58434 31288 58440 31300
rect 58492 31288 58498 31340
rect 55585 31263 55643 31269
rect 55585 31229 55597 31263
rect 55631 31229 55643 31263
rect 56226 31260 56232 31272
rect 56187 31232 56232 31260
rect 55585 31223 55643 31229
rect 55171 31164 55352 31192
rect 55600 31192 55628 31223
rect 56226 31220 56232 31232
rect 56284 31220 56290 31272
rect 57149 31195 57207 31201
rect 55600 31164 56456 31192
rect 55171 31161 55183 31164
rect 55125 31155 55183 31161
rect 21284 31096 21588 31124
rect 20680 31084 20686 31096
rect 23290 31084 23296 31136
rect 23348 31124 23354 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23348 31096 23949 31124
rect 23348 31084 23354 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 26510 31124 26516 31136
rect 26471 31096 26516 31124
rect 23937 31087 23995 31093
rect 26510 31084 26516 31096
rect 26568 31084 26574 31136
rect 55030 31084 55036 31136
rect 55088 31124 55094 31136
rect 55600 31124 55628 31164
rect 55766 31124 55772 31136
rect 55088 31096 55628 31124
rect 55727 31096 55772 31124
rect 55088 31084 55094 31096
rect 55766 31084 55772 31096
rect 55824 31084 55830 31136
rect 56428 31133 56456 31164
rect 57149 31161 57161 31195
rect 57195 31161 57207 31195
rect 57149 31155 57207 31161
rect 56413 31127 56471 31133
rect 56413 31093 56425 31127
rect 56459 31093 56471 31127
rect 56870 31124 56876 31136
rect 56831 31096 56876 31124
rect 56413 31087 56471 31093
rect 56870 31084 56876 31096
rect 56928 31124 56934 31136
rect 57164 31124 57192 31155
rect 57238 31152 57244 31204
rect 57296 31192 57302 31204
rect 57296 31164 57341 31192
rect 57296 31152 57302 31164
rect 56928 31096 57192 31124
rect 56928 31084 56934 31096
rect 1104 31034 58880 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 50326 31034
rect 50378 30982 50390 31034
rect 50442 30982 50454 31034
rect 50506 30982 50518 31034
rect 50570 30982 58880 31034
rect 1104 30960 58880 30982
rect 11422 30880 11428 30932
rect 11480 30920 11486 30932
rect 13633 30923 13691 30929
rect 13633 30920 13645 30923
rect 11480 30892 13645 30920
rect 11480 30880 11486 30892
rect 13633 30889 13645 30892
rect 13679 30920 13691 30923
rect 13906 30920 13912 30932
rect 13679 30892 13912 30920
rect 13679 30889 13691 30892
rect 13633 30883 13691 30889
rect 13906 30880 13912 30892
rect 13964 30880 13970 30932
rect 15378 30920 15384 30932
rect 15339 30892 15384 30920
rect 15378 30880 15384 30892
rect 15436 30920 15442 30932
rect 16390 30920 16396 30932
rect 15436 30892 16396 30920
rect 15436 30880 15442 30892
rect 16390 30880 16396 30892
rect 16448 30880 16454 30932
rect 18414 30920 18420 30932
rect 18375 30892 18420 30920
rect 18414 30880 18420 30892
rect 18472 30880 18478 30932
rect 20070 30880 20076 30932
rect 20128 30920 20134 30932
rect 21361 30923 21419 30929
rect 21361 30920 21373 30923
rect 20128 30892 21373 30920
rect 20128 30880 20134 30892
rect 21361 30889 21373 30892
rect 21407 30889 21419 30923
rect 21361 30883 21419 30889
rect 21913 30923 21971 30929
rect 21913 30889 21925 30923
rect 21959 30920 21971 30923
rect 22462 30920 22468 30932
rect 21959 30892 22468 30920
rect 21959 30889 21971 30892
rect 21913 30883 21971 30889
rect 22462 30880 22468 30892
rect 22520 30880 22526 30932
rect 25958 30920 25964 30932
rect 25919 30892 25964 30920
rect 25958 30880 25964 30892
rect 26016 30880 26022 30932
rect 28813 30923 28871 30929
rect 28813 30920 28825 30923
rect 26712 30892 28825 30920
rect 11164 30824 11928 30852
rect 1394 30784 1400 30796
rect 1355 30756 1400 30784
rect 1394 30744 1400 30756
rect 1452 30744 1458 30796
rect 10502 30784 10508 30796
rect 10463 30756 10508 30784
rect 10502 30744 10508 30756
rect 10560 30744 10566 30796
rect 11164 30793 11192 30824
rect 10965 30787 11023 30793
rect 10965 30753 10977 30787
rect 11011 30753 11023 30787
rect 10965 30747 11023 30753
rect 11149 30787 11207 30793
rect 11149 30753 11161 30787
rect 11195 30753 11207 30787
rect 11149 30747 11207 30753
rect 11793 30787 11851 30793
rect 11793 30753 11805 30787
rect 11839 30753 11851 30787
rect 11900 30784 11928 30824
rect 12434 30812 12440 30864
rect 12492 30852 12498 30864
rect 16200 30855 16258 30861
rect 12492 30824 12537 30852
rect 13832 30824 16160 30852
rect 12492 30812 12498 30824
rect 12986 30784 12992 30796
rect 11900 30756 12992 30784
rect 11793 30747 11851 30753
rect 10980 30716 11008 30747
rect 11514 30716 11520 30728
rect 10980 30688 11520 30716
rect 11514 30676 11520 30688
rect 11572 30676 11578 30728
rect 11808 30648 11836 30747
rect 12986 30744 12992 30756
rect 13044 30744 13050 30796
rect 13832 30793 13860 30824
rect 13817 30787 13875 30793
rect 13817 30753 13829 30787
rect 13863 30753 13875 30787
rect 13817 30747 13875 30753
rect 15197 30787 15255 30793
rect 15197 30753 15209 30787
rect 15243 30784 15255 30787
rect 15289 30787 15347 30793
rect 15289 30784 15301 30787
rect 15243 30756 15301 30784
rect 15243 30753 15255 30756
rect 15197 30747 15255 30753
rect 15289 30753 15301 30756
rect 15335 30753 15347 30787
rect 16132 30784 16160 30824
rect 16200 30821 16212 30855
rect 16246 30852 16258 30855
rect 17586 30852 17592 30864
rect 16246 30824 17592 30852
rect 16246 30821 16258 30824
rect 16200 30815 16258 30821
rect 17586 30812 17592 30824
rect 17644 30812 17650 30864
rect 18049 30855 18107 30861
rect 18049 30821 18061 30855
rect 18095 30852 18107 30855
rect 18598 30852 18604 30864
rect 18095 30824 18604 30852
rect 18095 30821 18107 30824
rect 18049 30815 18107 30821
rect 18598 30812 18604 30824
rect 18656 30852 18662 30864
rect 18969 30855 19027 30861
rect 18969 30852 18981 30855
rect 18656 30824 18981 30852
rect 18656 30812 18662 30824
rect 18969 30821 18981 30824
rect 19015 30821 19027 30855
rect 20530 30852 20536 30864
rect 18969 30815 19027 30821
rect 20088 30824 20536 30852
rect 20088 30796 20116 30824
rect 20530 30812 20536 30824
rect 20588 30812 20594 30864
rect 23032 30824 25268 30852
rect 16758 30784 16764 30796
rect 16132 30756 16764 30784
rect 15289 30747 15347 30753
rect 16758 30744 16764 30756
rect 16816 30744 16822 30796
rect 17954 30793 17960 30796
rect 17773 30787 17831 30793
rect 17773 30753 17785 30787
rect 17819 30753 17831 30787
rect 17773 30747 17831 30753
rect 17921 30787 17960 30793
rect 17921 30753 17933 30787
rect 17921 30747 17960 30753
rect 11885 30719 11943 30725
rect 11885 30685 11897 30719
rect 11931 30716 11943 30719
rect 12526 30716 12532 30728
rect 11931 30688 12532 30716
rect 11931 30685 11943 30688
rect 11885 30679 11943 30685
rect 12526 30676 12532 30688
rect 12584 30676 12590 30728
rect 12805 30719 12863 30725
rect 12805 30685 12817 30719
rect 12851 30716 12863 30719
rect 12894 30716 12900 30728
rect 12851 30688 12900 30716
rect 12851 30685 12863 30688
rect 12805 30679 12863 30685
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 14366 30676 14372 30728
rect 14424 30716 14430 30728
rect 15102 30716 15108 30728
rect 14424 30688 15108 30716
rect 14424 30676 14430 30688
rect 15102 30676 15108 30688
rect 15160 30716 15166 30728
rect 15933 30719 15991 30725
rect 15933 30716 15945 30719
rect 15160 30688 15945 30716
rect 15160 30676 15166 30688
rect 15933 30685 15945 30688
rect 15979 30685 15991 30719
rect 15933 30679 15991 30685
rect 12250 30648 12256 30660
rect 11808 30620 12256 30648
rect 12250 30608 12256 30620
rect 12308 30648 12314 30660
rect 12713 30651 12771 30657
rect 12713 30648 12725 30651
rect 12308 30620 12725 30648
rect 12308 30608 12314 30620
rect 12713 30617 12725 30620
rect 12759 30617 12771 30651
rect 17788 30648 17816 30747
rect 17954 30744 17960 30747
rect 18012 30744 18018 30796
rect 18138 30784 18144 30796
rect 18099 30756 18144 30784
rect 18138 30744 18144 30756
rect 18196 30744 18202 30796
rect 18322 30793 18328 30796
rect 18279 30787 18328 30793
rect 18279 30753 18291 30787
rect 18325 30753 18328 30787
rect 18279 30747 18328 30753
rect 18322 30744 18328 30747
rect 18380 30744 18386 30796
rect 18877 30787 18935 30793
rect 18877 30753 18889 30787
rect 18923 30753 18935 30787
rect 18877 30747 18935 30753
rect 19981 30787 20039 30793
rect 19981 30753 19993 30787
rect 20027 30784 20039 30787
rect 20070 30784 20076 30796
rect 20027 30756 20076 30784
rect 20027 30753 20039 30756
rect 19981 30747 20039 30753
rect 18156 30716 18184 30744
rect 18892 30716 18920 30747
rect 20070 30744 20076 30756
rect 20128 30744 20134 30796
rect 20254 30793 20260 30796
rect 20248 30747 20260 30793
rect 20312 30784 20318 30796
rect 20312 30756 20348 30784
rect 20254 30744 20260 30747
rect 20312 30744 20318 30756
rect 21634 30744 21640 30796
rect 21692 30784 21698 30796
rect 21821 30787 21879 30793
rect 21821 30784 21833 30787
rect 21692 30756 21833 30784
rect 21692 30744 21698 30756
rect 21821 30753 21833 30756
rect 21867 30753 21879 30787
rect 21821 30747 21879 30753
rect 22370 30744 22376 30796
rect 22428 30784 22434 30796
rect 23032 30793 23060 30824
rect 23017 30787 23075 30793
rect 23017 30784 23029 30787
rect 22428 30756 23029 30784
rect 22428 30744 22434 30756
rect 23017 30753 23029 30756
rect 23063 30753 23075 30787
rect 23017 30747 23075 30753
rect 23201 30787 23259 30793
rect 23201 30753 23213 30787
rect 23247 30753 23259 30787
rect 23201 30747 23259 30753
rect 18156 30688 18920 30716
rect 19426 30648 19432 30660
rect 17788 30620 19432 30648
rect 12713 30611 12771 30617
rect 19426 30608 19432 30620
rect 19484 30608 19490 30660
rect 22462 30608 22468 30660
rect 22520 30648 22526 30660
rect 23216 30648 23244 30747
rect 23290 30744 23296 30796
rect 23348 30784 23354 30796
rect 23569 30787 23627 30793
rect 23348 30756 23393 30784
rect 23348 30744 23354 30756
rect 23569 30753 23581 30787
rect 23615 30784 23627 30787
rect 23658 30784 23664 30796
rect 23615 30756 23664 30784
rect 23615 30753 23627 30756
rect 23569 30747 23627 30753
rect 23658 30744 23664 30756
rect 23716 30784 23722 30796
rect 25240 30793 25268 30824
rect 25332 30824 25820 30852
rect 25225 30787 25283 30793
rect 23716 30756 25176 30784
rect 23716 30744 23722 30756
rect 23385 30719 23443 30725
rect 23385 30685 23397 30719
rect 23431 30716 23443 30719
rect 23934 30716 23940 30728
rect 23431 30688 23940 30716
rect 23431 30685 23443 30688
rect 23385 30679 23443 30685
rect 23934 30676 23940 30688
rect 23992 30716 23998 30728
rect 24486 30716 24492 30728
rect 23992 30688 24492 30716
rect 23992 30676 23998 30688
rect 24486 30676 24492 30688
rect 24544 30676 24550 30728
rect 25148 30716 25176 30756
rect 25225 30753 25237 30787
rect 25271 30753 25283 30787
rect 25225 30747 25283 30753
rect 25332 30716 25360 30824
rect 25792 30793 25820 30824
rect 25409 30787 25467 30793
rect 25409 30753 25421 30787
rect 25455 30753 25467 30787
rect 25409 30747 25467 30753
rect 25504 30787 25562 30793
rect 25504 30753 25516 30787
rect 25550 30753 25562 30787
rect 25504 30747 25562 30753
rect 25777 30787 25835 30793
rect 25777 30753 25789 30787
rect 25823 30753 25835 30787
rect 25777 30747 25835 30753
rect 25148 30688 25360 30716
rect 25424 30648 25452 30747
rect 25516 30660 25544 30747
rect 26510 30744 26516 30796
rect 26568 30784 26574 30796
rect 26712 30793 26740 30892
rect 28813 30889 28825 30892
rect 28859 30889 28871 30923
rect 28813 30883 28871 30889
rect 54297 30923 54355 30929
rect 54297 30889 54309 30923
rect 54343 30920 54355 30923
rect 54570 30920 54576 30932
rect 54343 30892 54576 30920
rect 54343 30889 54355 30892
rect 54297 30883 54355 30889
rect 26605 30787 26663 30793
rect 26605 30784 26617 30787
rect 26568 30756 26617 30784
rect 26568 30744 26574 30756
rect 26605 30753 26617 30756
rect 26651 30753 26663 30787
rect 26605 30747 26663 30753
rect 26697 30787 26755 30793
rect 26697 30753 26709 30787
rect 26743 30753 26755 30787
rect 26970 30784 26976 30796
rect 26931 30756 26976 30784
rect 26697 30747 26755 30753
rect 26970 30744 26976 30756
rect 27028 30744 27034 30796
rect 27700 30787 27758 30793
rect 27700 30753 27712 30787
rect 27746 30784 27758 30787
rect 28828 30784 28856 30883
rect 54570 30880 54576 30892
rect 54628 30880 54634 30932
rect 54941 30923 54999 30929
rect 54941 30889 54953 30923
rect 54987 30920 54999 30923
rect 56410 30920 56416 30932
rect 54987 30892 56416 30920
rect 54987 30889 54999 30892
rect 54941 30883 54999 30889
rect 56410 30880 56416 30892
rect 56468 30880 56474 30932
rect 55766 30812 55772 30864
rect 55824 30852 55830 30864
rect 56873 30855 56931 30861
rect 56873 30852 56885 30855
rect 55824 30824 56885 30852
rect 55824 30812 55830 30824
rect 56873 30821 56885 30824
rect 56919 30821 56931 30855
rect 57790 30852 57796 30864
rect 57751 30824 57796 30852
rect 56873 30815 56931 30821
rect 57790 30812 57796 30824
rect 57848 30812 57854 30864
rect 29273 30787 29331 30793
rect 29273 30784 29285 30787
rect 27746 30756 28764 30784
rect 28828 30756 29285 30784
rect 27746 30753 27758 30756
rect 27700 30747 27758 30753
rect 25593 30719 25651 30725
rect 25593 30685 25605 30719
rect 25639 30716 25651 30719
rect 26528 30716 26556 30744
rect 25639 30688 26556 30716
rect 25639 30685 25651 30688
rect 25593 30679 25651 30685
rect 27246 30676 27252 30728
rect 27304 30716 27310 30728
rect 27433 30719 27491 30725
rect 27433 30716 27445 30719
rect 27304 30688 27445 30716
rect 27304 30676 27310 30688
rect 27433 30685 27445 30688
rect 27479 30685 27491 30719
rect 28736 30716 28764 30756
rect 29273 30753 29285 30756
rect 29319 30753 29331 30787
rect 29273 30747 29331 30753
rect 53834 30744 53840 30796
rect 53892 30784 53898 30796
rect 54481 30787 54539 30793
rect 54481 30784 54493 30787
rect 53892 30756 54493 30784
rect 53892 30744 53898 30756
rect 54481 30753 54493 30756
rect 54527 30753 54539 30787
rect 54481 30747 54539 30753
rect 55030 30744 55036 30796
rect 55088 30784 55094 30796
rect 55125 30787 55183 30793
rect 55125 30784 55137 30787
rect 55088 30756 55137 30784
rect 55088 30744 55094 30756
rect 55125 30753 55137 30756
rect 55171 30784 55183 30787
rect 55585 30787 55643 30793
rect 55585 30784 55597 30787
rect 55171 30756 55597 30784
rect 55171 30753 55183 30756
rect 55125 30747 55183 30753
rect 55585 30753 55597 30756
rect 55631 30753 55643 30787
rect 55585 30747 55643 30753
rect 29822 30716 29828 30728
rect 28736 30688 29828 30716
rect 27433 30679 27491 30685
rect 29822 30676 29828 30688
rect 29880 30676 29886 30728
rect 56781 30719 56839 30725
rect 56781 30685 56793 30719
rect 56827 30716 56839 30719
rect 56962 30716 56968 30728
rect 56827 30688 56968 30716
rect 56827 30685 56839 30688
rect 56781 30679 56839 30685
rect 56962 30676 56968 30688
rect 57020 30676 57026 30728
rect 22520 30620 25452 30648
rect 22520 30608 22526 30620
rect 25498 30608 25504 30660
rect 25556 30608 25562 30660
rect 53837 30651 53895 30657
rect 53837 30617 53849 30651
rect 53883 30648 53895 30651
rect 55769 30651 55827 30657
rect 53883 30620 55214 30648
rect 53883 30617 53895 30620
rect 53837 30611 53895 30617
rect 8754 30540 8760 30592
rect 8812 30580 8818 30592
rect 10321 30583 10379 30589
rect 10321 30580 10333 30583
rect 8812 30552 10333 30580
rect 8812 30540 8818 30552
rect 10321 30549 10333 30552
rect 10367 30549 10379 30583
rect 10321 30543 10379 30549
rect 10410 30540 10416 30592
rect 10468 30580 10474 30592
rect 10965 30583 11023 30589
rect 10965 30580 10977 30583
rect 10468 30552 10977 30580
rect 10468 30540 10474 30552
rect 10965 30549 10977 30552
rect 11011 30549 11023 30583
rect 10965 30543 11023 30549
rect 12602 30583 12660 30589
rect 12602 30549 12614 30583
rect 12648 30580 12660 30583
rect 12802 30580 12808 30592
rect 12648 30552 12808 30580
rect 12648 30549 12660 30552
rect 12602 30543 12660 30549
rect 12802 30540 12808 30552
rect 12860 30540 12866 30592
rect 13081 30583 13139 30589
rect 13081 30549 13093 30583
rect 13127 30580 13139 30583
rect 13722 30580 13728 30592
rect 13127 30552 13728 30580
rect 13127 30549 13139 30552
rect 13081 30543 13139 30549
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 15197 30583 15255 30589
rect 15197 30549 15209 30583
rect 15243 30580 15255 30583
rect 16666 30580 16672 30592
rect 15243 30552 16672 30580
rect 15243 30549 15255 30552
rect 15197 30543 15255 30549
rect 16666 30540 16672 30552
rect 16724 30580 16730 30592
rect 17313 30583 17371 30589
rect 17313 30580 17325 30583
rect 16724 30552 17325 30580
rect 16724 30540 16730 30552
rect 17313 30549 17325 30552
rect 17359 30580 17371 30583
rect 17494 30580 17500 30592
rect 17359 30552 17500 30580
rect 17359 30549 17371 30552
rect 17313 30543 17371 30549
rect 17494 30540 17500 30552
rect 17552 30540 17558 30592
rect 17954 30540 17960 30592
rect 18012 30580 18018 30592
rect 20714 30580 20720 30592
rect 18012 30552 20720 30580
rect 18012 30540 18018 30552
rect 20714 30540 20720 30552
rect 20772 30540 20778 30592
rect 23750 30580 23756 30592
rect 23711 30552 23756 30580
rect 23750 30540 23756 30552
rect 23808 30540 23814 30592
rect 26421 30583 26479 30589
rect 26421 30549 26433 30583
rect 26467 30580 26479 30583
rect 26694 30580 26700 30592
rect 26467 30552 26700 30580
rect 26467 30549 26479 30552
rect 26421 30543 26479 30549
rect 26694 30540 26700 30552
rect 26752 30540 26758 30592
rect 26786 30540 26792 30592
rect 26844 30580 26850 30592
rect 26881 30583 26939 30589
rect 26881 30580 26893 30583
rect 26844 30552 26893 30580
rect 26844 30540 26850 30552
rect 26881 30549 26893 30552
rect 26927 30580 26939 30583
rect 29365 30583 29423 30589
rect 29365 30580 29377 30583
rect 26927 30552 29377 30580
rect 26927 30549 26939 30552
rect 26881 30543 26939 30549
rect 29365 30549 29377 30552
rect 29411 30580 29423 30583
rect 30098 30580 30104 30592
rect 29411 30552 30104 30580
rect 29411 30549 29423 30552
rect 29365 30543 29423 30549
rect 30098 30540 30104 30552
rect 30156 30540 30162 30592
rect 55186 30580 55214 30620
rect 55769 30617 55781 30651
rect 55815 30648 55827 30651
rect 57238 30648 57244 30660
rect 55815 30620 57244 30648
rect 55815 30617 55827 30620
rect 55769 30611 55827 30617
rect 57238 30608 57244 30620
rect 57296 30608 57302 30660
rect 55674 30580 55680 30592
rect 55186 30552 55680 30580
rect 55674 30540 55680 30552
rect 55732 30540 55738 30592
rect 56597 30583 56655 30589
rect 56597 30549 56609 30583
rect 56643 30580 56655 30583
rect 56962 30580 56968 30592
rect 56643 30552 56968 30580
rect 56643 30549 56655 30552
rect 56597 30543 56655 30549
rect 56962 30540 56968 30552
rect 57020 30540 57026 30592
rect 1104 30490 58880 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 58880 30490
rect 1104 30416 58880 30438
rect 10321 30379 10379 30385
rect 10321 30345 10333 30379
rect 10367 30376 10379 30379
rect 10502 30376 10508 30388
rect 10367 30348 10508 30376
rect 10367 30345 10379 30348
rect 10321 30339 10379 30345
rect 1394 30172 1400 30184
rect 1355 30144 1400 30172
rect 1394 30132 1400 30144
rect 1452 30132 1458 30184
rect 9677 30175 9735 30181
rect 9677 30141 9689 30175
rect 9723 30172 9735 30175
rect 10336 30172 10364 30339
rect 10502 30336 10508 30348
rect 10560 30336 10566 30388
rect 12713 30379 12771 30385
rect 12713 30345 12725 30379
rect 12759 30376 12771 30379
rect 12802 30376 12808 30388
rect 12759 30348 12808 30376
rect 12759 30345 12771 30348
rect 12713 30339 12771 30345
rect 12802 30336 12808 30348
rect 12860 30376 12866 30388
rect 13630 30376 13636 30388
rect 12860 30348 13636 30376
rect 12860 30336 12866 30348
rect 13630 30336 13636 30348
rect 13688 30336 13694 30388
rect 13814 30376 13820 30388
rect 13775 30348 13820 30376
rect 13814 30336 13820 30348
rect 13872 30336 13878 30388
rect 18322 30376 18328 30388
rect 18235 30348 18328 30376
rect 18322 30336 18328 30348
rect 18380 30376 18386 30388
rect 20165 30379 20223 30385
rect 18380 30348 19012 30376
rect 18380 30336 18386 30348
rect 12526 30268 12532 30320
rect 12584 30317 12590 30320
rect 12584 30311 12633 30317
rect 12584 30277 12587 30311
rect 12621 30277 12633 30311
rect 12894 30308 12900 30320
rect 12584 30271 12633 30277
rect 12820 30280 12900 30308
rect 12584 30268 12590 30271
rect 11422 30240 11428 30252
rect 10520 30212 11428 30240
rect 10520 30181 10548 30212
rect 11422 30200 11428 30212
rect 11480 30200 11486 30252
rect 12250 30200 12256 30252
rect 12308 30240 12314 30252
rect 12820 30249 12848 30280
rect 12894 30268 12900 30280
rect 12952 30268 12958 30320
rect 15838 30268 15844 30320
rect 15896 30308 15902 30320
rect 16025 30311 16083 30317
rect 16025 30308 16037 30311
rect 15896 30280 16037 30308
rect 15896 30268 15902 30280
rect 16025 30277 16037 30280
rect 16071 30308 16083 30311
rect 17773 30311 17831 30317
rect 16071 30280 17264 30308
rect 16071 30277 16083 30280
rect 16025 30271 16083 30277
rect 12805 30243 12863 30249
rect 12308 30212 12756 30240
rect 12308 30200 12314 30212
rect 9723 30144 10364 30172
rect 10505 30175 10563 30181
rect 9723 30141 9735 30144
rect 9677 30135 9735 30141
rect 10505 30141 10517 30175
rect 10551 30141 10563 30175
rect 10962 30172 10968 30184
rect 10923 30144 10968 30172
rect 10505 30135 10563 30141
rect 10962 30132 10968 30144
rect 11020 30132 11026 30184
rect 12434 30132 12440 30184
rect 12492 30172 12498 30184
rect 12728 30172 12756 30212
rect 12805 30209 12817 30243
rect 12851 30209 12863 30243
rect 14093 30243 14151 30249
rect 14093 30240 14105 30243
rect 12805 30203 12863 30209
rect 12912 30212 14105 30240
rect 12912 30172 12940 30212
rect 14093 30209 14105 30212
rect 14139 30209 14151 30243
rect 16226 30243 16284 30249
rect 16226 30240 16238 30243
rect 14093 30203 14151 30209
rect 15672 30212 16238 30240
rect 12492 30144 12537 30172
rect 12728 30144 12940 30172
rect 12492 30132 12498 30144
rect 13170 30132 13176 30184
rect 13228 30172 13234 30184
rect 13633 30175 13691 30181
rect 13633 30172 13645 30175
rect 13228 30144 13645 30172
rect 13228 30132 13234 30144
rect 13633 30141 13645 30144
rect 13679 30141 13691 30175
rect 13633 30135 13691 30141
rect 15102 30132 15108 30184
rect 15160 30172 15166 30184
rect 15160 30144 15205 30172
rect 15160 30132 15166 30144
rect 15672 30104 15700 30212
rect 16226 30209 16238 30212
rect 16272 30240 16284 30243
rect 17126 30240 17132 30252
rect 16272 30212 17132 30240
rect 16272 30209 16284 30212
rect 16226 30203 16284 30209
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 17236 30240 17264 30280
rect 17773 30277 17785 30311
rect 17819 30308 17831 30311
rect 18138 30308 18144 30320
rect 17819 30280 18144 30308
rect 17819 30277 17831 30280
rect 17773 30271 17831 30277
rect 18138 30268 18144 30280
rect 18196 30268 18202 30320
rect 18984 30308 19012 30348
rect 20165 30345 20177 30379
rect 20211 30376 20223 30379
rect 20254 30376 20260 30388
rect 20211 30348 20260 30376
rect 20211 30345 20223 30348
rect 20165 30339 20223 30345
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 23658 30376 23664 30388
rect 20364 30348 23664 30376
rect 19518 30308 19524 30320
rect 18984 30280 19524 30308
rect 19518 30268 19524 30280
rect 19576 30268 19582 30320
rect 17862 30240 17868 30252
rect 17236 30212 17724 30240
rect 17823 30212 17868 30240
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 16117 30175 16175 30181
rect 16117 30141 16129 30175
rect 16163 30141 16175 30175
rect 16390 30172 16396 30184
rect 16351 30144 16396 30172
rect 16117 30135 16175 30141
rect 15212 30076 15700 30104
rect 9493 30039 9551 30045
rect 9493 30005 9505 30039
rect 9539 30036 9551 30039
rect 9582 30036 9588 30048
rect 9539 30008 9588 30036
rect 9539 30005 9551 30008
rect 9493 29999 9551 30005
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 11054 30036 11060 30048
rect 11015 30008 11060 30036
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 13078 30036 13084 30048
rect 13039 30008 13084 30036
rect 13078 29996 13084 30008
rect 13136 29996 13142 30048
rect 13354 29996 13360 30048
rect 13412 30036 13418 30048
rect 15212 30045 15240 30076
rect 15197 30039 15255 30045
rect 15197 30036 15209 30039
rect 13412 30008 15209 30036
rect 13412 29996 13418 30008
rect 15197 30005 15209 30008
rect 15243 30005 15255 30039
rect 15746 30036 15752 30048
rect 15707 30008 15752 30036
rect 15197 29999 15255 30005
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 15948 30036 15976 30135
rect 16132 30104 16160 30135
rect 16390 30132 16396 30144
rect 16448 30132 16454 30184
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 17313 30175 17371 30181
rect 17313 30172 17325 30175
rect 16632 30144 17325 30172
rect 16632 30132 16638 30144
rect 17313 30141 17325 30144
rect 17359 30141 17371 30175
rect 17494 30172 17500 30184
rect 17455 30144 17500 30172
rect 17313 30135 17371 30141
rect 17494 30132 17500 30144
rect 17552 30132 17558 30184
rect 17696 30172 17724 30212
rect 17862 30200 17868 30212
rect 17920 30200 17926 30252
rect 18785 30243 18843 30249
rect 18785 30240 18797 30243
rect 17963 30212 18797 30240
rect 17963 30172 17991 30212
rect 18785 30209 18797 30212
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 18506 30172 18512 30184
rect 17696 30144 17991 30172
rect 18467 30144 18512 30172
rect 18506 30132 18512 30144
rect 18564 30132 18570 30184
rect 18601 30175 18659 30181
rect 18601 30141 18613 30175
rect 18647 30172 18659 30175
rect 18690 30172 18696 30184
rect 18647 30144 18696 30172
rect 18647 30141 18659 30144
rect 18601 30135 18659 30141
rect 18690 30132 18696 30144
rect 18748 30132 18754 30184
rect 17862 30104 17868 30116
rect 16132 30076 17868 30104
rect 17862 30064 17868 30076
rect 17920 30064 17926 30116
rect 18800 30104 18828 30203
rect 18966 30200 18972 30252
rect 19024 30240 19030 30252
rect 19705 30243 19763 30249
rect 19705 30240 19717 30243
rect 19024 30212 19717 30240
rect 19024 30200 19030 30212
rect 19705 30209 19717 30212
rect 19751 30209 19763 30243
rect 19705 30203 19763 30209
rect 19797 30243 19855 30249
rect 19797 30209 19809 30243
rect 19843 30240 19855 30243
rect 19886 30240 19892 30252
rect 19843 30212 19892 30240
rect 19843 30209 19855 30212
rect 19797 30203 19855 30209
rect 19886 30200 19892 30212
rect 19944 30200 19950 30252
rect 20364 30240 20392 30348
rect 23658 30336 23664 30348
rect 23716 30336 23722 30388
rect 25498 30376 25504 30388
rect 25459 30348 25504 30376
rect 25498 30336 25504 30348
rect 25556 30336 25562 30388
rect 28445 30379 28503 30385
rect 28445 30345 28457 30379
rect 28491 30376 28503 30379
rect 31110 30376 31116 30388
rect 28491 30348 28856 30376
rect 28491 30345 28503 30348
rect 28445 30339 28503 30345
rect 20714 30268 20720 30320
rect 20772 30308 20778 30320
rect 20772 30280 20817 30308
rect 20772 30268 20778 30280
rect 20990 30268 20996 30320
rect 21048 30308 21054 30320
rect 21453 30311 21511 30317
rect 21453 30308 21465 30311
rect 21048 30280 21465 30308
rect 21048 30268 21054 30280
rect 21453 30277 21465 30280
rect 21499 30308 21511 30311
rect 22002 30308 22008 30320
rect 21499 30280 22008 30308
rect 21499 30277 21511 30280
rect 21453 30271 21511 30277
rect 22002 30268 22008 30280
rect 22060 30268 22066 30320
rect 24486 30268 24492 30320
rect 24544 30308 24550 30320
rect 24857 30311 24915 30317
rect 24857 30308 24869 30311
rect 24544 30280 24869 30308
rect 24544 30268 24550 30280
rect 24857 30277 24869 30280
rect 24903 30277 24915 30311
rect 24857 30271 24915 30277
rect 25961 30311 26019 30317
rect 25961 30277 25973 30311
rect 26007 30308 26019 30311
rect 26326 30308 26332 30320
rect 26007 30280 26332 30308
rect 26007 30277 26019 30280
rect 25961 30271 26019 30277
rect 26326 30268 26332 30280
rect 26384 30268 26390 30320
rect 26602 30268 26608 30320
rect 26660 30308 26666 30320
rect 26697 30311 26755 30317
rect 26697 30308 26709 30311
rect 26660 30280 26709 30308
rect 26660 30268 26666 30280
rect 26697 30277 26709 30280
rect 26743 30308 26755 30311
rect 26970 30308 26976 30320
rect 26743 30280 26976 30308
rect 26743 30277 26755 30280
rect 26697 30271 26755 30277
rect 26970 30268 26976 30280
rect 27028 30308 27034 30320
rect 28718 30308 28724 30320
rect 27028 30280 28724 30308
rect 27028 30268 27034 30280
rect 28718 30268 28724 30280
rect 28776 30268 28782 30320
rect 28828 30308 28856 30348
rect 28966 30348 29960 30376
rect 31071 30348 31116 30376
rect 28966 30308 28994 30348
rect 29822 30308 29828 30320
rect 28828 30280 28994 30308
rect 29783 30280 29828 30308
rect 29822 30268 29828 30280
rect 29880 30268 29886 30320
rect 29932 30308 29960 30348
rect 31110 30336 31116 30348
rect 31168 30336 31174 30388
rect 29932 30280 31708 30308
rect 27982 30240 27988 30252
rect 19996 30212 20392 30240
rect 26068 30212 27988 30240
rect 18874 30132 18880 30184
rect 18932 30172 18938 30184
rect 19429 30175 19487 30181
rect 18932 30144 18977 30172
rect 18932 30132 18938 30144
rect 19429 30141 19441 30175
rect 19475 30141 19487 30175
rect 19429 30135 19487 30141
rect 19334 30104 19340 30116
rect 18800 30076 19340 30104
rect 19334 30064 19340 30076
rect 19392 30064 19398 30116
rect 18874 30036 18880 30048
rect 15948 30008 18880 30036
rect 18874 29996 18880 30008
rect 18932 29996 18938 30048
rect 19444 30036 19472 30135
rect 19610 30132 19616 30184
rect 19668 30172 19674 30184
rect 19996 30181 20024 30212
rect 26068 30184 26096 30212
rect 27982 30200 27988 30212
rect 28040 30200 28046 30252
rect 30561 30243 30619 30249
rect 30561 30240 30573 30243
rect 28092 30212 30573 30240
rect 19981 30175 20039 30181
rect 19668 30144 19713 30172
rect 19668 30132 19674 30144
rect 19981 30141 19993 30175
rect 20027 30141 20039 30175
rect 19981 30135 20039 30141
rect 20625 30175 20683 30181
rect 20625 30141 20637 30175
rect 20671 30141 20683 30175
rect 20625 30135 20683 30141
rect 19518 30064 19524 30116
rect 19576 30104 19582 30116
rect 20640 30104 20668 30135
rect 20990 30132 20996 30184
rect 21048 30172 21054 30184
rect 21361 30175 21419 30181
rect 21361 30172 21373 30175
rect 21048 30144 21373 30172
rect 21048 30132 21054 30144
rect 21361 30141 21373 30144
rect 21407 30141 21419 30175
rect 21361 30135 21419 30141
rect 22278 30132 22284 30184
rect 22336 30172 22342 30184
rect 22833 30175 22891 30181
rect 22833 30172 22845 30175
rect 22336 30144 22845 30172
rect 22336 30132 22342 30144
rect 22833 30141 22845 30144
rect 22879 30172 22891 30175
rect 23198 30172 23204 30184
rect 22879 30144 23204 30172
rect 22879 30141 22891 30144
rect 22833 30135 22891 30141
rect 23198 30132 23204 30144
rect 23256 30132 23262 30184
rect 23477 30175 23535 30181
rect 23477 30141 23489 30175
rect 23523 30172 23535 30175
rect 23566 30172 23572 30184
rect 23523 30144 23572 30172
rect 23523 30141 23535 30144
rect 23477 30135 23535 30141
rect 23566 30132 23572 30144
rect 23624 30132 23630 30184
rect 23750 30181 23756 30184
rect 23744 30172 23756 30181
rect 23711 30144 23756 30172
rect 23744 30135 23756 30144
rect 23750 30132 23756 30135
rect 23808 30132 23814 30184
rect 25685 30175 25743 30181
rect 25685 30141 25697 30175
rect 25731 30141 25743 30175
rect 25685 30135 25743 30141
rect 19576 30076 20668 30104
rect 19576 30064 19582 30076
rect 22646 30064 22652 30116
rect 22704 30104 22710 30116
rect 24486 30104 24492 30116
rect 22704 30076 24492 30104
rect 22704 30064 22710 30076
rect 24486 30064 24492 30076
rect 24544 30064 24550 30116
rect 25700 30104 25728 30135
rect 25774 30132 25780 30184
rect 25832 30172 25838 30184
rect 26050 30172 26056 30184
rect 25832 30144 25877 30172
rect 25963 30144 26056 30172
rect 25832 30132 25838 30144
rect 26050 30132 26056 30144
rect 26108 30132 26114 30184
rect 26510 30132 26516 30184
rect 26568 30172 26574 30184
rect 26605 30175 26663 30181
rect 26605 30172 26617 30175
rect 26568 30144 26617 30172
rect 26568 30132 26574 30144
rect 26605 30141 26617 30144
rect 26651 30141 26663 30175
rect 26605 30135 26663 30141
rect 26694 30132 26700 30184
rect 26752 30172 26758 30184
rect 27793 30175 27851 30181
rect 27793 30172 27805 30175
rect 26752 30144 27805 30172
rect 26752 30132 26758 30144
rect 27793 30141 27805 30144
rect 27839 30141 27851 30175
rect 27793 30135 27851 30141
rect 26712 30104 26740 30132
rect 25700 30076 26740 30104
rect 27430 30064 27436 30116
rect 27488 30104 27494 30116
rect 28092 30104 28120 30212
rect 30561 30209 30573 30212
rect 30607 30209 30619 30243
rect 31680 30240 31708 30280
rect 31864 30280 36400 30308
rect 31864 30240 31892 30280
rect 31680 30212 31892 30240
rect 35452 30212 36216 30240
rect 30561 30203 30619 30209
rect 35452 30184 35480 30212
rect 28442 30132 28448 30184
rect 28500 30172 28506 30184
rect 28537 30175 28595 30181
rect 28537 30172 28549 30175
rect 28500 30144 28549 30172
rect 28500 30132 28506 30144
rect 28537 30141 28549 30144
rect 28583 30141 28595 30175
rect 28537 30135 28595 30141
rect 28626 30132 28632 30184
rect 28684 30172 28690 30184
rect 29181 30175 29239 30181
rect 29181 30172 29193 30175
rect 28684 30144 29193 30172
rect 28684 30132 28690 30144
rect 29181 30141 29193 30144
rect 29227 30141 29239 30175
rect 29822 30172 29828 30184
rect 29783 30144 29828 30172
rect 29181 30135 29239 30141
rect 29822 30132 29828 30144
rect 29880 30132 29886 30184
rect 30006 30132 30012 30184
rect 30064 30172 30070 30184
rect 30466 30172 30472 30184
rect 30064 30144 30109 30172
rect 30427 30144 30472 30172
rect 30064 30132 30070 30144
rect 30466 30132 30472 30144
rect 30524 30132 30530 30184
rect 30650 30172 30656 30184
rect 30611 30144 30656 30172
rect 30650 30132 30656 30144
rect 30708 30132 30714 30184
rect 31113 30175 31171 30181
rect 31113 30141 31125 30175
rect 31159 30141 31171 30175
rect 31113 30135 31171 30141
rect 31297 30175 31355 30181
rect 31297 30141 31309 30175
rect 31343 30172 31355 30175
rect 31478 30172 31484 30184
rect 31343 30144 31484 30172
rect 31343 30141 31355 30144
rect 31297 30135 31355 30141
rect 27488 30076 28120 30104
rect 27488 30064 27494 30076
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 29273 30107 29331 30113
rect 29273 30104 29285 30107
rect 28408 30076 29285 30104
rect 28408 30064 28414 30076
rect 29273 30073 29285 30076
rect 29319 30073 29331 30107
rect 30484 30104 30512 30132
rect 31128 30104 31156 30135
rect 31478 30132 31484 30144
rect 31536 30132 31542 30184
rect 35434 30172 35440 30184
rect 35395 30144 35440 30172
rect 35434 30132 35440 30144
rect 35492 30132 35498 30184
rect 36188 30181 36216 30212
rect 36372 30181 36400 30280
rect 50062 30268 50068 30320
rect 50120 30308 50126 30320
rect 55490 30308 55496 30320
rect 50120 30280 55496 30308
rect 50120 30268 50126 30280
rect 55490 30268 55496 30280
rect 55548 30268 55554 30320
rect 56870 30308 56876 30320
rect 55600 30280 56876 30308
rect 36538 30240 36544 30252
rect 36499 30212 36544 30240
rect 36538 30200 36544 30212
rect 36596 30200 36602 30252
rect 50154 30200 50160 30252
rect 50212 30240 50218 30252
rect 55600 30240 55628 30280
rect 56870 30268 56876 30280
rect 56928 30268 56934 30320
rect 57054 30308 57060 30320
rect 57015 30280 57060 30308
rect 57054 30268 57060 30280
rect 57112 30268 57118 30320
rect 50212 30212 55628 30240
rect 50212 30200 50218 30212
rect 55674 30200 55680 30252
rect 55732 30240 55738 30252
rect 57517 30243 57575 30249
rect 57517 30240 57529 30243
rect 55732 30212 57529 30240
rect 55732 30200 55738 30212
rect 57517 30209 57529 30212
rect 57563 30209 57575 30243
rect 57517 30203 57575 30209
rect 35529 30175 35587 30181
rect 35529 30141 35541 30175
rect 35575 30141 35587 30175
rect 35529 30135 35587 30141
rect 36173 30175 36231 30181
rect 36173 30141 36185 30175
rect 36219 30141 36231 30175
rect 36173 30135 36231 30141
rect 36357 30175 36415 30181
rect 36357 30141 36369 30175
rect 36403 30141 36415 30175
rect 36357 30135 36415 30141
rect 54757 30175 54815 30181
rect 54757 30141 54769 30175
rect 54803 30172 54815 30175
rect 54938 30172 54944 30184
rect 54803 30144 54944 30172
rect 54803 30141 54815 30144
rect 54757 30135 54815 30141
rect 35544 30104 35572 30135
rect 54938 30132 54944 30144
rect 54996 30132 55002 30184
rect 56134 30132 56140 30184
rect 56192 30172 56198 30184
rect 57701 30175 57759 30181
rect 57701 30172 57713 30175
rect 56192 30144 57713 30172
rect 56192 30132 56198 30144
rect 57701 30141 57713 30144
rect 57747 30141 57759 30175
rect 57701 30135 57759 30141
rect 30484 30076 31156 30104
rect 31726 30076 35572 30104
rect 35713 30107 35771 30113
rect 29273 30067 29331 30073
rect 22370 30036 22376 30048
rect 19444 30008 22376 30036
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 22738 29996 22744 30048
rect 22796 30036 22802 30048
rect 22925 30039 22983 30045
rect 22925 30036 22937 30039
rect 22796 30008 22937 30036
rect 22796 29996 22802 30008
rect 22925 30005 22937 30008
rect 22971 30036 22983 30039
rect 25406 30036 25412 30048
rect 22971 30008 25412 30036
rect 22971 30005 22983 30008
rect 22925 29999 22983 30005
rect 25406 29996 25412 30008
rect 25464 29996 25470 30048
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 27982 30036 27988 30048
rect 27939 30008 27988 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 27982 29996 27988 30008
rect 28040 29996 28046 30048
rect 28258 29996 28264 30048
rect 28316 30036 28322 30048
rect 28445 30039 28503 30045
rect 28445 30036 28457 30039
rect 28316 30008 28457 30036
rect 28316 29996 28322 30008
rect 28445 30005 28457 30008
rect 28491 30036 28503 30039
rect 28629 30039 28687 30045
rect 28629 30036 28641 30039
rect 28491 30008 28641 30036
rect 28491 30005 28503 30008
rect 28445 29999 28503 30005
rect 28629 30005 28641 30008
rect 28675 30005 28687 30039
rect 28629 29999 28687 30005
rect 28718 29996 28724 30048
rect 28776 30036 28782 30048
rect 30006 30036 30012 30048
rect 28776 30008 30012 30036
rect 28776 29996 28782 30008
rect 30006 29996 30012 30008
rect 30064 29996 30070 30048
rect 30098 29996 30104 30048
rect 30156 30036 30162 30048
rect 31726 30036 31754 30076
rect 35713 30073 35725 30107
rect 35759 30104 35771 30107
rect 55309 30107 55367 30113
rect 55309 30104 55321 30107
rect 35759 30076 55321 30104
rect 35759 30073 35771 30076
rect 35713 30067 35771 30073
rect 55309 30073 55321 30076
rect 55355 30073 55367 30107
rect 55309 30067 55367 30073
rect 55398 30064 55404 30116
rect 55456 30104 55462 30116
rect 55953 30107 56011 30113
rect 55456 30076 55501 30104
rect 55456 30064 55462 30076
rect 55953 30073 55965 30107
rect 55999 30104 56011 30107
rect 56873 30107 56931 30113
rect 55999 30076 56824 30104
rect 55999 30073 56011 30076
rect 55953 30067 56011 30073
rect 30156 30008 31754 30036
rect 54573 30039 54631 30045
rect 30156 29996 30162 30008
rect 54573 30005 54585 30039
rect 54619 30036 54631 30039
rect 56042 30036 56048 30048
rect 54619 30008 56048 30036
rect 54619 30005 54631 30008
rect 54573 29999 54631 30005
rect 56042 29996 56048 30008
rect 56100 29996 56106 30048
rect 56796 30036 56824 30076
rect 56873 30073 56885 30107
rect 56919 30104 56931 30107
rect 58161 30107 58219 30113
rect 58161 30104 58173 30107
rect 56919 30076 58173 30104
rect 56919 30073 56931 30076
rect 56873 30067 56931 30073
rect 58161 30073 58173 30076
rect 58207 30073 58219 30107
rect 58161 30067 58219 30073
rect 57514 30036 57520 30048
rect 56796 30008 57520 30036
rect 57514 29996 57520 30008
rect 57572 29996 57578 30048
rect 1104 29946 58880 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 50326 29946
rect 50378 29894 50390 29946
rect 50442 29894 50454 29946
rect 50506 29894 50518 29946
rect 50570 29894 58880 29946
rect 1104 29872 58880 29894
rect 11054 29792 11060 29844
rect 11112 29832 11118 29844
rect 15930 29832 15936 29844
rect 11112 29804 15936 29832
rect 11112 29792 11118 29804
rect 15930 29792 15936 29804
rect 15988 29792 15994 29844
rect 16117 29835 16175 29841
rect 16117 29801 16129 29835
rect 16163 29801 16175 29835
rect 16117 29795 16175 29801
rect 16669 29835 16727 29841
rect 16669 29801 16681 29835
rect 16715 29832 16727 29835
rect 17862 29832 17868 29844
rect 16715 29804 17868 29832
rect 16715 29801 16727 29804
rect 16669 29795 16727 29801
rect 12342 29764 12348 29776
rect 7300 29736 9720 29764
rect 12303 29736 12348 29764
rect 7300 29708 7328 29736
rect 1854 29696 1860 29708
rect 1815 29668 1860 29696
rect 1854 29656 1860 29668
rect 1912 29656 1918 29708
rect 6454 29696 6460 29708
rect 6415 29668 6460 29696
rect 6454 29656 6460 29668
rect 6512 29656 6518 29708
rect 7101 29699 7159 29705
rect 7101 29665 7113 29699
rect 7147 29696 7159 29699
rect 7190 29696 7196 29708
rect 7147 29668 7196 29696
rect 7147 29665 7159 29668
rect 7101 29659 7159 29665
rect 7190 29656 7196 29668
rect 7248 29656 7254 29708
rect 7282 29656 7288 29708
rect 7340 29696 7346 29708
rect 8113 29699 8171 29705
rect 7340 29668 7433 29696
rect 7340 29656 7346 29668
rect 8113 29665 8125 29699
rect 8159 29696 8171 29699
rect 8202 29696 8208 29708
rect 8159 29668 8208 29696
rect 8159 29665 8171 29668
rect 8113 29659 8171 29665
rect 8202 29656 8208 29668
rect 8260 29656 8266 29708
rect 9398 29656 9404 29708
rect 9456 29696 9462 29708
rect 9692 29705 9720 29736
rect 12342 29724 12348 29736
rect 12400 29724 12406 29776
rect 13648 29736 13952 29764
rect 9493 29699 9551 29705
rect 9493 29696 9505 29699
rect 9456 29668 9505 29696
rect 9456 29656 9462 29668
rect 9493 29665 9505 29668
rect 9539 29665 9551 29699
rect 9493 29659 9551 29665
rect 9677 29699 9735 29705
rect 9677 29665 9689 29699
rect 9723 29665 9735 29699
rect 9677 29659 9735 29665
rect 10772 29699 10830 29705
rect 10772 29665 10784 29699
rect 10818 29696 10830 29699
rect 11054 29696 11060 29708
rect 10818 29668 11060 29696
rect 10818 29665 10830 29668
rect 10772 29659 10830 29665
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 12526 29705 12532 29708
rect 12492 29699 12532 29705
rect 12492 29665 12504 29699
rect 12492 29659 12532 29665
rect 12526 29656 12532 29659
rect 12584 29656 12590 29708
rect 12802 29696 12808 29708
rect 12636 29668 12808 29696
rect 9582 29588 9588 29640
rect 9640 29628 9646 29640
rect 10505 29631 10563 29637
rect 10505 29628 10517 29631
rect 9640 29600 10517 29628
rect 9640 29588 9646 29600
rect 10505 29597 10517 29600
rect 10551 29597 10563 29631
rect 10505 29591 10563 29597
rect 12636 29572 12664 29668
rect 12802 29656 12808 29668
rect 12860 29656 12866 29708
rect 13648 29705 13676 29736
rect 13633 29699 13691 29705
rect 13633 29665 13645 29699
rect 13679 29665 13691 29699
rect 13633 29659 13691 29665
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29665 13875 29699
rect 13924 29696 13952 29736
rect 14734 29724 14740 29776
rect 14792 29764 14798 29776
rect 14982 29767 15040 29773
rect 14982 29764 14994 29767
rect 14792 29736 14994 29764
rect 14792 29724 14798 29736
rect 14982 29733 14994 29736
rect 15028 29733 15040 29767
rect 14982 29727 15040 29733
rect 15102 29724 15108 29776
rect 15160 29764 15166 29776
rect 16132 29764 16160 29795
rect 17862 29792 17868 29804
rect 17920 29792 17926 29844
rect 31570 29832 31576 29844
rect 17972 29804 31576 29832
rect 15160 29736 16620 29764
rect 15160 29724 15166 29736
rect 16592 29708 16620 29736
rect 16850 29724 16856 29776
rect 16908 29764 16914 29776
rect 17972 29773 18000 29804
rect 31570 29792 31576 29804
rect 31628 29792 31634 29844
rect 50154 29832 50160 29844
rect 31680 29804 50160 29832
rect 17957 29767 18015 29773
rect 16908 29736 17724 29764
rect 16908 29724 16914 29736
rect 17696 29708 17724 29736
rect 17957 29733 17969 29767
rect 18003 29733 18015 29767
rect 20073 29767 20131 29773
rect 20073 29764 20085 29767
rect 17957 29727 18015 29733
rect 18708 29736 20085 29764
rect 18708 29708 18736 29736
rect 20073 29733 20085 29736
rect 20119 29733 20131 29767
rect 20073 29727 20131 29733
rect 20898 29724 20904 29776
rect 20956 29764 20962 29776
rect 21146 29767 21204 29773
rect 21146 29764 21158 29767
rect 20956 29736 21158 29764
rect 20956 29724 20962 29736
rect 21146 29733 21158 29736
rect 21192 29733 21204 29767
rect 30736 29767 30794 29773
rect 21146 29727 21204 29733
rect 21264 29736 30696 29764
rect 15562 29696 15568 29708
rect 13924 29668 15568 29696
rect 13817 29659 13875 29665
rect 12713 29631 12771 29637
rect 12713 29597 12725 29631
rect 12759 29628 12771 29631
rect 12894 29628 12900 29640
rect 12759 29600 12900 29628
rect 12759 29597 12771 29600
rect 12713 29591 12771 29597
rect 12894 29588 12900 29600
rect 12952 29588 12958 29640
rect 13832 29628 13860 29659
rect 15562 29656 15568 29668
rect 15620 29696 15626 29708
rect 16390 29696 16396 29708
rect 15620 29668 16396 29696
rect 15620 29656 15626 29668
rect 16390 29656 16396 29668
rect 16448 29656 16454 29708
rect 16574 29696 16580 29708
rect 16535 29668 16580 29696
rect 16574 29656 16580 29668
rect 16632 29656 16638 29708
rect 16666 29656 16672 29708
rect 16724 29696 16730 29708
rect 16761 29699 16819 29705
rect 16761 29696 16773 29699
rect 16724 29668 16773 29696
rect 16724 29656 16730 29668
rect 16761 29665 16773 29668
rect 16807 29665 16819 29699
rect 17218 29696 17224 29708
rect 17179 29668 17224 29696
rect 16761 29659 16819 29665
rect 17218 29656 17224 29668
rect 17276 29656 17282 29708
rect 17678 29696 17684 29708
rect 17639 29668 17684 29696
rect 17678 29656 17684 29668
rect 17736 29656 17742 29708
rect 18598 29696 18604 29708
rect 18559 29668 18604 29696
rect 18598 29656 18604 29668
rect 18656 29656 18662 29708
rect 18690 29656 18696 29708
rect 18748 29696 18754 29708
rect 18877 29699 18935 29705
rect 18748 29668 18793 29696
rect 18748 29656 18754 29668
rect 18877 29665 18889 29699
rect 18923 29665 18935 29699
rect 18877 29659 18935 29665
rect 13998 29628 14004 29640
rect 13832 29600 14004 29628
rect 13998 29588 14004 29600
rect 14056 29588 14062 29640
rect 14366 29588 14372 29640
rect 14424 29628 14430 29640
rect 14737 29631 14795 29637
rect 14737 29628 14749 29631
rect 14424 29600 14749 29628
rect 14424 29588 14430 29600
rect 14737 29597 14749 29600
rect 14783 29597 14795 29631
rect 14737 29591 14795 29597
rect 15746 29588 15752 29640
rect 15804 29628 15810 29640
rect 18892 29628 18920 29659
rect 19150 29656 19156 29708
rect 19208 29696 19214 29708
rect 19981 29699 20039 29705
rect 19981 29696 19993 29699
rect 19208 29668 19993 29696
rect 19208 29656 19214 29668
rect 19981 29665 19993 29668
rect 20027 29665 20039 29699
rect 19981 29659 20039 29665
rect 20530 29656 20536 29708
rect 20588 29696 20594 29708
rect 21264 29696 21292 29736
rect 20588 29668 21292 29696
rect 20588 29656 20594 29668
rect 22646 29656 22652 29708
rect 22704 29696 22710 29708
rect 22741 29699 22799 29705
rect 22741 29696 22753 29699
rect 22704 29668 22753 29696
rect 22704 29656 22710 29668
rect 22741 29665 22753 29668
rect 22787 29665 22799 29699
rect 22741 29659 22799 29665
rect 22833 29699 22891 29705
rect 22833 29665 22845 29699
rect 22879 29696 22891 29699
rect 23474 29696 23480 29708
rect 22879 29668 23480 29696
rect 22879 29665 22891 29668
rect 22833 29659 22891 29665
rect 23474 29656 23480 29668
rect 23532 29696 23538 29708
rect 23845 29699 23903 29705
rect 23845 29696 23857 29699
rect 23532 29668 23857 29696
rect 23532 29656 23538 29668
rect 23845 29665 23857 29668
rect 23891 29665 23903 29699
rect 23845 29659 23903 29665
rect 24029 29699 24087 29705
rect 24029 29665 24041 29699
rect 24075 29696 24087 29699
rect 25038 29696 25044 29708
rect 24075 29668 25044 29696
rect 24075 29665 24087 29668
rect 24029 29659 24087 29665
rect 25038 29656 25044 29668
rect 25096 29656 25102 29708
rect 25225 29699 25283 29705
rect 25225 29665 25237 29699
rect 25271 29665 25283 29699
rect 25225 29659 25283 29665
rect 15804 29600 18920 29628
rect 15804 29588 15810 29600
rect 20070 29588 20076 29640
rect 20128 29628 20134 29640
rect 20901 29631 20959 29637
rect 20901 29628 20913 29631
rect 20128 29600 20913 29628
rect 20128 29588 20134 29600
rect 20901 29597 20913 29600
rect 20947 29597 20959 29631
rect 20901 29591 20959 29597
rect 22922 29588 22928 29640
rect 22980 29628 22986 29640
rect 23017 29631 23075 29637
rect 23017 29628 23029 29631
rect 22980 29600 23029 29628
rect 22980 29588 22986 29600
rect 23017 29597 23029 29600
rect 23063 29628 23075 29631
rect 23934 29628 23940 29640
rect 23063 29600 23940 29628
rect 23063 29597 23075 29600
rect 23017 29591 23075 29597
rect 23934 29588 23940 29600
rect 23992 29588 23998 29640
rect 24305 29631 24363 29637
rect 24305 29597 24317 29631
rect 24351 29628 24363 29631
rect 24946 29628 24952 29640
rect 24351 29600 24952 29628
rect 24351 29597 24363 29600
rect 24305 29591 24363 29597
rect 24946 29588 24952 29600
rect 25004 29588 25010 29640
rect 12618 29560 12624 29572
rect 12531 29532 12624 29560
rect 12618 29520 12624 29532
rect 12676 29520 12682 29572
rect 18506 29520 18512 29572
rect 18564 29560 18570 29572
rect 18785 29563 18843 29569
rect 18785 29560 18797 29563
rect 18564 29532 18797 29560
rect 18564 29520 18570 29532
rect 18785 29529 18797 29532
rect 18831 29560 18843 29563
rect 19426 29560 19432 29572
rect 18831 29532 19432 29560
rect 18831 29529 18843 29532
rect 18785 29523 18843 29529
rect 19426 29520 19432 29532
rect 19484 29520 19490 29572
rect 22278 29560 22284 29572
rect 22239 29532 22284 29560
rect 22278 29520 22284 29532
rect 22336 29520 22342 29572
rect 22646 29520 22652 29572
rect 22704 29560 22710 29572
rect 25240 29560 25268 29659
rect 26234 29656 26240 29708
rect 26292 29696 26298 29708
rect 26329 29699 26387 29705
rect 26329 29696 26341 29699
rect 26292 29668 26341 29696
rect 26292 29656 26298 29668
rect 26329 29665 26341 29668
rect 26375 29665 26387 29699
rect 26329 29659 26387 29665
rect 22704 29532 25268 29560
rect 26344 29560 26372 29659
rect 26418 29656 26424 29708
rect 26476 29696 26482 29708
rect 26602 29696 26608 29708
rect 26476 29668 26521 29696
rect 26563 29668 26608 29696
rect 26476 29656 26482 29668
rect 26602 29656 26608 29668
rect 26660 29656 26666 29708
rect 26694 29656 26700 29708
rect 26752 29696 26758 29708
rect 27341 29699 27399 29705
rect 26752 29668 26797 29696
rect 26752 29656 26758 29668
rect 27341 29665 27353 29699
rect 27387 29696 27399 29699
rect 27798 29696 27804 29708
rect 27387 29668 27804 29696
rect 27387 29665 27399 29668
rect 27341 29659 27399 29665
rect 27798 29656 27804 29668
rect 27856 29696 27862 29708
rect 27985 29699 28043 29705
rect 27985 29696 27997 29699
rect 27856 29668 27997 29696
rect 27856 29656 27862 29668
rect 27985 29665 27997 29668
rect 28031 29665 28043 29699
rect 28166 29696 28172 29708
rect 28079 29668 28172 29696
rect 27985 29659 28043 29665
rect 26436 29628 26464 29656
rect 28092 29628 28120 29668
rect 28166 29656 28172 29668
rect 28224 29656 28230 29708
rect 28258 29656 28264 29708
rect 28316 29696 28322 29708
rect 28537 29699 28595 29705
rect 28316 29668 28409 29696
rect 28316 29656 28322 29668
rect 28537 29665 28549 29699
rect 28583 29696 28595 29699
rect 28810 29696 28816 29708
rect 28583 29668 28816 29696
rect 28583 29665 28595 29668
rect 28537 29659 28595 29665
rect 28810 29656 28816 29668
rect 28868 29696 28874 29708
rect 28997 29699 29055 29705
rect 28997 29696 29009 29699
rect 28868 29668 29009 29696
rect 28868 29656 28874 29668
rect 28997 29665 29009 29668
rect 29043 29665 29055 29699
rect 30668 29696 30696 29736
rect 30736 29733 30748 29767
rect 30782 29764 30794 29767
rect 31110 29764 31116 29776
rect 30782 29736 31116 29764
rect 30782 29733 30794 29736
rect 30736 29727 30794 29733
rect 31110 29724 31116 29736
rect 31168 29724 31174 29776
rect 31680 29696 31708 29804
rect 50154 29792 50160 29804
rect 50212 29792 50218 29844
rect 54389 29835 54447 29841
rect 54389 29801 54401 29835
rect 54435 29832 54447 29835
rect 55398 29832 55404 29844
rect 54435 29804 55404 29832
rect 54435 29801 54447 29804
rect 54389 29795 54447 29801
rect 55398 29792 55404 29804
rect 55456 29792 55462 29844
rect 58618 29832 58624 29844
rect 55784 29804 58624 29832
rect 31754 29724 31760 29776
rect 31812 29764 31818 29776
rect 50062 29764 50068 29776
rect 31812 29736 50068 29764
rect 31812 29724 31818 29736
rect 50062 29724 50068 29736
rect 50120 29724 50126 29776
rect 54846 29724 54852 29776
rect 54904 29764 54910 29776
rect 55784 29773 55812 29804
rect 58618 29792 58624 29804
rect 58676 29792 58682 29844
rect 55217 29767 55275 29773
rect 55217 29764 55229 29767
rect 54904 29736 55229 29764
rect 54904 29724 54910 29736
rect 55217 29733 55229 29736
rect 55263 29733 55275 29767
rect 55217 29727 55275 29733
rect 55769 29767 55827 29773
rect 55769 29733 55781 29767
rect 55815 29733 55827 29767
rect 55769 29727 55827 29733
rect 56042 29724 56048 29776
rect 56100 29764 56106 29776
rect 56873 29767 56931 29773
rect 56873 29764 56885 29767
rect 56100 29736 56885 29764
rect 56100 29724 56106 29736
rect 56873 29733 56885 29736
rect 56919 29733 56931 29767
rect 56873 29727 56931 29733
rect 57425 29767 57483 29773
rect 57425 29733 57437 29767
rect 57471 29764 57483 29767
rect 57698 29764 57704 29776
rect 57471 29736 57704 29764
rect 57471 29733 57483 29736
rect 57425 29727 57483 29733
rect 57698 29724 57704 29736
rect 57756 29724 57762 29776
rect 30668 29668 31708 29696
rect 32309 29699 32367 29705
rect 28997 29659 29055 29665
rect 32309 29665 32321 29699
rect 32355 29665 32367 29699
rect 32309 29659 32367 29665
rect 53745 29699 53803 29705
rect 53745 29665 53757 29699
rect 53791 29696 53803 29699
rect 54478 29696 54484 29708
rect 53791 29668 54484 29696
rect 53791 29665 53803 29668
rect 53745 29659 53803 29665
rect 28276 29628 28304 29656
rect 28442 29628 28448 29640
rect 26436 29600 28120 29628
rect 28184 29600 28304 29628
rect 28403 29600 28448 29628
rect 28184 29560 28212 29600
rect 28442 29588 28448 29600
rect 28500 29588 28506 29640
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 30469 29631 30527 29637
rect 30469 29628 30481 29631
rect 30432 29600 30481 29628
rect 30432 29588 30438 29600
rect 30469 29597 30481 29600
rect 30515 29597 30527 29631
rect 30469 29591 30527 29597
rect 26344 29532 28212 29560
rect 22704 29520 22710 29532
rect 28258 29520 28264 29572
rect 28316 29560 28322 29572
rect 29089 29563 29147 29569
rect 29089 29560 29101 29563
rect 28316 29532 29101 29560
rect 28316 29520 28322 29532
rect 29089 29529 29101 29532
rect 29135 29529 29147 29563
rect 29089 29523 29147 29529
rect 31570 29520 31576 29572
rect 31628 29560 31634 29572
rect 31849 29563 31907 29569
rect 31849 29560 31861 29563
rect 31628 29532 31861 29560
rect 31628 29520 31634 29532
rect 31849 29529 31861 29532
rect 31895 29560 31907 29563
rect 32324 29560 32352 29659
rect 54478 29656 54484 29668
rect 54536 29656 54542 29708
rect 54573 29699 54631 29705
rect 54573 29665 54585 29699
rect 54619 29696 54631 29699
rect 54938 29696 54944 29708
rect 54619 29668 54944 29696
rect 54619 29665 54631 29668
rect 54573 29659 54631 29665
rect 54938 29656 54944 29668
rect 54996 29656 55002 29708
rect 57974 29696 57980 29708
rect 57935 29668 57980 29696
rect 57974 29656 57980 29668
rect 58032 29656 58038 29708
rect 50246 29588 50252 29640
rect 50304 29628 50310 29640
rect 55125 29631 55183 29637
rect 55125 29628 55137 29631
rect 50304 29600 55137 29628
rect 50304 29588 50310 29600
rect 55125 29597 55137 29600
rect 55171 29597 55183 29631
rect 56781 29631 56839 29637
rect 56781 29628 56793 29631
rect 55125 29591 55183 29597
rect 55600 29600 56793 29628
rect 31895 29532 32352 29560
rect 31895 29529 31907 29532
rect 31849 29523 31907 29529
rect 50338 29520 50344 29572
rect 50396 29560 50402 29572
rect 55600 29560 55628 29600
rect 56781 29597 56793 29600
rect 56827 29597 56839 29631
rect 56781 29591 56839 29597
rect 58158 29560 58164 29572
rect 50396 29532 55628 29560
rect 58119 29532 58164 29560
rect 50396 29520 50402 29532
rect 58158 29520 58164 29532
rect 58216 29520 58222 29572
rect 1946 29492 1952 29504
rect 1907 29464 1952 29492
rect 1946 29452 1952 29464
rect 2004 29452 2010 29504
rect 6546 29492 6552 29504
rect 6507 29464 6552 29492
rect 6546 29452 6552 29464
rect 6604 29452 6610 29504
rect 7098 29492 7104 29504
rect 7059 29464 7104 29492
rect 7098 29452 7104 29464
rect 7156 29452 7162 29504
rect 8110 29452 8116 29504
rect 8168 29492 8174 29504
rect 8205 29495 8263 29501
rect 8205 29492 8217 29495
rect 8168 29464 8217 29492
rect 8168 29452 8174 29464
rect 8205 29461 8217 29464
rect 8251 29461 8263 29495
rect 9490 29492 9496 29504
rect 9451 29464 9496 29492
rect 8205 29455 8263 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 11885 29495 11943 29501
rect 11885 29461 11897 29495
rect 11931 29492 11943 29495
rect 12066 29492 12072 29504
rect 11931 29464 12072 29492
rect 11931 29461 11943 29464
rect 11885 29455 11943 29461
rect 12066 29452 12072 29464
rect 12124 29452 12130 29504
rect 12989 29495 13047 29501
rect 12989 29461 13001 29495
rect 13035 29492 13047 29495
rect 13538 29492 13544 29504
rect 13035 29464 13544 29492
rect 13035 29461 13047 29464
rect 12989 29455 13047 29461
rect 13538 29452 13544 29464
rect 13596 29452 13602 29504
rect 13633 29495 13691 29501
rect 13633 29461 13645 29495
rect 13679 29492 13691 29495
rect 14734 29492 14740 29504
rect 13679 29464 14740 29492
rect 13679 29461 13691 29464
rect 13633 29455 13691 29461
rect 14734 29452 14740 29464
rect 14792 29452 14798 29504
rect 17310 29452 17316 29504
rect 17368 29492 17374 29504
rect 18417 29495 18475 29501
rect 18417 29492 18429 29495
rect 17368 29464 18429 29492
rect 17368 29452 17374 29464
rect 18417 29461 18429 29464
rect 18463 29461 18475 29495
rect 18417 29455 18475 29461
rect 18598 29452 18604 29504
rect 18656 29492 18662 29504
rect 21082 29492 21088 29504
rect 18656 29464 21088 29492
rect 18656 29452 18662 29464
rect 21082 29452 21088 29464
rect 21140 29452 21146 29504
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22888 29464 22937 29492
rect 22888 29452 22894 29464
rect 22925 29461 22937 29464
rect 22971 29492 22983 29495
rect 24026 29492 24032 29504
rect 22971 29464 24032 29492
rect 22971 29461 22983 29464
rect 22925 29455 22983 29461
rect 24026 29452 24032 29464
rect 24084 29452 24090 29504
rect 24213 29495 24271 29501
rect 24213 29461 24225 29495
rect 24259 29492 24271 29495
rect 24854 29492 24860 29504
rect 24259 29464 24860 29492
rect 24259 29461 24271 29464
rect 24213 29455 24271 29461
rect 24854 29452 24860 29464
rect 24912 29452 24918 29504
rect 25314 29492 25320 29504
rect 25275 29464 25320 29492
rect 25314 29452 25320 29464
rect 25372 29452 25378 29504
rect 25866 29452 25872 29504
rect 25924 29492 25930 29504
rect 26145 29495 26203 29501
rect 26145 29492 26157 29495
rect 25924 29464 26157 29492
rect 25924 29452 25930 29464
rect 26145 29461 26157 29464
rect 26191 29461 26203 29495
rect 26145 29455 26203 29461
rect 27338 29452 27344 29504
rect 27396 29492 27402 29504
rect 27433 29495 27491 29501
rect 27433 29492 27445 29495
rect 27396 29464 27445 29492
rect 27396 29452 27402 29464
rect 27433 29461 27445 29464
rect 27479 29461 27491 29495
rect 27433 29455 27491 29461
rect 28074 29452 28080 29504
rect 28132 29492 28138 29504
rect 30650 29492 30656 29504
rect 28132 29464 30656 29492
rect 28132 29452 28138 29464
rect 30650 29452 30656 29464
rect 30708 29452 30714 29504
rect 31754 29452 31760 29504
rect 31812 29492 31818 29504
rect 32401 29495 32459 29501
rect 32401 29492 32413 29495
rect 31812 29464 32413 29492
rect 31812 29452 31818 29464
rect 32401 29461 32413 29464
rect 32447 29492 32459 29495
rect 35618 29492 35624 29504
rect 32447 29464 35624 29492
rect 32447 29461 32459 29464
rect 32401 29455 32459 29461
rect 35618 29452 35624 29464
rect 35676 29452 35682 29504
rect 54478 29452 54484 29504
rect 54536 29492 54542 29504
rect 56502 29492 56508 29504
rect 54536 29464 56508 29492
rect 54536 29452 54542 29464
rect 56502 29452 56508 29464
rect 56560 29452 56566 29504
rect 1104 29402 58880 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 58880 29402
rect 1104 29328 58880 29350
rect 8202 29288 8208 29300
rect 8163 29260 8208 29288
rect 8202 29248 8208 29260
rect 8260 29248 8266 29300
rect 11514 29248 11520 29300
rect 11572 29288 11578 29300
rect 12161 29291 12219 29297
rect 12161 29288 12173 29291
rect 11572 29260 12173 29288
rect 11572 29248 11578 29260
rect 12161 29257 12173 29260
rect 12207 29257 12219 29291
rect 12161 29251 12219 29257
rect 12250 29248 12256 29300
rect 12308 29288 12314 29300
rect 13173 29291 13231 29297
rect 13173 29288 13185 29291
rect 12308 29260 13185 29288
rect 12308 29248 12314 29260
rect 13173 29257 13185 29260
rect 13219 29257 13231 29291
rect 13173 29251 13231 29257
rect 15930 29248 15936 29300
rect 15988 29288 15994 29300
rect 18506 29288 18512 29300
rect 15988 29260 18512 29288
rect 15988 29248 15994 29260
rect 18506 29248 18512 29260
rect 18564 29248 18570 29300
rect 18877 29291 18935 29297
rect 18877 29257 18889 29291
rect 18923 29288 18935 29291
rect 18966 29288 18972 29300
rect 18923 29260 18972 29288
rect 18923 29257 18935 29260
rect 18877 29251 18935 29257
rect 18966 29248 18972 29260
rect 19024 29248 19030 29300
rect 20438 29288 20444 29300
rect 20399 29260 20444 29288
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 21082 29288 21088 29300
rect 20732 29260 21088 29288
rect 10137 29223 10195 29229
rect 10137 29189 10149 29223
rect 10183 29189 10195 29223
rect 10137 29183 10195 29189
rect 8754 29152 8760 29164
rect 5920 29124 6960 29152
rect 8715 29124 8760 29152
rect 1857 29087 1915 29093
rect 1857 29053 1869 29087
rect 1903 29084 1915 29087
rect 2958 29084 2964 29096
rect 1903 29056 2964 29084
rect 1903 29053 1915 29056
rect 1857 29047 1915 29053
rect 2958 29044 2964 29056
rect 3016 29044 3022 29096
rect 5920 29093 5948 29124
rect 5721 29087 5779 29093
rect 5721 29053 5733 29087
rect 5767 29053 5779 29087
rect 5721 29047 5779 29053
rect 5905 29087 5963 29093
rect 5905 29053 5917 29087
rect 5951 29053 5963 29087
rect 6822 29084 6828 29096
rect 6783 29056 6828 29084
rect 5905 29047 5963 29053
rect 2038 29016 2044 29028
rect 1999 28988 2044 29016
rect 2038 28976 2044 28988
rect 2096 28976 2102 29028
rect 5736 29016 5764 29047
rect 6822 29044 6828 29056
rect 6880 29044 6886 29096
rect 6932 29084 6960 29124
rect 8754 29112 8760 29124
rect 8812 29112 8818 29164
rect 7098 29093 7104 29096
rect 6932 29056 7052 29084
rect 6914 29016 6920 29028
rect 5736 28988 6920 29016
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7024 29016 7052 29056
rect 7092 29047 7104 29093
rect 7156 29084 7162 29096
rect 9024 29087 9082 29093
rect 7156 29056 7192 29084
rect 7098 29044 7104 29047
rect 7156 29044 7162 29056
rect 9024 29053 9036 29087
rect 9070 29084 9082 29087
rect 9490 29084 9496 29096
rect 9070 29056 9496 29084
rect 9070 29053 9082 29056
rect 9024 29047 9082 29053
rect 9490 29044 9496 29056
rect 9548 29044 9554 29096
rect 10152 29084 10180 29183
rect 12986 29180 12992 29232
rect 13044 29220 13050 29232
rect 15105 29223 15163 29229
rect 13044 29192 15056 29220
rect 13044 29180 13050 29192
rect 11146 29112 11152 29164
rect 11204 29152 11210 29164
rect 13541 29155 13599 29161
rect 13541 29152 13553 29155
rect 11204 29124 13553 29152
rect 11204 29112 11210 29124
rect 13541 29121 13553 29124
rect 13587 29121 13599 29155
rect 15028 29152 15056 29192
rect 15105 29189 15117 29223
rect 15151 29220 15163 29223
rect 15286 29220 15292 29232
rect 15151 29192 15292 29220
rect 15151 29189 15163 29192
rect 15105 29183 15163 29189
rect 15286 29180 15292 29192
rect 15344 29180 15350 29232
rect 18690 29180 18696 29232
rect 18748 29220 18754 29232
rect 19337 29223 19395 29229
rect 19337 29220 19349 29223
rect 18748 29192 19349 29220
rect 18748 29180 18754 29192
rect 19337 29189 19349 29192
rect 19383 29189 19395 29223
rect 19337 29183 19395 29189
rect 15304 29152 15332 29180
rect 16393 29155 16451 29161
rect 15028 29124 15240 29152
rect 15304 29124 16160 29152
rect 13541 29115 13599 29121
rect 10597 29087 10655 29093
rect 10597 29084 10609 29087
rect 10152 29056 10609 29084
rect 10597 29053 10609 29056
rect 10643 29053 10655 29087
rect 12066 29084 12072 29096
rect 12027 29056 12072 29084
rect 10597 29047 10655 29053
rect 12066 29044 12072 29056
rect 12124 29044 12130 29096
rect 13078 29084 13084 29096
rect 13039 29056 13084 29084
rect 13078 29044 13084 29056
rect 13136 29084 13142 29096
rect 14277 29087 14335 29093
rect 14277 29084 14289 29087
rect 13136 29056 14289 29084
rect 13136 29044 13142 29056
rect 14277 29053 14289 29056
rect 14323 29053 14335 29087
rect 14277 29047 14335 29053
rect 15013 29087 15071 29093
rect 15013 29053 15025 29087
rect 15059 29084 15071 29087
rect 15102 29084 15108 29096
rect 15059 29056 15108 29084
rect 15059 29053 15071 29056
rect 15013 29047 15071 29053
rect 15102 29044 15108 29056
rect 15160 29044 15166 29096
rect 15212 29084 15240 29124
rect 16132 29093 16160 29124
rect 16393 29121 16405 29155
rect 16439 29152 16451 29155
rect 20530 29152 20536 29164
rect 16439 29124 20536 29152
rect 16439 29121 16451 29124
rect 16393 29115 16451 29121
rect 20530 29112 20536 29124
rect 20588 29112 20594 29164
rect 15657 29087 15715 29093
rect 15657 29084 15669 29087
rect 15212 29056 15669 29084
rect 15657 29053 15669 29056
rect 15703 29053 15715 29087
rect 15657 29047 15715 29053
rect 16117 29087 16175 29093
rect 16117 29053 16129 29087
rect 16163 29053 16175 29087
rect 17218 29084 17224 29096
rect 16117 29047 16175 29053
rect 17052 29056 17224 29084
rect 7282 29016 7288 29028
rect 7024 28988 7288 29016
rect 7282 28976 7288 28988
rect 7340 28976 7346 29028
rect 13814 28976 13820 29028
rect 13872 29016 13878 29028
rect 14093 29019 14151 29025
rect 14093 29016 14105 29019
rect 13872 28988 14105 29016
rect 13872 28976 13878 28988
rect 14093 28985 14105 28988
rect 14139 28985 14151 29019
rect 14458 29016 14464 29028
rect 14419 28988 14464 29016
rect 14093 28979 14151 28985
rect 14458 28976 14464 28988
rect 14516 28976 14522 29028
rect 15672 29016 15700 29047
rect 17052 29016 17080 29056
rect 17218 29044 17224 29056
rect 17276 29084 17282 29096
rect 17313 29087 17371 29093
rect 17313 29084 17325 29087
rect 17276 29056 17325 29084
rect 17276 29044 17282 29056
rect 17313 29053 17325 29056
rect 17359 29053 17371 29087
rect 17313 29047 17371 29053
rect 17773 29087 17831 29093
rect 17773 29053 17785 29087
rect 17819 29053 17831 29087
rect 17773 29047 17831 29053
rect 19061 29087 19119 29093
rect 19061 29053 19073 29087
rect 19107 29053 19119 29087
rect 19061 29047 19119 29053
rect 15672 28988 17080 29016
rect 17126 28976 17132 29028
rect 17184 29016 17190 29028
rect 17788 29016 17816 29047
rect 18046 29016 18052 29028
rect 17184 28988 17816 29016
rect 18007 28988 18052 29016
rect 17184 28976 17190 28988
rect 18046 28976 18052 28988
rect 18104 28976 18110 29028
rect 19076 29016 19104 29047
rect 19150 29044 19156 29096
rect 19208 29084 19214 29096
rect 19426 29084 19432 29096
rect 19208 29056 19253 29084
rect 19387 29056 19432 29084
rect 19208 29044 19214 29056
rect 19426 29044 19432 29056
rect 19484 29044 19490 29096
rect 20732 29093 20760 29260
rect 21082 29248 21088 29260
rect 21140 29248 21146 29300
rect 21818 29248 21824 29300
rect 21876 29288 21882 29300
rect 22554 29288 22560 29300
rect 21876 29260 22560 29288
rect 21876 29248 21882 29260
rect 22554 29248 22560 29260
rect 22612 29248 22618 29300
rect 24397 29291 24455 29297
rect 24397 29288 24409 29291
rect 22664 29260 24409 29288
rect 20898 29220 20904 29232
rect 20824 29192 20904 29220
rect 20824 29093 20852 29192
rect 20898 29180 20904 29192
rect 20956 29180 20962 29232
rect 22664 29164 22692 29260
rect 24397 29257 24409 29260
rect 24443 29257 24455 29291
rect 24397 29251 24455 29257
rect 24578 29248 24584 29300
rect 24636 29288 24642 29300
rect 25041 29291 25099 29297
rect 25041 29288 25053 29291
rect 24636 29260 25053 29288
rect 24636 29248 24642 29260
rect 25041 29257 25053 29260
rect 25087 29257 25099 29291
rect 25041 29251 25099 29257
rect 27801 29291 27859 29297
rect 27801 29257 27813 29291
rect 27847 29288 27859 29291
rect 27890 29288 27896 29300
rect 27847 29260 27896 29288
rect 27847 29257 27859 29260
rect 27801 29251 27859 29257
rect 27890 29248 27896 29260
rect 27948 29288 27954 29300
rect 28626 29288 28632 29300
rect 27948 29260 28632 29288
rect 27948 29248 27954 29260
rect 28626 29248 28632 29260
rect 28684 29248 28690 29300
rect 28810 29248 28816 29300
rect 28868 29288 28874 29300
rect 30193 29291 30251 29297
rect 30193 29288 30205 29291
rect 28868 29260 30205 29288
rect 28868 29248 28874 29260
rect 30193 29257 30205 29260
rect 30239 29257 30251 29291
rect 50338 29288 50344 29300
rect 30193 29251 30251 29257
rect 35728 29260 50344 29288
rect 22995 29223 23053 29229
rect 22995 29189 23007 29223
rect 23041 29220 23053 29223
rect 24213 29223 24271 29229
rect 23041 29192 24164 29220
rect 23041 29189 23053 29192
rect 22995 29183 23053 29189
rect 22646 29112 22652 29164
rect 22704 29112 22710 29164
rect 23106 29152 23112 29164
rect 23067 29124 23112 29152
rect 23106 29112 23112 29124
rect 23164 29112 23170 29164
rect 23198 29112 23204 29164
rect 23256 29152 23262 29164
rect 23256 29124 23301 29152
rect 23256 29112 23262 29124
rect 20697 29087 20760 29093
rect 20697 29053 20709 29087
rect 20743 29056 20760 29087
rect 20806 29087 20864 29093
rect 20743 29053 20755 29056
rect 20697 29047 20755 29053
rect 20806 29053 20818 29087
rect 20852 29053 20864 29087
rect 20806 29047 20864 29053
rect 20898 29044 20904 29096
rect 20956 29084 20962 29096
rect 21082 29084 21088 29096
rect 20956 29056 21001 29084
rect 21043 29056 21088 29084
rect 20956 29044 20962 29056
rect 21082 29044 21088 29056
rect 21140 29044 21146 29096
rect 23290 29084 23296 29096
rect 23251 29056 23296 29084
rect 23290 29044 23296 29056
rect 23348 29044 23354 29096
rect 24136 29093 24164 29192
rect 24213 29189 24225 29223
rect 24259 29220 24271 29223
rect 24946 29220 24952 29232
rect 24259 29192 24952 29220
rect 24259 29189 24271 29192
rect 24213 29183 24271 29189
rect 24946 29180 24952 29192
rect 25004 29220 25010 29232
rect 25774 29220 25780 29232
rect 25004 29192 25780 29220
rect 25004 29180 25010 29192
rect 25774 29180 25780 29192
rect 25832 29180 25838 29232
rect 26326 29180 26332 29232
rect 26384 29220 26390 29232
rect 27522 29220 27528 29232
rect 26384 29192 27528 29220
rect 26384 29180 26390 29192
rect 27522 29180 27528 29192
rect 27580 29220 27586 29232
rect 33318 29220 33324 29232
rect 27580 29192 28028 29220
rect 27580 29180 27586 29192
rect 24305 29155 24363 29161
rect 24305 29121 24317 29155
rect 24351 29152 24363 29155
rect 24854 29152 24860 29164
rect 24351 29124 24860 29152
rect 24351 29121 24363 29124
rect 24305 29115 24363 29121
rect 24854 29112 24860 29124
rect 24912 29112 24918 29164
rect 26605 29155 26663 29161
rect 26605 29152 26617 29155
rect 25062 29124 26617 29152
rect 25062 29096 25090 29124
rect 26605 29121 26617 29124
rect 26651 29121 26663 29155
rect 28000 29152 28028 29192
rect 33305 29180 33324 29220
rect 33376 29180 33382 29232
rect 35728 29229 35756 29260
rect 50338 29248 50344 29260
rect 50396 29248 50402 29300
rect 54846 29288 54852 29300
rect 54807 29260 54852 29288
rect 54846 29248 54852 29260
rect 54904 29248 54910 29300
rect 56134 29288 56140 29300
rect 56095 29260 56140 29288
rect 56134 29248 56140 29260
rect 56192 29248 56198 29300
rect 57974 29288 57980 29300
rect 57935 29260 57980 29288
rect 57974 29248 57980 29260
rect 58032 29248 58038 29300
rect 35713 29223 35771 29229
rect 35713 29189 35725 29223
rect 35759 29189 35771 29223
rect 35713 29183 35771 29189
rect 55214 29180 55220 29232
rect 55272 29220 55278 29232
rect 55677 29223 55735 29229
rect 55677 29220 55689 29223
rect 55272 29192 55689 29220
rect 55272 29180 55278 29192
rect 55677 29189 55689 29192
rect 55723 29189 55735 29223
rect 55677 29183 55735 29189
rect 57057 29223 57115 29229
rect 57057 29189 57069 29223
rect 57103 29220 57115 29223
rect 57146 29220 57152 29232
rect 57103 29192 57152 29220
rect 57103 29189 57115 29192
rect 57057 29183 57115 29189
rect 57146 29180 57152 29192
rect 57204 29180 57210 29232
rect 28261 29155 28319 29161
rect 28261 29152 28273 29155
rect 28000 29124 28120 29152
rect 26605 29115 26663 29121
rect 24121 29087 24179 29093
rect 24121 29053 24133 29087
rect 24167 29053 24179 29087
rect 24486 29084 24492 29096
rect 24447 29056 24492 29084
rect 24121 29047 24179 29053
rect 24486 29044 24492 29056
rect 24544 29084 24550 29096
rect 24544 29056 24992 29084
rect 24544 29044 24550 29056
rect 20530 29016 20536 29028
rect 19076 28988 20536 29016
rect 20530 28976 20536 28988
rect 20588 28976 20594 29028
rect 21266 28976 21272 29028
rect 21324 29016 21330 29028
rect 22646 29016 22652 29028
rect 21324 28988 22652 29016
rect 21324 28976 21330 28988
rect 22646 28976 22652 28988
rect 22704 28976 22710 29028
rect 22922 29016 22928 29028
rect 22883 28988 22928 29016
rect 22922 28976 22928 28988
rect 22980 28976 22986 29028
rect 23474 28976 23480 29028
rect 23532 28976 23538 29028
rect 23750 28976 23756 29028
rect 23808 29016 23814 29028
rect 24578 29016 24584 29028
rect 23808 28988 24584 29016
rect 23808 28976 23814 28988
rect 24578 28976 24584 28988
rect 24636 28976 24642 29028
rect 5810 28948 5816 28960
rect 5771 28920 5816 28948
rect 5810 28908 5816 28920
rect 5868 28908 5874 28960
rect 9766 28908 9772 28960
rect 9824 28948 9830 28960
rect 10134 28948 10140 28960
rect 9824 28920 10140 28948
rect 9824 28908 9830 28920
rect 10134 28908 10140 28920
rect 10192 28948 10198 28960
rect 10689 28951 10747 28957
rect 10689 28948 10701 28951
rect 10192 28920 10701 28948
rect 10192 28908 10198 28920
rect 10689 28917 10701 28920
rect 10735 28917 10747 28951
rect 10689 28911 10747 28917
rect 16482 28908 16488 28960
rect 16540 28948 16546 28960
rect 20806 28948 20812 28960
rect 16540 28920 20812 28948
rect 16540 28908 16546 28920
rect 20806 28908 20812 28920
rect 20864 28908 20870 28960
rect 20990 28908 20996 28960
rect 21048 28948 21054 28960
rect 22554 28948 22560 28960
rect 21048 28920 22560 28948
rect 21048 28908 21054 28920
rect 22554 28908 22560 28920
rect 22612 28948 22618 28960
rect 23290 28948 23296 28960
rect 22612 28920 23296 28948
rect 22612 28908 22618 28920
rect 23290 28908 23296 28920
rect 23348 28908 23354 28960
rect 23492 28948 23520 28976
rect 23842 28948 23848 28960
rect 23492 28920 23848 28948
rect 23842 28908 23848 28920
rect 23900 28908 23906 28960
rect 24964 28948 24992 29056
rect 25038 29044 25044 29096
rect 25096 29084 25102 29096
rect 25225 29087 25283 29093
rect 25096 29056 25189 29084
rect 25096 29044 25102 29056
rect 25225 29053 25237 29087
rect 25271 29053 25283 29087
rect 25866 29084 25872 29096
rect 25827 29056 25872 29084
rect 25225 29047 25283 29053
rect 25240 28948 25268 29047
rect 25866 29044 25872 29056
rect 25924 29044 25930 29096
rect 26053 29087 26111 29093
rect 26053 29053 26065 29087
rect 26099 29053 26111 29087
rect 26053 29047 26111 29053
rect 26068 29016 26096 29047
rect 26142 29044 26148 29096
rect 26200 29084 26206 29096
rect 26326 29093 26332 29096
rect 26283 29087 26332 29093
rect 26200 29056 26245 29084
rect 26200 29044 26206 29056
rect 26283 29053 26295 29087
rect 26329 29053 26332 29087
rect 26283 29047 26332 29053
rect 26326 29044 26332 29047
rect 26384 29044 26390 29096
rect 26418 29044 26424 29096
rect 26476 29084 26482 29096
rect 26476 29056 26521 29084
rect 26476 29044 26482 29056
rect 26694 29044 26700 29096
rect 26752 29084 26758 29096
rect 27982 29084 27988 29096
rect 26752 29056 27844 29084
rect 27943 29056 27988 29084
rect 26752 29044 26758 29056
rect 27706 29016 27712 29028
rect 26068 28988 27712 29016
rect 27706 28976 27712 28988
rect 27764 28976 27770 29028
rect 27816 29016 27844 29056
rect 27982 29044 27988 29056
rect 28040 29044 28046 29096
rect 28092 29093 28120 29124
rect 28184 29124 28273 29152
rect 28077 29087 28135 29093
rect 28077 29053 28089 29087
rect 28123 29053 28135 29087
rect 28077 29047 28135 29053
rect 28184 29016 28212 29124
rect 28261 29121 28273 29124
rect 28307 29121 28319 29155
rect 28261 29115 28319 29121
rect 31202 29112 31208 29164
rect 31260 29152 31266 29164
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31260 29124 32137 29152
rect 31260 29112 31266 29124
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 28353 29087 28411 29093
rect 28353 29053 28365 29087
rect 28399 29084 28411 29087
rect 28718 29084 28724 29096
rect 28399 29056 28724 29084
rect 28399 29053 28411 29056
rect 28353 29047 28411 29053
rect 28718 29044 28724 29056
rect 28776 29044 28782 29096
rect 28813 29087 28871 29093
rect 28813 29053 28825 29087
rect 28859 29084 28871 29087
rect 30374 29084 30380 29096
rect 28859 29056 30380 29084
rect 28859 29053 28871 29056
rect 28813 29047 28871 29053
rect 30374 29044 30380 29056
rect 30432 29044 30438 29096
rect 30929 29087 30987 29093
rect 30929 29084 30941 29087
rect 30852 29056 30941 29084
rect 27816 28988 28212 29016
rect 28994 28976 29000 29028
rect 29052 29025 29058 29028
rect 29052 29019 29116 29025
rect 29052 28985 29070 29019
rect 29104 28985 29116 29019
rect 30852 29016 30880 29056
rect 30929 29053 30941 29056
rect 30975 29053 30987 29087
rect 31570 29084 31576 29096
rect 31531 29056 31576 29084
rect 30929 29047 30987 29053
rect 31570 29044 31576 29056
rect 31628 29044 31634 29096
rect 33305 29093 33333 29180
rect 36633 29155 36691 29161
rect 36633 29121 36645 29155
rect 36679 29152 36691 29155
rect 50246 29152 50252 29164
rect 36679 29124 50252 29152
rect 36679 29121 36691 29124
rect 36633 29115 36691 29121
rect 50246 29112 50252 29124
rect 50304 29112 50310 29164
rect 54389 29155 54447 29161
rect 54389 29121 54401 29155
rect 54435 29152 54447 29155
rect 57517 29155 57575 29161
rect 57517 29152 57529 29155
rect 54435 29124 57529 29152
rect 54435 29121 54447 29124
rect 54389 29115 54447 29121
rect 57517 29121 57529 29124
rect 57563 29121 57575 29155
rect 57517 29115 57575 29121
rect 31757 29087 31815 29093
rect 31757 29053 31769 29087
rect 31803 29084 31815 29087
rect 33275 29087 33333 29093
rect 31803 29056 32352 29084
rect 31803 29053 31815 29056
rect 31757 29047 31815 29053
rect 31110 29016 31116 29028
rect 30852 28988 31116 29016
rect 29052 28979 29116 28985
rect 29052 28976 29058 28979
rect 31110 28976 31116 28988
rect 31168 29016 31174 29028
rect 31772 29016 31800 29047
rect 31168 28988 31800 29016
rect 31168 28976 31174 28988
rect 24964 28920 25268 28948
rect 27614 28908 27620 28960
rect 27672 28948 27678 28960
rect 28350 28948 28356 28960
rect 27672 28920 28356 28948
rect 27672 28908 27678 28920
rect 28350 28908 28356 28920
rect 28408 28908 28414 28960
rect 31021 28951 31079 28957
rect 31021 28917 31033 28951
rect 31067 28948 31079 28951
rect 31478 28948 31484 28960
rect 31067 28920 31484 28948
rect 31067 28917 31079 28920
rect 31021 28911 31079 28917
rect 31478 28908 31484 28920
rect 31536 28908 31542 28960
rect 32030 28948 32036 28960
rect 31991 28920 32036 28948
rect 32030 28908 32036 28920
rect 32088 28908 32094 28960
rect 32324 28948 32352 29056
rect 33275 29053 33287 29087
rect 33321 29053 33333 29087
rect 33410 29084 33416 29096
rect 33371 29056 33416 29084
rect 33275 29047 33333 29053
rect 33410 29044 33416 29056
rect 33468 29044 33474 29096
rect 33505 29087 33563 29093
rect 33505 29053 33517 29087
rect 33551 29053 33563 29087
rect 33686 29084 33692 29096
rect 33647 29056 33692 29084
rect 33505 29047 33563 29053
rect 33045 29019 33103 29025
rect 33045 28985 33057 29019
rect 33091 29016 33103 29019
rect 33134 29016 33140 29028
rect 33091 28988 33140 29016
rect 33091 28985 33103 28988
rect 33045 28979 33103 28985
rect 33134 28976 33140 28988
rect 33192 28976 33198 29028
rect 33428 28948 33456 29044
rect 33520 29006 33548 29047
rect 33686 29044 33692 29056
rect 33744 29044 33750 29096
rect 35434 29084 35440 29096
rect 35395 29056 35440 29084
rect 35434 29044 35440 29056
rect 35492 29044 35498 29096
rect 35618 29084 35624 29096
rect 35579 29056 35624 29084
rect 35618 29044 35624 29056
rect 35676 29044 35682 29096
rect 36265 29087 36323 29093
rect 36265 29053 36277 29087
rect 36311 29053 36323 29087
rect 36446 29084 36452 29096
rect 36407 29056 36452 29084
rect 36265 29047 36323 29053
rect 35452 29016 35480 29044
rect 36280 29016 36308 29047
rect 36446 29044 36452 29056
rect 36504 29044 36510 29096
rect 55033 29087 55091 29093
rect 55033 29053 55045 29087
rect 55079 29084 55091 29087
rect 55214 29084 55220 29096
rect 55079 29056 55220 29084
rect 55079 29053 55091 29056
rect 55033 29047 55091 29053
rect 55214 29044 55220 29056
rect 55272 29044 55278 29096
rect 55493 29087 55551 29093
rect 55493 29053 55505 29087
rect 55539 29084 55551 29087
rect 55674 29084 55680 29096
rect 55539 29056 55680 29084
rect 55539 29053 55551 29056
rect 55493 29047 55551 29053
rect 55674 29044 55680 29056
rect 55732 29084 55738 29096
rect 56226 29084 56232 29096
rect 55732 29056 56232 29084
rect 55732 29044 55738 29056
rect 56226 29044 56232 29056
rect 56284 29044 56290 29096
rect 56321 29087 56379 29093
rect 56321 29053 56333 29087
rect 56367 29084 56379 29087
rect 57422 29084 57428 29096
rect 56367 29056 57428 29084
rect 56367 29053 56379 29056
rect 56321 29047 56379 29053
rect 57422 29044 57428 29056
rect 57480 29044 57486 29096
rect 57698 29084 57704 29096
rect 57659 29056 57704 29084
rect 57698 29044 57704 29056
rect 57756 29044 57762 29096
rect 33502 28954 33508 29006
rect 33560 28954 33566 29006
rect 35452 28988 36308 29016
rect 56873 29019 56931 29025
rect 56873 28985 56885 29019
rect 56919 29016 56931 29019
rect 57330 29016 57336 29028
rect 56919 28988 57336 29016
rect 56919 28985 56931 28988
rect 56873 28979 56931 28985
rect 57330 28976 57336 28988
rect 57388 28976 57394 29028
rect 32324 28920 33456 28948
rect 1104 28858 58880 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 50326 28858
rect 50378 28806 50390 28858
rect 50442 28806 50454 28858
rect 50506 28806 50518 28858
rect 50570 28806 58880 28858
rect 1104 28784 58880 28806
rect 6454 28704 6460 28756
rect 6512 28744 6518 28756
rect 6549 28747 6607 28753
rect 6549 28744 6561 28747
rect 6512 28716 6561 28744
rect 6512 28704 6518 28716
rect 6549 28713 6561 28716
rect 6595 28713 6607 28747
rect 6549 28707 6607 28713
rect 7190 28704 7196 28756
rect 7248 28744 7254 28756
rect 7653 28747 7711 28753
rect 7653 28744 7665 28747
rect 7248 28716 7665 28744
rect 7248 28704 7254 28716
rect 7653 28713 7665 28716
rect 7699 28713 7711 28747
rect 9674 28744 9680 28756
rect 7653 28707 7711 28713
rect 9646 28704 9680 28744
rect 9732 28704 9738 28756
rect 12250 28744 12256 28756
rect 10796 28716 12256 28744
rect 5436 28679 5494 28685
rect 5436 28645 5448 28679
rect 5482 28676 5494 28679
rect 5810 28676 5816 28688
rect 5482 28648 5816 28676
rect 5482 28645 5494 28648
rect 5436 28639 5494 28645
rect 5810 28636 5816 28648
rect 5868 28636 5874 28688
rect 9646 28676 9674 28704
rect 10796 28676 10824 28716
rect 12250 28704 12256 28716
rect 12308 28704 12314 28756
rect 16592 28716 20944 28744
rect 7852 28648 9674 28676
rect 10520 28648 10824 28676
rect 10873 28679 10931 28685
rect 1489 28611 1547 28617
rect 1489 28577 1501 28611
rect 1535 28608 1547 28611
rect 2777 28611 2835 28617
rect 2777 28608 2789 28611
rect 1535 28580 2789 28608
rect 1535 28577 1547 28580
rect 1489 28571 1547 28577
rect 2777 28577 2789 28580
rect 2823 28577 2835 28611
rect 2777 28571 2835 28577
rect 4525 28611 4583 28617
rect 4525 28577 4537 28611
rect 4571 28577 4583 28611
rect 4706 28608 4712 28620
rect 4667 28580 4712 28608
rect 4525 28571 4583 28577
rect 1670 28540 1676 28552
rect 1631 28512 1676 28540
rect 1670 28500 1676 28512
rect 1728 28500 1734 28552
rect 4540 28540 4568 28571
rect 4706 28568 4712 28580
rect 4764 28568 4770 28620
rect 5169 28611 5227 28617
rect 5169 28577 5181 28611
rect 5215 28608 5227 28611
rect 6822 28608 6828 28620
rect 5215 28580 6828 28608
rect 5215 28577 5227 28580
rect 5169 28571 5227 28577
rect 6822 28568 6828 28580
rect 6880 28568 6886 28620
rect 7006 28608 7012 28620
rect 6967 28580 7012 28608
rect 7006 28568 7012 28580
rect 7064 28568 7070 28620
rect 7193 28611 7251 28617
rect 7193 28577 7205 28611
rect 7239 28608 7251 28611
rect 7282 28608 7288 28620
rect 7239 28580 7288 28608
rect 7239 28577 7251 28580
rect 7193 28571 7251 28577
rect 7282 28568 7288 28580
rect 7340 28568 7346 28620
rect 7852 28617 7880 28648
rect 7837 28611 7895 28617
rect 7837 28577 7849 28611
rect 7883 28577 7895 28611
rect 7837 28571 7895 28577
rect 7929 28611 7987 28617
rect 7929 28577 7941 28611
rect 7975 28577 7987 28611
rect 8202 28608 8208 28620
rect 8163 28580 8208 28608
rect 7929 28571 7987 28577
rect 4540 28512 5120 28540
rect 1854 28472 1860 28484
rect 1815 28444 1860 28472
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 4525 28475 4583 28481
rect 4525 28472 4537 28475
rect 2746 28444 4537 28472
rect 2590 28364 2596 28416
rect 2648 28404 2654 28416
rect 2746 28404 2774 28444
rect 4525 28441 4537 28444
rect 4571 28441 4583 28475
rect 4525 28435 4583 28441
rect 2648 28376 2774 28404
rect 5092 28404 5120 28512
rect 7558 28500 7564 28552
rect 7616 28540 7622 28552
rect 7944 28540 7972 28571
rect 8202 28568 8208 28580
rect 8260 28568 8266 28620
rect 9677 28611 9735 28617
rect 9677 28577 9689 28611
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 9769 28611 9827 28617
rect 9769 28577 9781 28611
rect 9815 28608 9827 28611
rect 9950 28608 9956 28620
rect 9815 28580 9956 28608
rect 9815 28577 9827 28580
rect 9769 28571 9827 28577
rect 7616 28512 7972 28540
rect 9692 28540 9720 28571
rect 9950 28568 9956 28580
rect 10008 28568 10014 28620
rect 10045 28611 10103 28617
rect 10045 28577 10057 28611
rect 10091 28608 10103 28611
rect 10134 28608 10140 28620
rect 10091 28580 10140 28608
rect 10091 28577 10103 28580
rect 10045 28571 10103 28577
rect 10134 28568 10140 28580
rect 10192 28568 10198 28620
rect 10520 28540 10548 28648
rect 10873 28645 10885 28679
rect 10919 28676 10931 28679
rect 11054 28676 11060 28688
rect 10919 28648 11060 28676
rect 10919 28645 10931 28648
rect 10873 28639 10931 28645
rect 11054 28636 11060 28648
rect 11112 28636 11118 28688
rect 12894 28676 12900 28688
rect 12544 28648 12900 28676
rect 11149 28611 11207 28617
rect 11149 28577 11161 28611
rect 11195 28608 11207 28611
rect 11330 28608 11336 28620
rect 11195 28580 11336 28608
rect 11195 28577 11207 28580
rect 11149 28571 11207 28577
rect 11330 28568 11336 28580
rect 11388 28568 11394 28620
rect 11514 28608 11520 28620
rect 11475 28580 11520 28608
rect 11514 28568 11520 28580
rect 11572 28568 11578 28620
rect 12544 28617 12572 28648
rect 12894 28636 12900 28648
rect 12952 28636 12958 28688
rect 13446 28636 13452 28688
rect 13504 28676 13510 28688
rect 13541 28679 13599 28685
rect 13541 28676 13553 28679
rect 13504 28648 13553 28676
rect 13504 28636 13510 28648
rect 13541 28645 13553 28648
rect 13587 28645 13599 28679
rect 13541 28639 13599 28645
rect 14918 28636 14924 28688
rect 14976 28685 14982 28688
rect 14976 28679 15040 28685
rect 14976 28645 14994 28679
rect 15028 28645 15040 28679
rect 14976 28639 15040 28645
rect 14976 28636 14982 28639
rect 12529 28611 12587 28617
rect 12529 28577 12541 28611
rect 12575 28577 12587 28611
rect 12710 28608 12716 28620
rect 12671 28580 12716 28608
rect 12529 28571 12587 28577
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 12989 28611 13047 28617
rect 12989 28577 13001 28611
rect 13035 28608 13047 28611
rect 16482 28608 16488 28620
rect 13035 28580 16488 28608
rect 13035 28577 13047 28580
rect 12989 28571 13047 28577
rect 16482 28568 16488 28580
rect 16540 28568 16546 28620
rect 16592 28617 16620 28716
rect 20248 28679 20306 28685
rect 16776 28648 20116 28676
rect 16776 28617 16804 28648
rect 16577 28611 16635 28617
rect 16577 28577 16589 28611
rect 16623 28577 16635 28611
rect 16577 28571 16635 28577
rect 16761 28611 16819 28617
rect 16761 28577 16773 28611
rect 16807 28577 16819 28611
rect 17218 28608 17224 28620
rect 17179 28580 17224 28608
rect 16761 28571 16819 28577
rect 17218 28568 17224 28580
rect 17276 28568 17282 28620
rect 17770 28608 17776 28620
rect 17731 28580 17776 28608
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 18598 28608 18604 28620
rect 18380 28580 18604 28608
rect 18380 28568 18386 28580
rect 18598 28568 18604 28580
rect 18656 28608 18662 28620
rect 18693 28611 18751 28617
rect 18693 28608 18705 28611
rect 18656 28580 18705 28608
rect 18656 28568 18662 28580
rect 18693 28577 18705 28580
rect 18739 28577 18751 28611
rect 18693 28571 18751 28577
rect 18785 28611 18843 28617
rect 18785 28577 18797 28611
rect 18831 28577 18843 28611
rect 18785 28571 18843 28577
rect 10686 28540 10692 28552
rect 9692 28512 10548 28540
rect 10647 28512 10692 28540
rect 7616 28500 7622 28512
rect 10686 28500 10692 28512
rect 10744 28500 10750 28552
rect 11241 28543 11299 28549
rect 11241 28509 11253 28543
rect 11287 28509 11299 28543
rect 11422 28540 11428 28552
rect 11383 28512 11428 28540
rect 11241 28503 11299 28509
rect 9766 28472 9772 28484
rect 6932 28444 9772 28472
rect 6932 28404 6960 28444
rect 9766 28432 9772 28444
rect 9824 28432 9830 28484
rect 11256 28472 11284 28503
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 12618 28540 12624 28552
rect 12579 28512 12624 28540
rect 12618 28500 12624 28512
rect 12676 28500 12682 28552
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28540 12863 28543
rect 12851 28512 13308 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 12345 28475 12403 28481
rect 12345 28472 12357 28475
rect 11256 28444 12357 28472
rect 12345 28441 12357 28444
rect 12391 28441 12403 28475
rect 12345 28435 12403 28441
rect 13280 28416 13308 28512
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 14737 28543 14795 28549
rect 14737 28540 14749 28543
rect 14424 28512 14749 28540
rect 14424 28500 14430 28512
rect 14737 28509 14749 28512
rect 14783 28509 14795 28543
rect 17862 28540 17868 28552
rect 17823 28512 17868 28540
rect 14737 28503 14795 28509
rect 17862 28500 17868 28512
rect 17920 28500 17926 28552
rect 17954 28500 17960 28552
rect 18012 28540 18018 28552
rect 18800 28540 18828 28571
rect 18874 28568 18880 28620
rect 18932 28608 18938 28620
rect 19058 28608 19064 28620
rect 18932 28580 18977 28608
rect 19019 28580 19064 28608
rect 18932 28568 18938 28580
rect 19058 28568 19064 28580
rect 19116 28568 19122 28620
rect 19150 28568 19156 28620
rect 19208 28608 19214 28620
rect 19981 28611 20039 28617
rect 19981 28608 19993 28611
rect 19208 28580 19993 28608
rect 19208 28568 19214 28580
rect 19981 28577 19993 28580
rect 20027 28577 20039 28611
rect 20088 28608 20116 28648
rect 20248 28645 20260 28679
rect 20294 28676 20306 28679
rect 20438 28676 20444 28688
rect 20294 28648 20444 28676
rect 20294 28645 20306 28648
rect 20248 28639 20306 28645
rect 20438 28636 20444 28648
rect 20496 28636 20502 28688
rect 20916 28676 20944 28716
rect 20990 28704 20996 28756
rect 21048 28744 21054 28756
rect 21361 28747 21419 28753
rect 21361 28744 21373 28747
rect 21048 28716 21373 28744
rect 21048 28704 21054 28716
rect 21361 28713 21373 28716
rect 21407 28713 21419 28747
rect 21818 28744 21824 28756
rect 21779 28716 21824 28744
rect 21361 28707 21419 28713
rect 21818 28704 21824 28716
rect 21876 28704 21882 28756
rect 22922 28744 22928 28756
rect 22883 28716 22928 28744
rect 22922 28704 22928 28716
rect 22980 28704 22986 28756
rect 24854 28704 24860 28756
rect 24912 28744 24918 28756
rect 26145 28747 26203 28753
rect 26145 28744 26157 28747
rect 24912 28716 26157 28744
rect 24912 28704 24918 28716
rect 26145 28713 26157 28716
rect 26191 28713 26203 28747
rect 26145 28707 26203 28713
rect 28077 28747 28135 28753
rect 28077 28713 28089 28747
rect 28123 28713 28135 28747
rect 28077 28707 28135 28713
rect 28537 28747 28595 28753
rect 28537 28713 28549 28747
rect 28583 28744 28595 28747
rect 28994 28744 29000 28756
rect 28583 28716 29000 28744
rect 28583 28713 28595 28716
rect 28537 28707 28595 28713
rect 22830 28676 22836 28688
rect 20916 28648 22836 28676
rect 22830 28636 22836 28648
rect 22888 28636 22894 28688
rect 23750 28676 23756 28688
rect 23124 28648 23756 28676
rect 21174 28608 21180 28620
rect 20088 28580 21180 28608
rect 19981 28571 20039 28577
rect 21174 28568 21180 28580
rect 21232 28568 21238 28620
rect 22002 28608 22008 28620
rect 21963 28580 22008 28608
rect 22002 28568 22008 28580
rect 22060 28568 22066 28620
rect 22097 28611 22155 28617
rect 22097 28577 22109 28611
rect 22143 28577 22155 28611
rect 22097 28571 22155 28577
rect 22373 28611 22431 28617
rect 22373 28577 22385 28611
rect 22419 28608 22431 28611
rect 22554 28608 22560 28620
rect 22419 28580 22560 28608
rect 22419 28577 22431 28580
rect 22373 28571 22431 28577
rect 19334 28540 19340 28552
rect 18012 28512 19340 28540
rect 18012 28500 18018 28512
rect 19334 28500 19340 28512
rect 19392 28500 19398 28552
rect 22112 28540 22140 28571
rect 22554 28568 22560 28580
rect 22612 28568 22618 28620
rect 23124 28617 23152 28648
rect 23750 28636 23756 28648
rect 23808 28636 23814 28688
rect 24026 28636 24032 28688
rect 24084 28676 24090 28688
rect 27341 28679 27399 28685
rect 24084 28648 26740 28676
rect 24084 28636 24090 28648
rect 23109 28611 23167 28617
rect 23109 28577 23121 28611
rect 23155 28577 23167 28611
rect 23109 28571 23167 28577
rect 23201 28611 23259 28617
rect 23201 28577 23213 28611
rect 23247 28577 23259 28611
rect 23474 28608 23480 28620
rect 23435 28580 23480 28608
rect 23201 28571 23259 28577
rect 22278 28540 22284 28552
rect 22066 28512 22140 28540
rect 22239 28512 22284 28540
rect 15746 28432 15752 28484
rect 15804 28472 15810 28484
rect 22066 28472 22094 28512
rect 22278 28500 22284 28512
rect 22336 28500 22342 28552
rect 23216 28540 23244 28571
rect 23474 28568 23480 28580
rect 23532 28568 23538 28620
rect 23934 28608 23940 28620
rect 23895 28580 23940 28608
rect 23934 28568 23940 28580
rect 23992 28568 23998 28620
rect 25501 28611 25559 28617
rect 25501 28577 25513 28611
rect 25547 28608 25559 28611
rect 25682 28608 25688 28620
rect 25547 28580 25688 28608
rect 25547 28577 25559 28580
rect 25501 28571 25559 28577
rect 25682 28568 25688 28580
rect 25740 28568 25746 28620
rect 26712 28617 26740 28648
rect 27341 28645 27353 28679
rect 27387 28676 27399 28679
rect 27798 28676 27804 28688
rect 27387 28648 27421 28676
rect 27759 28648 27804 28676
rect 27387 28645 27399 28648
rect 27341 28639 27399 28645
rect 26697 28611 26755 28617
rect 25792 28580 26648 28608
rect 24029 28543 24087 28549
rect 24029 28540 24041 28543
rect 23216 28512 24041 28540
rect 24029 28509 24041 28512
rect 24075 28509 24087 28543
rect 25792 28540 25820 28580
rect 24029 28503 24087 28509
rect 25700 28512 25820 28540
rect 25869 28543 25927 28549
rect 22738 28472 22744 28484
rect 15804 28444 19334 28472
rect 15804 28432 15810 28444
rect 5092 28376 6960 28404
rect 7009 28407 7067 28413
rect 2648 28364 2654 28376
rect 7009 28373 7021 28407
rect 7055 28404 7067 28407
rect 7098 28404 7104 28416
rect 7055 28376 7104 28404
rect 7055 28373 7067 28376
rect 7009 28367 7067 28373
rect 7098 28364 7104 28376
rect 7156 28364 7162 28416
rect 8110 28404 8116 28416
rect 8071 28376 8116 28404
rect 8110 28364 8116 28376
rect 8168 28364 8174 28416
rect 9398 28364 9404 28416
rect 9456 28404 9462 28416
rect 9493 28407 9551 28413
rect 9493 28404 9505 28407
rect 9456 28376 9505 28404
rect 9456 28364 9462 28376
rect 9493 28373 9505 28376
rect 9539 28373 9551 28407
rect 9950 28404 9956 28416
rect 9911 28376 9956 28404
rect 9493 28367 9551 28373
rect 9950 28364 9956 28376
rect 10008 28364 10014 28416
rect 13262 28364 13268 28416
rect 13320 28404 13326 28416
rect 13633 28407 13691 28413
rect 13633 28404 13645 28407
rect 13320 28376 13645 28404
rect 13320 28364 13326 28376
rect 13633 28373 13645 28376
rect 13679 28373 13691 28407
rect 13633 28367 13691 28373
rect 15102 28364 15108 28416
rect 15160 28404 15166 28416
rect 16117 28407 16175 28413
rect 16117 28404 16129 28407
rect 15160 28376 16129 28404
rect 15160 28364 15166 28376
rect 16117 28373 16129 28376
rect 16163 28373 16175 28407
rect 16117 28367 16175 28373
rect 16574 28364 16580 28416
rect 16632 28404 16638 28416
rect 16669 28407 16727 28413
rect 16669 28404 16681 28407
rect 16632 28376 16681 28404
rect 16632 28364 16638 28376
rect 16669 28373 16681 28376
rect 16715 28373 16727 28407
rect 16669 28367 16727 28373
rect 18230 28364 18236 28416
rect 18288 28404 18294 28416
rect 18417 28407 18475 28413
rect 18417 28404 18429 28407
rect 18288 28376 18429 28404
rect 18288 28364 18294 28376
rect 18417 28373 18429 28376
rect 18463 28373 18475 28407
rect 19306 28404 19334 28444
rect 22066 28444 22744 28472
rect 22066 28404 22094 28444
rect 22738 28432 22744 28444
rect 22796 28432 22802 28484
rect 23934 28432 23940 28484
rect 23992 28472 23998 28484
rect 25700 28472 25728 28512
rect 25869 28509 25881 28543
rect 25915 28540 25927 28543
rect 26050 28540 26056 28552
rect 25915 28512 26056 28540
rect 25915 28509 25927 28512
rect 25869 28503 25927 28509
rect 26050 28500 26056 28512
rect 26108 28500 26114 28552
rect 26620 28540 26648 28580
rect 26697 28577 26709 28611
rect 26743 28577 26755 28611
rect 26878 28608 26884 28620
rect 26839 28580 26884 28608
rect 26697 28571 26755 28577
rect 26878 28568 26884 28580
rect 26936 28568 26942 28620
rect 27356 28608 27384 28639
rect 27798 28636 27804 28648
rect 27856 28636 27862 28688
rect 28092 28676 28120 28707
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 30374 28704 30380 28756
rect 30432 28744 30438 28756
rect 32309 28747 32367 28753
rect 30432 28716 31754 28744
rect 30432 28704 30438 28716
rect 31018 28676 31024 28688
rect 28092 28648 29224 28676
rect 27614 28617 27620 28620
rect 27433 28611 27491 28617
rect 27433 28608 27445 28611
rect 27264 28580 27445 28608
rect 27264 28540 27292 28580
rect 27433 28577 27445 28580
rect 27479 28577 27491 28611
rect 27433 28571 27491 28577
rect 27571 28611 27620 28617
rect 27571 28577 27583 28611
rect 27617 28577 27620 28611
rect 27571 28571 27620 28577
rect 27614 28568 27620 28571
rect 27672 28568 27678 28620
rect 27709 28611 27767 28617
rect 27709 28577 27721 28611
rect 27755 28577 27767 28611
rect 27709 28571 27767 28577
rect 26620 28512 27292 28540
rect 27338 28500 27344 28552
rect 27396 28540 27402 28552
rect 27724 28540 27752 28571
rect 27890 28568 27896 28620
rect 27948 28617 27954 28620
rect 27948 28608 27956 28617
rect 28767 28611 28825 28617
rect 28767 28608 28779 28611
rect 27948 28580 27993 28608
rect 28460 28580 28779 28608
rect 27948 28571 27956 28580
rect 27948 28568 27954 28571
rect 27396 28512 27752 28540
rect 27396 28500 27402 28512
rect 23992 28444 25728 28472
rect 25777 28475 25835 28481
rect 23992 28432 23998 28444
rect 25777 28441 25789 28475
rect 25823 28472 25835 28475
rect 27356 28472 27384 28500
rect 25823 28444 27384 28472
rect 25823 28441 25835 28444
rect 25777 28435 25835 28441
rect 27798 28432 27804 28484
rect 27856 28472 27862 28484
rect 28460 28472 28488 28580
rect 28767 28577 28779 28580
rect 28813 28577 28825 28611
rect 28767 28571 28825 28577
rect 28905 28611 28963 28617
rect 28905 28577 28917 28611
rect 28951 28577 28963 28611
rect 28905 28571 28963 28577
rect 28534 28500 28540 28552
rect 28592 28540 28598 28552
rect 28920 28540 28948 28571
rect 28994 28568 29000 28620
rect 29052 28608 29058 28620
rect 29196 28617 29224 28648
rect 30944 28648 31024 28676
rect 30944 28617 30972 28648
rect 31018 28636 31024 28648
rect 31076 28636 31082 28688
rect 31202 28676 31208 28688
rect 31163 28648 31208 28676
rect 31202 28636 31208 28648
rect 31260 28636 31266 28688
rect 31726 28676 31754 28716
rect 32309 28713 32321 28747
rect 32355 28744 32367 28747
rect 33686 28744 33692 28756
rect 32355 28716 33692 28744
rect 32355 28713 32367 28716
rect 32309 28707 32367 28713
rect 33686 28704 33692 28716
rect 33744 28704 33750 28756
rect 34425 28747 34483 28753
rect 34425 28713 34437 28747
rect 34471 28713 34483 28747
rect 58066 28744 58072 28756
rect 34425 28707 34483 28713
rect 55784 28716 58072 28744
rect 32858 28676 32864 28688
rect 31726 28648 32864 28676
rect 32858 28636 32864 28648
rect 32916 28636 32922 28688
rect 33226 28636 33232 28688
rect 33284 28685 33290 28688
rect 33284 28679 33348 28685
rect 33284 28645 33302 28679
rect 33336 28645 33348 28679
rect 33284 28639 33348 28645
rect 33284 28636 33290 28639
rect 33410 28636 33416 28688
rect 33468 28676 33474 28688
rect 34440 28676 34468 28707
rect 33468 28648 34468 28676
rect 55217 28679 55275 28685
rect 33468 28636 33474 28648
rect 55217 28645 55229 28679
rect 55263 28676 55275 28679
rect 55306 28676 55312 28688
rect 55263 28648 55312 28676
rect 55263 28645 55275 28648
rect 55217 28639 55275 28645
rect 55306 28636 55312 28648
rect 55364 28636 55370 28688
rect 55784 28685 55812 28716
rect 58066 28704 58072 28716
rect 58124 28704 58130 28756
rect 55769 28679 55827 28685
rect 55769 28645 55781 28679
rect 55815 28645 55827 28679
rect 55769 28639 55827 28645
rect 56226 28636 56232 28688
rect 56284 28676 56290 28688
rect 56873 28679 56931 28685
rect 56873 28676 56885 28679
rect 56284 28648 56885 28676
rect 56284 28636 56290 28648
rect 56873 28645 56885 28648
rect 56919 28645 56931 28679
rect 58158 28676 58164 28688
rect 58119 28648 58164 28676
rect 56873 28639 56931 28645
rect 58158 28636 58164 28648
rect 58216 28636 58222 28688
rect 29181 28611 29239 28617
rect 29052 28580 29097 28608
rect 29052 28568 29058 28580
rect 29181 28577 29193 28611
rect 29227 28577 29239 28611
rect 29181 28571 29239 28577
rect 30929 28611 30987 28617
rect 30929 28577 30941 28611
rect 30975 28577 30987 28611
rect 31110 28608 31116 28620
rect 31071 28580 31116 28608
rect 30929 28571 30987 28577
rect 31110 28568 31116 28580
rect 31168 28568 31174 28620
rect 31654 28611 31712 28617
rect 31654 28608 31666 28611
rect 31588 28580 31666 28608
rect 28592 28512 28948 28540
rect 31588 28540 31616 28580
rect 31654 28577 31666 28580
rect 31700 28577 31712 28611
rect 31654 28571 31712 28577
rect 31754 28568 31760 28620
rect 31812 28608 31818 28620
rect 31938 28608 31944 28620
rect 31812 28580 31857 28608
rect 31899 28580 31944 28608
rect 31812 28568 31818 28580
rect 31938 28568 31944 28580
rect 31996 28568 32002 28620
rect 32030 28568 32036 28620
rect 32088 28608 32094 28620
rect 32171 28611 32229 28617
rect 32088 28580 32133 28608
rect 32088 28568 32094 28580
rect 32171 28577 32183 28611
rect 32217 28608 32229 28611
rect 33778 28608 33784 28620
rect 32217 28580 33784 28608
rect 32217 28577 32229 28580
rect 32171 28571 32229 28577
rect 33778 28568 33784 28580
rect 33836 28568 33842 28620
rect 35710 28608 35716 28620
rect 35671 28580 35716 28608
rect 35710 28568 35716 28580
rect 35768 28568 35774 28620
rect 54389 28611 54447 28617
rect 54389 28577 54401 28611
rect 54435 28577 54447 28611
rect 54389 28571 54447 28577
rect 57977 28611 58035 28617
rect 57977 28577 57989 28611
rect 58023 28608 58035 28611
rect 58066 28608 58072 28620
rect 58023 28580 58072 28608
rect 58023 28577 58035 28580
rect 57977 28571 58035 28577
rect 32582 28540 32588 28552
rect 31588 28512 32588 28540
rect 28592 28500 28598 28512
rect 31294 28472 31300 28484
rect 27856 28444 31300 28472
rect 27856 28432 27862 28444
rect 31294 28432 31300 28444
rect 31352 28432 31358 28484
rect 19306 28376 22094 28404
rect 18417 28367 18475 28373
rect 23198 28364 23204 28416
rect 23256 28404 23262 28416
rect 23385 28407 23443 28413
rect 23385 28404 23397 28407
rect 23256 28376 23397 28404
rect 23256 28364 23262 28376
rect 23385 28373 23397 28376
rect 23431 28373 23443 28407
rect 23385 28367 23443 28373
rect 25590 28364 25596 28416
rect 25648 28413 25654 28416
rect 25648 28407 25697 28413
rect 25648 28373 25651 28407
rect 25685 28373 25697 28407
rect 25648 28367 25697 28373
rect 25648 28364 25654 28367
rect 25866 28364 25872 28416
rect 25924 28404 25930 28416
rect 26697 28407 26755 28413
rect 26697 28404 26709 28407
rect 25924 28376 26709 28404
rect 25924 28364 25930 28376
rect 26697 28373 26709 28376
rect 26743 28373 26755 28407
rect 26697 28367 26755 28373
rect 27341 28407 27399 28413
rect 27341 28373 27353 28407
rect 27387 28404 27399 28407
rect 31588 28404 31616 28512
rect 32582 28500 32588 28512
rect 32640 28500 32646 28552
rect 32858 28500 32864 28552
rect 32916 28540 32922 28552
rect 33045 28543 33103 28549
rect 33045 28540 33057 28543
rect 32916 28512 33057 28540
rect 32916 28500 32922 28512
rect 33045 28509 33057 28512
rect 33091 28509 33103 28543
rect 33045 28503 33103 28509
rect 54404 28472 54432 28571
rect 58066 28568 58072 28580
rect 58124 28568 58130 28620
rect 55122 28540 55128 28552
rect 55083 28512 55128 28540
rect 55122 28500 55128 28512
rect 55180 28500 55186 28552
rect 56778 28540 56784 28552
rect 56739 28512 56784 28540
rect 56778 28500 56784 28512
rect 56836 28500 56842 28552
rect 57425 28543 57483 28549
rect 57425 28509 57437 28543
rect 57471 28540 57483 28543
rect 58710 28540 58716 28552
rect 57471 28512 58716 28540
rect 57471 28509 57483 28512
rect 57425 28503 57483 28509
rect 58710 28500 58716 28512
rect 58768 28500 58774 28552
rect 55582 28472 55588 28484
rect 54404 28444 55588 28472
rect 55582 28432 55588 28444
rect 55640 28432 55646 28484
rect 27387 28376 31616 28404
rect 27387 28373 27399 28376
rect 27341 28367 27399 28373
rect 35434 28364 35440 28416
rect 35492 28404 35498 28416
rect 35897 28407 35955 28413
rect 35897 28404 35909 28407
rect 35492 28376 35909 28404
rect 35492 28364 35498 28376
rect 35897 28373 35909 28376
rect 35943 28373 35955 28407
rect 35897 28367 35955 28373
rect 1104 28314 58880 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 58880 28314
rect 1104 28240 58880 28262
rect 2958 28200 2964 28212
rect 2919 28172 2964 28200
rect 2958 28160 2964 28172
rect 3016 28160 3022 28212
rect 6914 28160 6920 28212
rect 6972 28200 6978 28212
rect 7101 28203 7159 28209
rect 7101 28200 7113 28203
rect 6972 28172 7113 28200
rect 6972 28160 6978 28172
rect 7101 28169 7113 28172
rect 7147 28169 7159 28203
rect 15746 28200 15752 28212
rect 7101 28163 7159 28169
rect 7300 28172 15752 28200
rect 2590 28064 2596 28076
rect 2551 28036 2596 28064
rect 2590 28024 2596 28036
rect 2648 28024 2654 28076
rect 4448 28036 6224 28064
rect 2774 27956 2780 28008
rect 2832 27996 2838 28008
rect 4448 28005 4476 28036
rect 4433 27999 4491 28005
rect 2832 27968 2877 27996
rect 2832 27956 2838 27968
rect 4433 27965 4445 27999
rect 4479 27965 4491 27999
rect 4433 27959 4491 27965
rect 4617 27999 4675 28005
rect 4617 27965 4629 27999
rect 4663 27996 4675 27999
rect 4706 27996 4712 28008
rect 4663 27968 4712 27996
rect 4663 27965 4675 27968
rect 4617 27959 4675 27965
rect 4706 27956 4712 27968
rect 4764 27956 4770 28008
rect 5074 27996 5080 28008
rect 5035 27968 5080 27996
rect 5074 27956 5080 27968
rect 5132 27956 5138 28008
rect 5261 27999 5319 28005
rect 5261 27965 5273 27999
rect 5307 27965 5319 27999
rect 5261 27959 5319 27965
rect 1854 27928 1860 27940
rect 1815 27900 1860 27928
rect 1854 27888 1860 27900
rect 1912 27888 1918 27940
rect 4724 27928 4752 27956
rect 5270 27928 5298 27959
rect 4724 27900 5298 27928
rect 6196 27928 6224 28036
rect 7300 28005 7328 28172
rect 15746 28160 15752 28172
rect 15804 28160 15810 28212
rect 17678 28160 17684 28212
rect 17736 28200 17742 28212
rect 17736 28172 18920 28200
rect 17736 28160 17742 28172
rect 11149 28135 11207 28141
rect 11149 28101 11161 28135
rect 11195 28132 11207 28135
rect 11238 28132 11244 28144
rect 11195 28104 11244 28132
rect 11195 28101 11207 28104
rect 11149 28095 11207 28101
rect 11238 28092 11244 28104
rect 11296 28132 11302 28144
rect 11422 28132 11428 28144
rect 11296 28104 11428 28132
rect 11296 28092 11302 28104
rect 11422 28092 11428 28104
rect 11480 28092 11486 28144
rect 15654 28132 15660 28144
rect 15028 28104 15660 28132
rect 7561 28067 7619 28073
rect 7561 28033 7573 28067
rect 7607 28064 7619 28067
rect 8110 28064 8116 28076
rect 7607 28036 8116 28064
rect 7607 28033 7619 28036
rect 7561 28027 7619 28033
rect 8110 28024 8116 28036
rect 8168 28024 8174 28076
rect 9582 28024 9588 28076
rect 9640 28064 9646 28076
rect 12986 28064 12992 28076
rect 9640 28036 12756 28064
rect 12947 28036 12992 28064
rect 9640 28024 9646 28036
rect 7285 27999 7343 28005
rect 7285 27965 7297 27999
rect 7331 27965 7343 27999
rect 7285 27959 7343 27965
rect 7377 27999 7435 28005
rect 7377 27965 7389 27999
rect 7423 27996 7435 27999
rect 7466 27996 7472 28008
rect 7423 27968 7472 27996
rect 7423 27965 7435 27968
rect 7377 27959 7435 27965
rect 7466 27956 7472 27968
rect 7524 27956 7530 28008
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27965 7711 27999
rect 7653 27959 7711 27965
rect 8573 27999 8631 28005
rect 8573 27965 8585 27999
rect 8619 27996 8631 27999
rect 8662 27996 8668 28008
rect 8619 27968 8668 27996
rect 8619 27965 8631 27968
rect 8573 27959 8631 27965
rect 6546 27928 6552 27940
rect 6196 27900 6552 27928
rect 6546 27888 6552 27900
rect 6604 27928 6610 27940
rect 7668 27928 7696 27959
rect 8662 27956 8668 27968
rect 8720 27956 8726 28008
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11146 27996 11152 28008
rect 11011 27968 11152 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11146 27956 11152 27968
rect 11204 27996 11210 28008
rect 11790 27996 11796 28008
rect 11204 27968 11796 27996
rect 11204 27956 11210 27968
rect 11790 27956 11796 27968
rect 11848 27956 11854 28008
rect 12066 27996 12072 28008
rect 12027 27968 12072 27996
rect 12066 27956 12072 27968
rect 12124 27956 12130 28008
rect 12728 28005 12756 28036
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 15028 28064 15056 28104
rect 15654 28092 15660 28104
rect 15712 28092 15718 28144
rect 15930 28092 15936 28144
rect 15988 28132 15994 28144
rect 17954 28132 17960 28144
rect 15988 28104 17960 28132
rect 15988 28092 15994 28104
rect 17954 28092 17960 28104
rect 18012 28092 18018 28144
rect 18892 28132 18920 28172
rect 19058 28160 19064 28212
rect 19116 28200 19122 28212
rect 19981 28203 20039 28209
rect 19981 28200 19993 28203
rect 19116 28172 19993 28200
rect 19116 28160 19122 28172
rect 19981 28169 19993 28172
rect 20027 28169 20039 28203
rect 19981 28163 20039 28169
rect 21082 28160 21088 28212
rect 21140 28200 21146 28212
rect 21269 28203 21327 28209
rect 21269 28200 21281 28203
rect 21140 28172 21281 28200
rect 21140 28160 21146 28172
rect 21269 28169 21281 28172
rect 21315 28169 21327 28203
rect 21269 28163 21327 28169
rect 23106 28160 23112 28212
rect 23164 28200 23170 28212
rect 23385 28203 23443 28209
rect 23385 28200 23397 28203
rect 23164 28172 23397 28200
rect 23164 28160 23170 28172
rect 23385 28169 23397 28172
rect 23431 28169 23443 28203
rect 25866 28200 25872 28212
rect 23385 28163 23443 28169
rect 24044 28172 25872 28200
rect 18892 28104 19288 28132
rect 15749 28067 15807 28073
rect 15749 28064 15761 28067
rect 13188 28036 15056 28064
rect 15120 28036 15761 28064
rect 13188 28008 13216 28036
rect 15120 28008 15148 28036
rect 15749 28033 15761 28036
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 15838 28024 15844 28076
rect 15896 28064 15902 28076
rect 17405 28067 17463 28073
rect 15896 28036 16436 28064
rect 15896 28024 15902 28036
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27996 12771 27999
rect 13170 27996 13176 28008
rect 12759 27968 13176 27996
rect 12759 27965 12771 27968
rect 12713 27959 12771 27965
rect 13170 27956 13176 27968
rect 13228 27956 13234 28008
rect 13722 27996 13728 28008
rect 13683 27968 13728 27996
rect 13722 27956 13728 27968
rect 13780 27956 13786 28008
rect 14458 27996 14464 28008
rect 14419 27968 14464 27996
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 15102 27996 15108 28008
rect 15063 27968 15108 27996
rect 15102 27956 15108 27968
rect 15160 27956 15166 28008
rect 15194 27956 15200 28008
rect 15252 27996 15258 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 15252 27968 15301 27996
rect 15252 27956 15258 27968
rect 15289 27965 15301 27968
rect 15335 27996 15347 27999
rect 15930 27996 15936 28008
rect 15335 27968 15936 27996
rect 15335 27965 15347 27968
rect 15289 27959 15347 27965
rect 15930 27956 15936 27968
rect 15988 27956 15994 28008
rect 16301 27999 16359 28005
rect 16301 27965 16313 27999
rect 16347 27965 16359 27999
rect 16301 27959 16359 27965
rect 6604 27900 7696 27928
rect 6604 27888 6610 27900
rect 8478 27888 8484 27940
rect 8536 27928 8542 27940
rect 8818 27931 8876 27937
rect 8818 27928 8830 27931
rect 8536 27900 8830 27928
rect 8536 27888 8542 27900
rect 8818 27897 8830 27900
rect 8864 27897 8876 27931
rect 8818 27891 8876 27897
rect 10042 27888 10048 27940
rect 10100 27928 10106 27940
rect 13906 27928 13912 27940
rect 10100 27900 13912 27928
rect 10100 27888 10106 27900
rect 13906 27888 13912 27900
rect 13964 27888 13970 27940
rect 14553 27931 14611 27937
rect 14553 27897 14565 27931
rect 14599 27928 14611 27931
rect 15470 27928 15476 27940
rect 14599 27900 15476 27928
rect 14599 27897 14611 27900
rect 14553 27891 14611 27897
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 16316 27928 16344 27959
rect 15580 27900 16344 27928
rect 15580 27872 15608 27900
rect 1946 27860 1952 27872
rect 1907 27832 1952 27860
rect 1946 27820 1952 27832
rect 2004 27820 2010 27872
rect 4525 27863 4583 27869
rect 4525 27829 4537 27863
rect 4571 27860 4583 27863
rect 4890 27860 4896 27872
rect 4571 27832 4896 27860
rect 4571 27829 4583 27832
rect 4525 27823 4583 27829
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 5074 27820 5080 27872
rect 5132 27860 5138 27872
rect 5169 27863 5227 27869
rect 5169 27860 5181 27863
rect 5132 27832 5181 27860
rect 5132 27820 5138 27832
rect 5169 27829 5181 27832
rect 5215 27829 5227 27863
rect 5169 27823 5227 27829
rect 9953 27863 10011 27869
rect 9953 27829 9965 27863
rect 9999 27860 10011 27863
rect 10594 27860 10600 27872
rect 9999 27832 10600 27860
rect 9999 27829 10011 27832
rect 9953 27823 10011 27829
rect 10594 27820 10600 27832
rect 10652 27820 10658 27872
rect 12161 27863 12219 27869
rect 12161 27829 12173 27863
rect 12207 27860 12219 27863
rect 13998 27860 14004 27872
rect 12207 27832 14004 27860
rect 12207 27829 12219 27832
rect 12161 27823 12219 27829
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 15197 27863 15255 27869
rect 15197 27829 15209 27863
rect 15243 27860 15255 27863
rect 15562 27860 15568 27872
rect 15243 27832 15568 27860
rect 15243 27829 15255 27832
rect 15197 27823 15255 27829
rect 15562 27820 15568 27832
rect 15620 27820 15626 27872
rect 16206 27860 16212 27872
rect 16167 27832 16212 27860
rect 16206 27820 16212 27832
rect 16264 27820 16270 27872
rect 16408 27860 16436 28036
rect 17405 28033 17417 28067
rect 17451 28064 17463 28067
rect 19260 28064 19288 28104
rect 19334 28092 19340 28144
rect 19392 28132 19398 28144
rect 19392 28104 19437 28132
rect 19392 28092 19398 28104
rect 20530 28092 20536 28144
rect 20588 28132 20594 28144
rect 23937 28135 23995 28141
rect 23937 28132 23949 28135
rect 20588 28104 23949 28132
rect 20588 28092 20594 28104
rect 23937 28101 23949 28104
rect 23983 28101 23995 28135
rect 23937 28095 23995 28101
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 17451 28036 18092 28064
rect 19260 28036 19901 28064
rect 17451 28033 17463 28036
rect 17405 28027 17463 28033
rect 18064 28008 18092 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 20073 28067 20131 28073
rect 20073 28033 20085 28067
rect 20119 28033 20131 28067
rect 20073 28027 20131 28033
rect 20180 28036 20944 28064
rect 17310 27996 17316 28008
rect 17271 27968 17316 27996
rect 17310 27956 17316 27968
rect 17368 27996 17374 28008
rect 17586 27996 17592 28008
rect 17368 27968 17592 27996
rect 17368 27956 17374 27968
rect 17586 27956 17592 27968
rect 17644 27956 17650 28008
rect 17954 27996 17960 28008
rect 17915 27968 17960 27996
rect 17954 27956 17960 27968
rect 18012 27956 18018 28008
rect 18046 27956 18052 28008
rect 18104 27956 18110 28008
rect 18230 28005 18236 28008
rect 18224 27996 18236 28005
rect 18191 27968 18236 27996
rect 18224 27959 18236 27968
rect 18230 27956 18236 27959
rect 18288 27956 18294 28008
rect 18598 27956 18604 28008
rect 18656 27996 18662 28008
rect 19797 27999 19855 28005
rect 19797 27996 19809 27999
rect 18656 27968 19809 27996
rect 18656 27956 18662 27968
rect 19797 27965 19809 27968
rect 19843 27965 19855 27999
rect 19797 27959 19855 27965
rect 16482 27888 16488 27940
rect 16540 27928 16546 27940
rect 20088 27928 20116 28027
rect 16540 27900 20116 27928
rect 16540 27888 16546 27900
rect 20180 27860 20208 28036
rect 20622 27996 20628 28008
rect 20583 27968 20628 27996
rect 20622 27956 20628 27968
rect 20680 27956 20686 28008
rect 20714 27956 20720 28008
rect 20772 27996 20778 28008
rect 20916 27996 20944 28036
rect 23382 28024 23388 28076
rect 23440 28064 23446 28076
rect 24044 28064 24072 28172
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 25961 28203 26019 28209
rect 25961 28169 25973 28203
rect 26007 28200 26019 28203
rect 26142 28200 26148 28212
rect 26007 28172 26148 28200
rect 26007 28169 26019 28172
rect 25961 28163 26019 28169
rect 26142 28160 26148 28172
rect 26200 28160 26206 28212
rect 27522 28160 27528 28212
rect 27580 28200 27586 28212
rect 28353 28203 28411 28209
rect 28353 28200 28365 28203
rect 27580 28172 28365 28200
rect 27580 28160 27586 28172
rect 28353 28169 28365 28172
rect 28399 28169 28411 28203
rect 55306 28200 55312 28212
rect 28353 28163 28411 28169
rect 31128 28172 34560 28200
rect 55267 28172 55312 28200
rect 24765 28135 24823 28141
rect 24765 28101 24777 28135
rect 24811 28132 24823 28135
rect 26234 28132 26240 28144
rect 24811 28104 26240 28132
rect 24811 28101 24823 28104
rect 24765 28095 24823 28101
rect 26234 28092 26240 28104
rect 26292 28092 26298 28144
rect 26326 28092 26332 28144
rect 26384 28132 26390 28144
rect 26602 28132 26608 28144
rect 26384 28104 26608 28132
rect 26384 28092 26390 28104
rect 26602 28092 26608 28104
rect 26660 28132 26666 28144
rect 28074 28132 28080 28144
rect 26660 28104 28080 28132
rect 26660 28092 26666 28104
rect 28074 28092 28080 28104
rect 28132 28092 28138 28144
rect 23440 28036 24072 28064
rect 24489 28067 24547 28073
rect 23440 28024 23446 28036
rect 24489 28033 24501 28067
rect 24535 28064 24547 28067
rect 24535 28036 25084 28064
rect 24535 28033 24547 28036
rect 24489 28027 24547 28033
rect 21090 27999 21148 28005
rect 21090 27996 21102 27999
rect 20772 27968 20817 27996
rect 20916 27968 21102 27996
rect 20772 27956 20778 27968
rect 21090 27965 21102 27968
rect 21136 27965 21148 27999
rect 21090 27959 21148 27965
rect 22278 27956 22284 28008
rect 22336 27996 22342 28008
rect 22833 27999 22891 28005
rect 22833 27996 22845 27999
rect 22336 27968 22845 27996
rect 22336 27956 22342 27968
rect 22833 27965 22845 27968
rect 22879 27965 22891 27999
rect 23198 27996 23204 28008
rect 23159 27968 23204 27996
rect 22833 27959 22891 27965
rect 23198 27956 23204 27968
rect 23256 27956 23262 28008
rect 23842 27996 23848 28008
rect 23803 27968 23848 27996
rect 23842 27956 23848 27968
rect 23900 27956 23906 28008
rect 25056 28005 25084 28036
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 25280 28036 26004 28064
rect 25280 28024 25286 28036
rect 24673 27999 24731 28005
rect 24673 27965 24685 27999
rect 24719 27996 24731 27999
rect 25041 27999 25099 28005
rect 24719 27968 24992 27996
rect 24719 27965 24731 27968
rect 24673 27959 24731 27965
rect 20901 27931 20959 27937
rect 20901 27897 20913 27931
rect 20947 27897 20959 27931
rect 20901 27891 20959 27897
rect 20993 27931 21051 27937
rect 20993 27897 21005 27931
rect 21039 27928 21051 27931
rect 21358 27928 21364 27940
rect 21039 27900 21364 27928
rect 21039 27897 21051 27900
rect 20993 27891 21051 27897
rect 16408 27832 20208 27860
rect 20916 27860 20944 27891
rect 21358 27888 21364 27900
rect 21416 27928 21422 27940
rect 21818 27928 21824 27940
rect 21416 27900 21824 27928
rect 21416 27888 21422 27900
rect 21818 27888 21824 27900
rect 21876 27888 21882 27940
rect 22554 27888 22560 27940
rect 22612 27928 22618 27940
rect 23017 27931 23075 27937
rect 23017 27928 23029 27931
rect 22612 27900 23029 27928
rect 22612 27888 22618 27900
rect 23017 27897 23029 27900
rect 23063 27897 23075 27931
rect 23017 27891 23075 27897
rect 23109 27931 23167 27937
rect 23109 27897 23121 27931
rect 23155 27928 23167 27931
rect 23474 27928 23480 27940
rect 23155 27900 23480 27928
rect 23155 27897 23167 27900
rect 23109 27891 23167 27897
rect 23474 27888 23480 27900
rect 23532 27888 23538 27940
rect 24964 27937 24992 27968
rect 25041 27965 25053 27999
rect 25087 27996 25099 27999
rect 25682 27996 25688 28008
rect 25087 27968 25688 27996
rect 25087 27965 25099 27968
rect 25041 27959 25099 27965
rect 25682 27956 25688 27968
rect 25740 27956 25746 28008
rect 25976 27996 26004 28036
rect 26050 28024 26056 28076
rect 26108 28064 26114 28076
rect 26108 28036 26464 28064
rect 26108 28024 26114 28036
rect 26142 27996 26148 28008
rect 25976 27968 26148 27996
rect 26142 27956 26148 27968
rect 26200 27956 26206 28008
rect 26237 27999 26295 28005
rect 26237 27965 26249 27999
rect 26283 27996 26295 27999
rect 26326 27996 26332 28008
rect 26283 27968 26332 27996
rect 26283 27965 26295 27968
rect 26237 27959 26295 27965
rect 26326 27956 26332 27968
rect 26384 27956 26390 28008
rect 26436 28005 26464 28036
rect 26421 27999 26479 28005
rect 26421 27965 26433 27999
rect 26467 27965 26479 27999
rect 26421 27959 26479 27965
rect 26513 27999 26571 28005
rect 26513 27965 26525 27999
rect 26559 27996 26571 27999
rect 27338 27996 27344 28008
rect 26559 27968 27344 27996
rect 26559 27965 26571 27968
rect 26513 27959 26571 27965
rect 27338 27956 27344 27968
rect 27396 27956 27402 28008
rect 27801 27999 27859 28005
rect 27801 27965 27813 27999
rect 27847 27965 27859 27999
rect 28074 27996 28080 28008
rect 28035 27968 28080 27996
rect 27801 27959 27859 27965
rect 24949 27931 25007 27937
rect 24949 27897 24961 27931
rect 24995 27928 25007 27931
rect 26050 27928 26056 27940
rect 24995 27900 26056 27928
rect 24995 27897 25007 27900
rect 24949 27891 25007 27897
rect 26050 27888 26056 27900
rect 26108 27928 26114 27940
rect 27816 27928 27844 27959
rect 28074 27956 28080 27968
rect 28132 27956 28138 28008
rect 28169 27999 28227 28005
rect 28169 27965 28181 27999
rect 28215 27965 28227 27999
rect 28169 27959 28227 27965
rect 29089 27999 29147 28005
rect 29089 27965 29101 27999
rect 29135 27996 29147 27999
rect 30374 27996 30380 28008
rect 29135 27968 30380 27996
rect 29135 27965 29147 27968
rect 29089 27959 29147 27965
rect 27982 27928 27988 27940
rect 26108 27900 27844 27928
rect 27943 27900 27988 27928
rect 26108 27888 26114 27900
rect 27982 27888 27988 27900
rect 28040 27888 28046 27940
rect 25314 27860 25320 27872
rect 20916 27832 25320 27860
rect 25314 27820 25320 27832
rect 25372 27820 25378 27872
rect 26142 27820 26148 27872
rect 26200 27860 26206 27872
rect 28184 27860 28212 27959
rect 30374 27956 30380 27968
rect 30432 27956 30438 28008
rect 30834 27956 30840 28008
rect 30892 27996 30898 28008
rect 31128 28005 31156 28172
rect 31202 28092 31208 28144
rect 31260 28132 31266 28144
rect 31260 28104 31340 28132
rect 31260 28092 31266 28104
rect 31312 28073 31340 28104
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28033 31355 28067
rect 31297 28027 31355 28033
rect 31389 28067 31447 28073
rect 31389 28033 31401 28067
rect 31435 28064 31447 28067
rect 31662 28064 31668 28076
rect 31435 28036 31668 28064
rect 31435 28033 31447 28036
rect 31389 28027 31447 28033
rect 31662 28024 31668 28036
rect 31720 28024 31726 28076
rect 31754 28024 31760 28076
rect 31812 28064 31818 28076
rect 33778 28064 33784 28076
rect 31812 28036 33272 28064
rect 33739 28036 33784 28064
rect 31812 28024 31818 28036
rect 31113 27999 31171 28005
rect 31113 27996 31125 27999
rect 30892 27968 31125 27996
rect 30892 27956 30898 27968
rect 31113 27965 31125 27968
rect 31159 27965 31171 27999
rect 31113 27959 31171 27965
rect 31202 27956 31208 28008
rect 31260 27996 31266 28008
rect 31260 27968 31305 27996
rect 31260 27956 31266 27968
rect 31478 27956 31484 28008
rect 31536 27996 31542 28008
rect 31573 27999 31631 28005
rect 31573 27996 31585 27999
rect 31536 27968 31585 27996
rect 31536 27956 31542 27968
rect 31573 27965 31585 27968
rect 31619 27965 31631 27999
rect 31573 27959 31631 27965
rect 32030 27956 32036 28008
rect 32088 27996 32094 28008
rect 33045 27999 33103 28005
rect 33045 27996 33057 27999
rect 32088 27968 33057 27996
rect 32088 27956 32094 27968
rect 33045 27965 33057 27968
rect 33091 27965 33103 27999
rect 33244 27996 33272 28036
rect 33778 28024 33784 28036
rect 33836 28024 33842 28076
rect 33689 27999 33747 28005
rect 33689 27996 33701 27999
rect 33244 27968 33701 27996
rect 33045 27959 33103 27965
rect 33689 27965 33701 27968
rect 33735 27965 33747 27999
rect 34330 27996 34336 28008
rect 34291 27968 34336 27996
rect 33689 27959 33747 27965
rect 34330 27956 34336 27968
rect 34388 27956 34394 28008
rect 34532 28005 34560 28172
rect 55306 28160 55312 28172
rect 55364 28160 55370 28212
rect 56226 28200 56232 28212
rect 56187 28172 56232 28200
rect 56226 28160 56232 28172
rect 56284 28160 56290 28212
rect 57241 28203 57299 28209
rect 57241 28169 57253 28203
rect 57287 28200 57299 28203
rect 57698 28200 57704 28212
rect 57287 28172 57704 28200
rect 57287 28169 57299 28172
rect 57241 28163 57299 28169
rect 57698 28160 57704 28172
rect 57756 28160 57762 28212
rect 35713 28067 35771 28073
rect 35713 28033 35725 28067
rect 35759 28064 35771 28067
rect 56778 28064 56784 28076
rect 35759 28036 56784 28064
rect 35759 28033 35771 28036
rect 35713 28027 35771 28033
rect 56778 28024 56784 28036
rect 56836 28024 56842 28076
rect 34517 27999 34575 28005
rect 34517 27965 34529 27999
rect 34563 27965 34575 27999
rect 35434 27996 35440 28008
rect 35395 27968 35440 27996
rect 34517 27959 34575 27965
rect 35434 27956 35440 27968
rect 35492 27956 35498 28008
rect 35526 27956 35532 28008
rect 35584 27996 35590 28008
rect 36262 27996 36268 28008
rect 35584 27968 35629 27996
rect 36223 27968 36268 27996
rect 35584 27956 35590 27968
rect 36262 27956 36268 27968
rect 36320 27956 36326 28008
rect 36357 27999 36415 28005
rect 36357 27965 36369 27999
rect 36403 27965 36415 27999
rect 36357 27959 36415 27965
rect 29356 27931 29414 27937
rect 29356 27897 29368 27931
rect 29402 27928 29414 27931
rect 34425 27931 34483 27937
rect 34425 27928 34437 27931
rect 29402 27900 34437 27928
rect 29402 27897 29414 27900
rect 29356 27891 29414 27897
rect 34425 27897 34437 27900
rect 34471 27897 34483 27931
rect 34425 27891 34483 27897
rect 34606 27888 34612 27940
rect 34664 27928 34670 27940
rect 36372 27928 36400 27959
rect 55214 27956 55220 28008
rect 55272 27996 55278 28008
rect 55493 27999 55551 28005
rect 55493 27996 55505 27999
rect 55272 27968 55505 27996
rect 55272 27956 55278 27968
rect 55493 27965 55505 27968
rect 55539 27996 55551 27999
rect 56413 27999 56471 28005
rect 56413 27996 56425 27999
rect 55539 27968 56425 27996
rect 55539 27965 55551 27968
rect 55493 27959 55551 27965
rect 56413 27965 56425 27968
rect 56459 27965 56471 27999
rect 57422 27996 57428 28008
rect 57383 27968 57428 27996
rect 56413 27959 56471 27965
rect 57422 27956 57428 27968
rect 57480 27956 57486 28008
rect 34664 27900 36400 27928
rect 36541 27931 36599 27937
rect 34664 27888 34670 27900
rect 36541 27897 36553 27931
rect 36587 27928 36599 27931
rect 55122 27928 55128 27940
rect 36587 27900 55128 27928
rect 36587 27897 36599 27900
rect 36541 27891 36599 27897
rect 55122 27888 55128 27900
rect 55180 27888 55186 27940
rect 57974 27928 57980 27940
rect 57935 27900 57980 27928
rect 57974 27888 57980 27900
rect 58032 27888 58038 27940
rect 58158 27928 58164 27940
rect 58119 27900 58164 27928
rect 58158 27888 58164 27900
rect 58216 27888 58222 27940
rect 29086 27860 29092 27872
rect 26200 27832 29092 27860
rect 26200 27820 26206 27832
rect 29086 27820 29092 27832
rect 29144 27860 29150 27872
rect 30282 27860 30288 27872
rect 29144 27832 30288 27860
rect 29144 27820 29150 27832
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 30374 27820 30380 27872
rect 30432 27860 30438 27872
rect 30469 27863 30527 27869
rect 30469 27860 30481 27863
rect 30432 27832 30481 27860
rect 30432 27820 30438 27832
rect 30469 27829 30481 27832
rect 30515 27829 30527 27863
rect 30926 27860 30932 27872
rect 30887 27832 30932 27860
rect 30469 27823 30527 27829
rect 30926 27820 30932 27832
rect 30984 27820 30990 27872
rect 31478 27820 31484 27872
rect 31536 27860 31542 27872
rect 31662 27860 31668 27872
rect 31536 27832 31668 27860
rect 31536 27820 31542 27832
rect 31662 27820 31668 27832
rect 31720 27820 31726 27872
rect 31938 27820 31944 27872
rect 31996 27860 32002 27872
rect 33137 27863 33195 27869
rect 33137 27860 33149 27863
rect 31996 27832 33149 27860
rect 31996 27820 32002 27832
rect 33137 27829 33149 27832
rect 33183 27829 33195 27863
rect 33137 27823 33195 27829
rect 1104 27770 58880 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 50326 27770
rect 50378 27718 50390 27770
rect 50442 27718 50454 27770
rect 50506 27718 50518 27770
rect 50570 27718 58880 27770
rect 1104 27696 58880 27718
rect 1670 27616 1676 27668
rect 1728 27656 1734 27668
rect 2501 27659 2559 27665
rect 2501 27656 2513 27659
rect 1728 27628 2513 27656
rect 1728 27616 1734 27628
rect 2501 27625 2513 27628
rect 2547 27625 2559 27659
rect 2501 27619 2559 27625
rect 2774 27616 2780 27668
rect 2832 27656 2838 27668
rect 3145 27659 3203 27665
rect 3145 27656 3157 27659
rect 2832 27628 3157 27656
rect 2832 27616 2838 27628
rect 3145 27625 3157 27628
rect 3191 27625 3203 27659
rect 3145 27619 3203 27625
rect 5276 27628 5580 27656
rect 5276 27588 5304 27628
rect 5442 27588 5448 27600
rect 4632 27560 5304 27588
rect 5403 27560 5448 27588
rect 1857 27523 1915 27529
rect 1857 27489 1869 27523
rect 1903 27520 1915 27523
rect 2498 27520 2504 27532
rect 1903 27492 2504 27520
rect 1903 27489 1915 27492
rect 1857 27483 1915 27489
rect 2498 27480 2504 27492
rect 2556 27480 2562 27532
rect 2685 27523 2743 27529
rect 2685 27489 2697 27523
rect 2731 27520 2743 27523
rect 3326 27520 3332 27532
rect 2731 27492 3332 27520
rect 2731 27489 2743 27492
rect 2685 27483 2743 27489
rect 3326 27480 3332 27492
rect 3384 27480 3390 27532
rect 4632 27529 4660 27560
rect 5442 27548 5448 27560
rect 5500 27548 5506 27600
rect 5552 27588 5580 27628
rect 7006 27616 7012 27668
rect 7064 27656 7070 27668
rect 7193 27659 7251 27665
rect 7193 27656 7205 27659
rect 7064 27628 7205 27656
rect 7064 27616 7070 27628
rect 7193 27625 7205 27628
rect 7239 27625 7251 27659
rect 7193 27619 7251 27625
rect 12434 27616 12440 27668
rect 12492 27656 12498 27668
rect 13722 27656 13728 27668
rect 12492 27628 13728 27656
rect 12492 27616 12498 27628
rect 13722 27616 13728 27628
rect 13780 27616 13786 27668
rect 16206 27616 16212 27668
rect 16264 27656 16270 27668
rect 16485 27659 16543 27665
rect 16485 27656 16497 27659
rect 16264 27628 16497 27656
rect 16264 27616 16270 27628
rect 16485 27625 16497 27628
rect 16531 27656 16543 27659
rect 18598 27656 18604 27668
rect 16531 27628 18604 27656
rect 16531 27625 16543 27628
rect 16485 27619 16543 27625
rect 18598 27616 18604 27628
rect 18656 27616 18662 27668
rect 18874 27616 18880 27668
rect 18932 27656 18938 27668
rect 20990 27656 20996 27668
rect 18932 27628 20996 27656
rect 18932 27616 18938 27628
rect 20990 27616 20996 27628
rect 21048 27616 21054 27668
rect 21174 27616 21180 27668
rect 21232 27656 21238 27668
rect 26878 27656 26884 27668
rect 21232 27628 26884 27656
rect 21232 27616 21238 27628
rect 9490 27588 9496 27600
rect 5552 27560 9496 27588
rect 9490 27548 9496 27560
rect 9548 27548 9554 27600
rect 9858 27548 9864 27600
rect 9916 27588 9922 27600
rect 9916 27560 10180 27588
rect 9916 27548 9922 27560
rect 4617 27523 4675 27529
rect 4617 27489 4629 27523
rect 4663 27489 4675 27523
rect 4617 27483 4675 27489
rect 7377 27523 7435 27529
rect 7377 27489 7389 27523
rect 7423 27489 7435 27523
rect 7377 27483 7435 27489
rect 7469 27523 7527 27529
rect 7469 27489 7481 27523
rect 7515 27520 7527 27523
rect 7558 27520 7564 27532
rect 7515 27492 7564 27520
rect 7515 27489 7527 27492
rect 7469 27483 7527 27489
rect 5353 27455 5411 27461
rect 5353 27421 5365 27455
rect 5399 27452 5411 27455
rect 5626 27452 5632 27464
rect 5399 27424 5632 27452
rect 5399 27421 5411 27424
rect 5353 27415 5411 27421
rect 5626 27412 5632 27424
rect 5684 27412 5690 27464
rect 6365 27455 6423 27461
rect 6365 27421 6377 27455
rect 6411 27452 6423 27455
rect 6454 27452 6460 27464
rect 6411 27424 6460 27452
rect 6411 27421 6423 27424
rect 6365 27415 6423 27421
rect 6454 27412 6460 27424
rect 6512 27412 6518 27464
rect 7392 27384 7420 27483
rect 7558 27480 7564 27492
rect 7616 27480 7622 27532
rect 7742 27520 7748 27532
rect 7703 27492 7748 27520
rect 7742 27480 7748 27492
rect 7800 27480 7806 27532
rect 8297 27523 8355 27529
rect 8297 27489 8309 27523
rect 8343 27520 8355 27523
rect 8386 27520 8392 27532
rect 8343 27492 8392 27520
rect 8343 27489 8355 27492
rect 8297 27483 8355 27489
rect 8386 27480 8392 27492
rect 8444 27480 8450 27532
rect 9674 27520 9680 27532
rect 9635 27492 9680 27520
rect 9674 27480 9680 27492
rect 9732 27480 9738 27532
rect 9766 27480 9772 27532
rect 9824 27520 9830 27532
rect 10042 27520 10048 27532
rect 9824 27492 9869 27520
rect 10003 27492 10048 27520
rect 9824 27480 9830 27492
rect 10042 27480 10048 27492
rect 10100 27480 10106 27532
rect 10152 27520 10180 27560
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 11020 27560 15240 27588
rect 11020 27548 11026 27560
rect 11057 27523 11115 27529
rect 11057 27520 11069 27523
rect 10152 27492 11069 27520
rect 11057 27489 11069 27492
rect 11103 27489 11115 27523
rect 11057 27483 11115 27489
rect 11146 27480 11152 27532
rect 11204 27520 11210 27532
rect 11313 27523 11371 27529
rect 11313 27520 11325 27523
rect 11204 27492 11325 27520
rect 11204 27480 11210 27492
rect 11313 27489 11325 27492
rect 11359 27489 11371 27523
rect 11313 27483 11371 27489
rect 13449 27523 13507 27529
rect 13449 27489 13461 27523
rect 13495 27520 13507 27523
rect 14642 27520 14648 27532
rect 13495 27492 14648 27520
rect 13495 27489 13507 27492
rect 13449 27483 13507 27489
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 8110 27452 8116 27464
rect 7699 27424 8116 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 8110 27412 8116 27424
rect 8168 27412 8174 27464
rect 9950 27452 9956 27464
rect 9600 27424 9812 27452
rect 9911 27424 9956 27452
rect 9600 27384 9628 27424
rect 7392 27356 9628 27384
rect 9784 27384 9812 27424
rect 9950 27412 9956 27424
rect 10008 27412 10014 27464
rect 12618 27412 12624 27464
rect 12676 27452 12682 27464
rect 13722 27452 13728 27464
rect 12676 27424 13728 27452
rect 12676 27412 12682 27424
rect 13722 27412 13728 27424
rect 13780 27412 13786 27464
rect 15212 27461 15240 27560
rect 15470 27548 15476 27600
rect 15528 27588 15534 27600
rect 20257 27591 20315 27597
rect 15528 27560 20116 27588
rect 15528 27548 15534 27560
rect 15378 27520 15384 27532
rect 15339 27492 15384 27520
rect 15378 27480 15384 27492
rect 15436 27480 15442 27532
rect 15562 27520 15568 27532
rect 15523 27492 15568 27520
rect 15562 27480 15568 27492
rect 15620 27480 15626 27532
rect 15841 27523 15899 27529
rect 15841 27489 15853 27523
rect 15887 27489 15899 27523
rect 15841 27483 15899 27489
rect 16301 27523 16359 27529
rect 16301 27489 16313 27523
rect 16347 27489 16359 27523
rect 16301 27483 16359 27489
rect 16577 27523 16635 27529
rect 16577 27489 16589 27523
rect 16623 27520 16635 27523
rect 17034 27520 17040 27532
rect 16623 27492 17040 27520
rect 16623 27489 16635 27492
rect 16577 27483 16635 27489
rect 15197 27455 15255 27461
rect 15197 27421 15209 27455
rect 15243 27421 15255 27455
rect 15197 27415 15255 27421
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 15657 27455 15715 27461
rect 15657 27452 15669 27455
rect 15344 27424 15669 27452
rect 15344 27412 15350 27424
rect 15657 27421 15669 27424
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 9784 27356 11100 27384
rect 1394 27276 1400 27328
rect 1452 27316 1458 27328
rect 1949 27319 2007 27325
rect 1949 27316 1961 27319
rect 1452 27288 1961 27316
rect 1452 27276 1458 27288
rect 1949 27285 1961 27288
rect 1995 27285 2007 27319
rect 1949 27279 2007 27285
rect 4706 27276 4712 27328
rect 4764 27316 4770 27328
rect 4801 27319 4859 27325
rect 4801 27316 4813 27319
rect 4764 27288 4813 27316
rect 4764 27276 4770 27288
rect 4801 27285 4813 27288
rect 4847 27285 4859 27319
rect 4801 27279 4859 27285
rect 7282 27276 7288 27328
rect 7340 27316 7346 27328
rect 8202 27316 8208 27328
rect 7340 27288 8208 27316
rect 7340 27276 7346 27288
rect 8202 27276 8208 27288
rect 8260 27316 8266 27328
rect 8389 27319 8447 27325
rect 8389 27316 8401 27319
rect 8260 27288 8401 27316
rect 8260 27276 8266 27288
rect 8389 27285 8401 27288
rect 8435 27285 8447 27319
rect 9490 27316 9496 27328
rect 9451 27288 9496 27316
rect 8389 27279 8447 27285
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 9674 27276 9680 27328
rect 9732 27316 9738 27328
rect 10962 27316 10968 27328
rect 9732 27288 10968 27316
rect 9732 27276 9738 27288
rect 10962 27276 10968 27288
rect 11020 27276 11026 27328
rect 11072 27316 11100 27356
rect 12526 27344 12532 27396
rect 12584 27384 12590 27396
rect 13633 27387 13691 27393
rect 13633 27384 13645 27387
rect 12584 27356 13645 27384
rect 12584 27344 12590 27356
rect 13633 27353 13645 27356
rect 13679 27353 13691 27387
rect 13633 27347 13691 27353
rect 13814 27344 13820 27396
rect 13872 27384 13878 27396
rect 15304 27384 15332 27412
rect 15470 27384 15476 27396
rect 13872 27356 15332 27384
rect 15431 27356 15476 27384
rect 13872 27344 13878 27356
rect 15470 27344 15476 27356
rect 15528 27344 15534 27396
rect 12250 27316 12256 27328
rect 11072 27288 12256 27316
rect 12250 27276 12256 27288
rect 12308 27276 12314 27328
rect 12342 27276 12348 27328
rect 12400 27316 12406 27328
rect 12437 27319 12495 27325
rect 12437 27316 12449 27319
rect 12400 27288 12449 27316
rect 12400 27276 12406 27288
rect 12437 27285 12449 27288
rect 12483 27285 12495 27319
rect 13538 27316 13544 27328
rect 13499 27288 13544 27316
rect 12437 27279 12495 27285
rect 13538 27276 13544 27288
rect 13596 27276 13602 27328
rect 14550 27276 14556 27328
rect 14608 27316 14614 27328
rect 15856 27316 15884 27483
rect 16316 27452 16344 27483
rect 17034 27480 17040 27492
rect 17092 27480 17098 27532
rect 17402 27529 17408 27532
rect 17221 27523 17279 27529
rect 17221 27489 17233 27523
rect 17267 27489 17279 27523
rect 17221 27483 17279 27489
rect 17359 27523 17408 27529
rect 17359 27489 17371 27523
rect 17405 27489 17408 27523
rect 17359 27483 17408 27489
rect 17126 27452 17132 27464
rect 16316 27424 17132 27452
rect 17126 27412 17132 27424
rect 17184 27412 17190 27464
rect 16301 27387 16359 27393
rect 16301 27353 16313 27387
rect 16347 27384 16359 27387
rect 16482 27384 16488 27396
rect 16347 27356 16488 27384
rect 16347 27353 16359 27356
rect 16301 27347 16359 27353
rect 16482 27344 16488 27356
rect 16540 27344 16546 27396
rect 17236 27384 17264 27483
rect 17402 27480 17408 27483
rect 17460 27480 17466 27532
rect 17586 27520 17592 27532
rect 17547 27492 17592 27520
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 18046 27520 18052 27532
rect 17696 27492 18052 27520
rect 17696 27452 17724 27492
rect 18046 27480 18052 27492
rect 18104 27520 18110 27532
rect 18233 27523 18291 27529
rect 18233 27520 18245 27523
rect 18104 27492 18245 27520
rect 18104 27480 18110 27492
rect 18233 27489 18245 27492
rect 18279 27489 18291 27523
rect 18233 27483 18291 27489
rect 18417 27523 18475 27529
rect 18417 27489 18429 27523
rect 18463 27520 18475 27523
rect 18598 27520 18604 27532
rect 18463 27492 18604 27520
rect 18463 27489 18475 27492
rect 18417 27483 18475 27489
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 20088 27529 20116 27560
rect 20257 27557 20269 27591
rect 20303 27588 20315 27591
rect 22278 27588 22284 27600
rect 20303 27560 22284 27588
rect 20303 27557 20315 27560
rect 20257 27551 20315 27557
rect 22278 27548 22284 27560
rect 22336 27548 22342 27600
rect 22480 27597 22508 27628
rect 26878 27616 26884 27628
rect 26936 27616 26942 27668
rect 29086 27656 29092 27668
rect 29047 27628 29092 27656
rect 29086 27616 29092 27628
rect 29144 27616 29150 27668
rect 34606 27656 34612 27668
rect 31864 27628 34612 27656
rect 22465 27591 22523 27597
rect 22465 27557 22477 27591
rect 22511 27557 22523 27591
rect 23566 27588 23572 27600
rect 22465 27551 22523 27557
rect 22664 27560 23572 27588
rect 19981 27523 20039 27529
rect 19981 27489 19993 27523
rect 20027 27489 20039 27523
rect 19981 27483 20039 27489
rect 20074 27523 20132 27529
rect 20074 27489 20086 27523
rect 20120 27489 20132 27523
rect 20074 27483 20132 27489
rect 17420 27424 17724 27452
rect 17420 27384 17448 27424
rect 17862 27412 17868 27464
rect 17920 27452 17926 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 17920 27424 18337 27452
rect 17920 27412 17926 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18506 27452 18512 27464
rect 18467 27424 18512 27452
rect 18325 27415 18383 27421
rect 18506 27412 18512 27424
rect 18564 27412 18570 27464
rect 19996 27452 20024 27483
rect 20162 27480 20168 27532
rect 20220 27520 20226 27532
rect 20349 27523 20407 27529
rect 20349 27520 20361 27523
rect 20220 27492 20361 27520
rect 20220 27480 20226 27492
rect 20349 27489 20361 27492
rect 20395 27489 20407 27523
rect 20349 27483 20407 27489
rect 20438 27480 20444 27532
rect 20496 27529 20502 27532
rect 20496 27520 20504 27529
rect 21174 27520 21180 27532
rect 20496 27492 20541 27520
rect 21135 27492 21180 27520
rect 20496 27483 20504 27492
rect 20496 27480 20502 27483
rect 21174 27480 21180 27492
rect 21232 27480 21238 27532
rect 21358 27520 21364 27532
rect 21319 27492 21364 27520
rect 21358 27480 21364 27492
rect 21416 27480 21422 27532
rect 21821 27523 21879 27529
rect 21821 27489 21833 27523
rect 21867 27489 21879 27523
rect 21821 27483 21879 27489
rect 21266 27452 21272 27464
rect 19306 27424 20760 27452
rect 21227 27424 21272 27452
rect 16592 27356 17172 27384
rect 17236 27356 17448 27384
rect 17497 27387 17555 27393
rect 14608 27288 15884 27316
rect 14608 27276 14614 27288
rect 16114 27276 16120 27328
rect 16172 27316 16178 27328
rect 16592 27316 16620 27356
rect 17034 27316 17040 27328
rect 16172 27288 16620 27316
rect 16995 27288 17040 27316
rect 16172 27276 16178 27288
rect 17034 27276 17040 27288
rect 17092 27276 17098 27328
rect 17144 27316 17172 27356
rect 17497 27353 17509 27387
rect 17543 27384 17555 27387
rect 17586 27384 17592 27396
rect 17543 27356 17592 27384
rect 17543 27353 17555 27356
rect 17497 27347 17555 27353
rect 17586 27344 17592 27356
rect 17644 27344 17650 27396
rect 19306 27384 19334 27424
rect 17696 27356 19334 27384
rect 17696 27316 17724 27356
rect 18046 27316 18052 27328
rect 17144 27288 17724 27316
rect 18007 27288 18052 27316
rect 18046 27276 18052 27288
rect 18104 27276 18110 27328
rect 18138 27276 18144 27328
rect 18196 27316 18202 27328
rect 20438 27316 20444 27328
rect 18196 27288 20444 27316
rect 18196 27276 18202 27288
rect 20438 27276 20444 27288
rect 20496 27276 20502 27328
rect 20622 27316 20628 27328
rect 20583 27288 20628 27316
rect 20622 27276 20628 27288
rect 20680 27276 20686 27328
rect 20732 27316 20760 27424
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 21836 27452 21864 27483
rect 22002 27480 22008 27532
rect 22060 27520 22066 27532
rect 22664 27529 22692 27560
rect 23566 27548 23572 27560
rect 23624 27548 23630 27600
rect 24213 27591 24271 27597
rect 24213 27557 24225 27591
rect 24259 27588 24271 27591
rect 24762 27588 24768 27600
rect 24259 27560 24768 27588
rect 24259 27557 24271 27560
rect 24213 27551 24271 27557
rect 22649 27523 22707 27529
rect 22649 27520 22661 27523
rect 22060 27492 22661 27520
rect 22060 27480 22066 27492
rect 22649 27489 22661 27492
rect 22695 27489 22707 27523
rect 22649 27483 22707 27489
rect 22741 27523 22799 27529
rect 22741 27489 22753 27523
rect 22787 27520 22799 27523
rect 23017 27523 23075 27529
rect 22787 27492 22867 27520
rect 22787 27489 22799 27492
rect 22741 27483 22799 27489
rect 21376 27424 21864 27452
rect 21174 27344 21180 27396
rect 21232 27384 21238 27396
rect 21376 27384 21404 27424
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 21968 27424 22013 27452
rect 21968 27412 21974 27424
rect 21232 27356 21404 27384
rect 21232 27344 21238 27356
rect 21450 27344 21456 27396
rect 21508 27384 21514 27396
rect 22839 27384 22867 27492
rect 23017 27489 23029 27523
rect 23063 27520 23075 27523
rect 23474 27520 23480 27532
rect 23063 27492 23480 27520
rect 23063 27489 23075 27492
rect 23017 27483 23075 27489
rect 23474 27480 23480 27492
rect 23532 27480 23538 27532
rect 24118 27520 24124 27532
rect 24079 27492 24124 27520
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 23198 27452 23204 27464
rect 22971 27424 23204 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 23198 27412 23204 27424
rect 23256 27452 23262 27464
rect 24136 27452 24164 27480
rect 23256 27424 24164 27452
rect 23256 27412 23262 27424
rect 24228 27384 24256 27551
rect 24762 27548 24768 27560
rect 24820 27548 24826 27600
rect 26053 27591 26111 27597
rect 26053 27557 26065 27591
rect 26099 27588 26111 27591
rect 27982 27588 27988 27600
rect 26099 27560 27988 27588
rect 26099 27557 26111 27560
rect 26053 27551 26111 27557
rect 27982 27548 27988 27560
rect 28040 27548 28046 27600
rect 30374 27548 30380 27600
rect 30432 27588 30438 27600
rect 30432 27560 31616 27588
rect 30432 27548 30438 27560
rect 25685 27523 25743 27529
rect 25685 27489 25697 27523
rect 25731 27489 25743 27523
rect 25685 27483 25743 27489
rect 25869 27523 25927 27529
rect 25869 27489 25881 27523
rect 25915 27520 25927 27523
rect 26142 27520 26148 27532
rect 25915 27492 26148 27520
rect 25915 27489 25927 27492
rect 25869 27483 25927 27489
rect 25700 27452 25728 27483
rect 26142 27480 26148 27492
rect 26200 27520 26206 27532
rect 26513 27523 26571 27529
rect 26513 27520 26525 27523
rect 26200 27492 26525 27520
rect 26200 27480 26206 27492
rect 26513 27489 26525 27492
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 26602 27480 26608 27532
rect 26660 27520 26666 27532
rect 27430 27529 27436 27532
rect 27424 27520 27436 27529
rect 26660 27492 26705 27520
rect 27391 27492 27436 27520
rect 26660 27480 26666 27492
rect 27424 27483 27436 27492
rect 27430 27480 27436 27483
rect 27488 27480 27494 27532
rect 28997 27523 29055 27529
rect 28997 27520 29009 27523
rect 28552 27492 29009 27520
rect 25700 27424 27108 27452
rect 25682 27384 25688 27396
rect 21508 27356 24256 27384
rect 25643 27356 25688 27384
rect 21508 27344 21514 27356
rect 25682 27344 25688 27356
rect 25740 27344 25746 27396
rect 25866 27344 25872 27396
rect 25924 27384 25930 27396
rect 26418 27384 26424 27396
rect 25924 27356 26424 27384
rect 25924 27344 25930 27356
rect 26418 27344 26424 27356
rect 26476 27344 26482 27396
rect 25958 27316 25964 27328
rect 20732 27288 25964 27316
rect 25958 27276 25964 27288
rect 26016 27276 26022 27328
rect 27080 27316 27108 27424
rect 27154 27412 27160 27464
rect 27212 27452 27218 27464
rect 27212 27424 27257 27452
rect 27212 27412 27218 27424
rect 28552 27325 28580 27492
rect 28997 27489 29009 27492
rect 29043 27489 29055 27523
rect 28997 27483 29055 27489
rect 30190 27480 30196 27532
rect 30248 27520 30254 27532
rect 30834 27520 30840 27532
rect 30248 27492 30840 27520
rect 30248 27480 30254 27492
rect 30834 27480 30840 27492
rect 30892 27480 30898 27532
rect 31588 27529 31616 27560
rect 31662 27548 31668 27600
rect 31720 27588 31726 27600
rect 31864 27588 31892 27628
rect 34606 27616 34612 27628
rect 34664 27616 34670 27668
rect 57974 27616 57980 27668
rect 58032 27656 58038 27668
rect 58161 27659 58219 27665
rect 58161 27656 58173 27659
rect 58032 27628 58173 27656
rect 58032 27616 58038 27628
rect 58161 27625 58173 27628
rect 58207 27625 58219 27659
rect 58161 27619 58219 27625
rect 31720 27560 31892 27588
rect 31720 27548 31726 27560
rect 31573 27523 31631 27529
rect 31573 27489 31585 27523
rect 31619 27489 31631 27523
rect 31573 27483 31631 27489
rect 32585 27523 32643 27529
rect 32585 27489 32597 27523
rect 32631 27520 32643 27523
rect 32950 27520 32956 27532
rect 32631 27492 32956 27520
rect 32631 27489 32643 27492
rect 32585 27483 32643 27489
rect 32950 27480 32956 27492
rect 33008 27480 33014 27532
rect 33042 27480 33048 27532
rect 33100 27520 33106 27532
rect 33669 27523 33727 27529
rect 33669 27520 33681 27523
rect 33100 27492 33681 27520
rect 33100 27480 33106 27492
rect 33669 27489 33681 27492
rect 33715 27489 33727 27523
rect 35710 27520 35716 27532
rect 35671 27492 35716 27520
rect 33669 27483 33727 27489
rect 35710 27480 35716 27492
rect 35768 27480 35774 27532
rect 55582 27520 55588 27532
rect 55543 27492 55588 27520
rect 55582 27480 55588 27492
rect 55640 27480 55646 27532
rect 56042 27480 56048 27532
rect 56100 27520 56106 27532
rect 56873 27523 56931 27529
rect 56873 27520 56885 27523
rect 56100 27492 56885 27520
rect 56100 27480 56106 27492
rect 56873 27489 56885 27492
rect 56919 27489 56931 27523
rect 56873 27483 56931 27489
rect 31113 27455 31171 27461
rect 31113 27421 31125 27455
rect 31159 27452 31171 27455
rect 32030 27452 32036 27464
rect 31159 27424 32036 27452
rect 31159 27421 31171 27424
rect 31113 27415 31171 27421
rect 32030 27412 32036 27424
rect 32088 27412 32094 27464
rect 32858 27412 32864 27464
rect 32916 27452 32922 27464
rect 33410 27452 33416 27464
rect 32916 27424 33416 27452
rect 32916 27412 32922 27424
rect 33410 27412 33416 27424
rect 33468 27412 33474 27464
rect 56778 27412 56784 27464
rect 56836 27452 56842 27464
rect 57517 27455 57575 27461
rect 57517 27452 57529 27455
rect 56836 27424 57529 27452
rect 56836 27412 56842 27424
rect 57517 27421 57529 27424
rect 57563 27421 57575 27455
rect 57698 27452 57704 27464
rect 57659 27424 57704 27452
rect 57517 27415 57575 27421
rect 57698 27412 57704 27424
rect 57756 27412 57762 27464
rect 31021 27387 31079 27393
rect 31021 27353 31033 27387
rect 31067 27384 31079 27387
rect 31754 27384 31760 27396
rect 31067 27356 31760 27384
rect 31067 27353 31079 27356
rect 31021 27347 31079 27353
rect 31754 27344 31760 27356
rect 31812 27344 31818 27396
rect 28537 27319 28595 27325
rect 28537 27316 28549 27319
rect 27080 27288 28549 27316
rect 28537 27285 28549 27288
rect 28583 27285 28595 27319
rect 28537 27279 28595 27285
rect 30006 27276 30012 27328
rect 30064 27316 30070 27328
rect 30929 27319 30987 27325
rect 30929 27316 30941 27319
rect 30064 27288 30941 27316
rect 30064 27276 30070 27288
rect 30929 27285 30941 27288
rect 30975 27316 30987 27319
rect 31202 27316 31208 27328
rect 30975 27288 31208 27316
rect 30975 27285 30987 27288
rect 30929 27279 30987 27285
rect 31202 27276 31208 27288
rect 31260 27316 31266 27328
rect 31662 27316 31668 27328
rect 31260 27288 31668 27316
rect 31260 27276 31266 27288
rect 31662 27276 31668 27288
rect 31720 27276 31726 27328
rect 32677 27319 32735 27325
rect 32677 27285 32689 27319
rect 32723 27316 32735 27319
rect 32858 27316 32864 27328
rect 32723 27288 32864 27316
rect 32723 27285 32735 27288
rect 32677 27279 32735 27285
rect 32858 27276 32864 27288
rect 32916 27276 32922 27328
rect 34790 27316 34796 27328
rect 34751 27288 34796 27316
rect 34790 27276 34796 27288
rect 34848 27276 34854 27328
rect 35897 27319 35955 27325
rect 35897 27285 35909 27319
rect 35943 27316 35955 27319
rect 36354 27316 36360 27328
rect 35943 27288 36360 27316
rect 35943 27285 35955 27288
rect 35897 27279 35955 27285
rect 36354 27276 36360 27288
rect 36412 27276 36418 27328
rect 56962 27316 56968 27328
rect 56923 27288 56968 27316
rect 56962 27276 56968 27288
rect 57020 27276 57026 27328
rect 1104 27226 58880 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 58880 27226
rect 1104 27152 58880 27174
rect 1854 27112 1860 27124
rect 1815 27084 1860 27112
rect 1854 27072 1860 27084
rect 1912 27072 1918 27124
rect 5442 27112 5448 27124
rect 5403 27084 5448 27112
rect 5442 27072 5448 27084
rect 5500 27072 5506 27124
rect 5626 27072 5632 27124
rect 5684 27112 5690 27124
rect 10410 27112 10416 27124
rect 5684 27084 10416 27112
rect 5684 27072 5690 27084
rect 10410 27072 10416 27084
rect 10468 27072 10474 27124
rect 11146 27112 11152 27124
rect 11107 27084 11152 27112
rect 11146 27072 11152 27084
rect 11204 27072 11210 27124
rect 14090 27112 14096 27124
rect 11532 27084 14096 27112
rect 2593 27047 2651 27053
rect 2593 27044 2605 27047
rect 1688 27016 2605 27044
rect 1688 26985 1716 27016
rect 2593 27013 2605 27016
rect 2639 27013 2651 27047
rect 2593 27007 2651 27013
rect 8110 27004 8116 27056
rect 8168 27044 8174 27056
rect 8941 27047 8999 27053
rect 8941 27044 8953 27047
rect 8168 27016 8953 27044
rect 8168 27004 8174 27016
rect 8941 27013 8953 27016
rect 8987 27044 8999 27047
rect 9950 27044 9956 27056
rect 8987 27016 9956 27044
rect 8987 27013 8999 27016
rect 8941 27007 8999 27013
rect 9950 27004 9956 27016
rect 10008 27004 10014 27056
rect 11238 27044 11244 27056
rect 10612 27016 11244 27044
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26945 1731 26979
rect 3326 26976 3332 26988
rect 1673 26939 1731 26945
rect 2792 26948 3332 26976
rect 2792 26917 2820 26948
rect 3326 26936 3332 26948
rect 3384 26976 3390 26988
rect 5442 26976 5448 26988
rect 3384 26948 5448 26976
rect 3384 26936 3390 26948
rect 5442 26936 5448 26948
rect 5500 26936 5506 26988
rect 6822 26976 6828 26988
rect 6783 26948 6828 26976
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 7926 26936 7932 26988
rect 7984 26976 7990 26988
rect 9858 26976 9864 26988
rect 7984 26948 9864 26976
rect 7984 26936 7990 26948
rect 9858 26936 9864 26948
rect 9916 26936 9922 26988
rect 1489 26911 1547 26917
rect 1489 26877 1501 26911
rect 1535 26877 1547 26911
rect 1489 26871 1547 26877
rect 2777 26911 2835 26917
rect 2777 26877 2789 26911
rect 2823 26877 2835 26911
rect 3418 26908 3424 26920
rect 3331 26880 3424 26908
rect 2777 26871 2835 26877
rect 1504 26840 1532 26871
rect 3418 26868 3424 26880
rect 3476 26908 3482 26920
rect 4065 26911 4123 26917
rect 4065 26908 4077 26911
rect 3476 26880 4077 26908
rect 3476 26868 3482 26880
rect 4065 26877 4077 26880
rect 4111 26877 4123 26911
rect 4522 26908 4528 26920
rect 4483 26880 4528 26908
rect 4065 26871 4123 26877
rect 4522 26868 4528 26880
rect 4580 26868 4586 26920
rect 4706 26908 4712 26920
rect 4667 26880 4712 26908
rect 4706 26868 4712 26880
rect 4764 26868 4770 26920
rect 5258 26908 5264 26920
rect 5219 26880 5264 26908
rect 5258 26868 5264 26880
rect 5316 26908 5322 26920
rect 7098 26917 7104 26920
rect 7092 26908 7104 26917
rect 5316 26880 6960 26908
rect 7059 26880 7104 26908
rect 5316 26868 5322 26880
rect 5350 26840 5356 26852
rect 1504 26812 5356 26840
rect 5350 26800 5356 26812
rect 5408 26800 5414 26852
rect 6932 26840 6960 26880
rect 7092 26871 7104 26880
rect 7098 26868 7104 26871
rect 7156 26868 7162 26920
rect 8386 26868 8392 26920
rect 8444 26908 8450 26920
rect 10134 26908 10140 26920
rect 8444 26880 10140 26908
rect 8444 26868 8450 26880
rect 10134 26868 10140 26880
rect 10192 26868 10198 26920
rect 10410 26908 10416 26920
rect 10371 26880 10416 26908
rect 10410 26868 10416 26880
rect 10468 26868 10474 26920
rect 10612 26917 10640 27016
rect 11238 27004 11244 27016
rect 11296 27004 11302 27056
rect 10689 26979 10747 26985
rect 10689 26945 10701 26979
rect 10735 26976 10747 26979
rect 11532 26976 11560 27084
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 17310 27072 17316 27124
rect 17368 27112 17374 27124
rect 17862 27112 17868 27124
rect 17368 27084 17868 27112
rect 17368 27072 17374 27084
rect 17862 27072 17868 27084
rect 17920 27072 17926 27124
rect 17954 27072 17960 27124
rect 18012 27112 18018 27124
rect 21085 27115 21143 27121
rect 21085 27112 21097 27115
rect 18012 27084 21097 27112
rect 18012 27072 18018 27084
rect 21085 27081 21097 27084
rect 21131 27112 21143 27115
rect 21450 27112 21456 27124
rect 21131 27084 21456 27112
rect 21131 27081 21143 27084
rect 21085 27075 21143 27081
rect 21450 27072 21456 27084
rect 21508 27072 21514 27124
rect 24029 27115 24087 27121
rect 24029 27081 24041 27115
rect 24075 27112 24087 27115
rect 24118 27112 24124 27124
rect 24075 27084 24124 27112
rect 24075 27081 24087 27084
rect 24029 27075 24087 27081
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 24670 27112 24676 27124
rect 24631 27084 24676 27112
rect 24670 27072 24676 27084
rect 24728 27072 24734 27124
rect 25866 27112 25872 27124
rect 25332 27084 25872 27112
rect 11606 27004 11612 27056
rect 11664 27044 11670 27056
rect 12897 27047 12955 27053
rect 12897 27044 12909 27047
rect 11664 27016 12909 27044
rect 11664 27004 11670 27016
rect 12897 27013 12909 27016
rect 12943 27013 12955 27047
rect 14277 27047 14335 27053
rect 14277 27044 14289 27047
rect 12897 27007 12955 27013
rect 13280 27016 14289 27044
rect 12342 26976 12348 26988
rect 10735 26948 11560 26976
rect 11992 26948 12348 26976
rect 10735 26945 10747 26948
rect 10689 26939 10747 26945
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26877 10655 26911
rect 10597 26871 10655 26877
rect 10781 26911 10839 26917
rect 10781 26877 10793 26911
rect 10827 26877 10839 26911
rect 10781 26871 10839 26877
rect 8110 26840 8116 26852
rect 6932 26812 8116 26840
rect 8110 26800 8116 26812
rect 8168 26800 8174 26852
rect 8570 26800 8576 26852
rect 8628 26840 8634 26852
rect 8757 26843 8815 26849
rect 8757 26840 8769 26843
rect 8628 26812 8769 26840
rect 8628 26800 8634 26812
rect 8757 26809 8769 26812
rect 8803 26840 8815 26843
rect 9769 26843 9827 26849
rect 9769 26840 9781 26843
rect 8803 26812 9781 26840
rect 8803 26809 8815 26812
rect 8757 26803 8815 26809
rect 9769 26809 9781 26812
rect 9815 26809 9827 26843
rect 9769 26803 9827 26809
rect 9953 26843 10011 26849
rect 9953 26809 9965 26843
rect 9999 26840 10011 26843
rect 10226 26840 10232 26852
rect 9999 26812 10232 26840
rect 9999 26809 10011 26812
rect 9953 26803 10011 26809
rect 10226 26800 10232 26812
rect 10284 26840 10290 26852
rect 10796 26840 10824 26871
rect 10962 26868 10968 26920
rect 11020 26908 11026 26920
rect 11992 26908 12020 26948
rect 12342 26936 12348 26948
rect 12400 26936 12406 26988
rect 12618 26936 12624 26988
rect 12676 26976 12682 26988
rect 12989 26979 13047 26985
rect 12989 26976 13001 26979
rect 12676 26948 13001 26976
rect 12676 26936 12682 26948
rect 12989 26945 13001 26948
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 11020 26880 12020 26908
rect 12069 26911 12127 26917
rect 11020 26868 11026 26880
rect 12069 26877 12081 26911
rect 12115 26908 12127 26911
rect 12434 26908 12440 26920
rect 12115 26880 12440 26908
rect 12115 26877 12127 26880
rect 12069 26871 12127 26877
rect 12434 26868 12440 26880
rect 12492 26868 12498 26920
rect 12710 26908 12716 26920
rect 12671 26880 12716 26908
rect 12710 26868 12716 26880
rect 12768 26868 12774 26920
rect 12805 26911 12863 26917
rect 12805 26877 12817 26911
rect 12851 26908 12863 26911
rect 13280 26908 13308 27016
rect 12851 26880 13308 26908
rect 12851 26877 12863 26880
rect 12805 26871 12863 26877
rect 13354 26868 13360 26920
rect 13412 26908 13418 26920
rect 13449 26911 13507 26917
rect 13449 26908 13461 26911
rect 13412 26880 13461 26908
rect 13412 26868 13418 26880
rect 13449 26877 13461 26880
rect 13495 26877 13507 26911
rect 13449 26871 13507 26877
rect 13538 26868 13544 26920
rect 13596 26908 13602 26920
rect 13648 26908 13676 27016
rect 14277 27013 14289 27016
rect 14323 27044 14335 27047
rect 15105 27047 15163 27053
rect 15105 27044 15117 27047
rect 14323 27016 15117 27044
rect 14323 27013 14335 27016
rect 14277 27007 14335 27013
rect 15105 27013 15117 27016
rect 15151 27013 15163 27047
rect 15105 27007 15163 27013
rect 15470 27004 15476 27056
rect 15528 27044 15534 27056
rect 16301 27047 16359 27053
rect 16301 27044 16313 27047
rect 15528 27016 16313 27044
rect 15528 27004 15534 27016
rect 16301 27013 16313 27016
rect 16347 27044 16359 27047
rect 17770 27044 17776 27056
rect 16347 27016 17776 27044
rect 16347 27013 16359 27016
rect 16301 27007 16359 27013
rect 17770 27004 17776 27016
rect 17828 27004 17834 27056
rect 13728 26979 13786 26985
rect 13728 26945 13740 26979
rect 13774 26976 13786 26979
rect 13814 26976 13820 26988
rect 13774 26948 13820 26976
rect 13774 26945 13786 26948
rect 13728 26939 13786 26945
rect 13814 26936 13820 26948
rect 13872 26976 13878 26988
rect 14461 26979 14519 26985
rect 14461 26976 14473 26979
rect 13872 26948 14473 26976
rect 13872 26936 13878 26948
rect 14461 26945 14473 26948
rect 14507 26945 14519 26979
rect 14461 26939 14519 26945
rect 14642 26936 14648 26988
rect 14700 26976 14706 26988
rect 17034 26976 17040 26988
rect 14700 26948 17040 26976
rect 14700 26936 14706 26948
rect 17034 26936 17040 26948
rect 17092 26936 17098 26988
rect 17218 26936 17224 26988
rect 17276 26976 17282 26988
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 17276 26948 17325 26976
rect 17276 26936 17282 26948
rect 17313 26945 17325 26948
rect 17359 26976 17371 26979
rect 17678 26976 17684 26988
rect 17359 26948 17684 26976
rect 17359 26945 17371 26948
rect 17313 26939 17371 26945
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 17880 26976 17908 27072
rect 17880 26948 18368 26976
rect 14182 26908 14188 26920
rect 13596 26880 13689 26908
rect 14143 26880 14188 26908
rect 13596 26868 13602 26880
rect 14182 26868 14188 26880
rect 14240 26868 14246 26920
rect 14921 26911 14979 26917
rect 14921 26877 14933 26911
rect 14967 26877 14979 26911
rect 14921 26871 14979 26877
rect 15565 26911 15623 26917
rect 15565 26877 15577 26911
rect 15611 26877 15623 26911
rect 15565 26871 15623 26877
rect 15657 26911 15715 26917
rect 15657 26877 15669 26911
rect 15703 26908 15715 26911
rect 15838 26908 15844 26920
rect 15703 26880 15844 26908
rect 15703 26877 15715 26880
rect 15657 26871 15715 26877
rect 10284 26812 10824 26840
rect 10284 26800 10290 26812
rect 2038 26732 2044 26784
rect 2096 26772 2102 26784
rect 3237 26775 3295 26781
rect 3237 26772 3249 26775
rect 2096 26744 3249 26772
rect 2096 26732 2102 26744
rect 3237 26741 3249 26744
rect 3283 26741 3295 26775
rect 3878 26772 3884 26784
rect 3839 26744 3884 26772
rect 3237 26735 3295 26741
rect 3878 26732 3884 26744
rect 3936 26732 3942 26784
rect 4154 26732 4160 26784
rect 4212 26772 4218 26784
rect 4617 26775 4675 26781
rect 4617 26772 4629 26775
rect 4212 26744 4629 26772
rect 4212 26732 4218 26744
rect 4617 26741 4629 26744
rect 4663 26741 4675 26775
rect 4617 26735 4675 26741
rect 7466 26732 7472 26784
rect 7524 26772 7530 26784
rect 8205 26775 8263 26781
rect 8205 26772 8217 26775
rect 7524 26744 8217 26772
rect 7524 26732 7530 26744
rect 8205 26741 8217 26744
rect 8251 26741 8263 26775
rect 10796 26772 10824 26812
rect 11422 26800 11428 26852
rect 11480 26840 11486 26852
rect 13725 26843 13783 26849
rect 13725 26840 13737 26843
rect 11480 26812 13737 26840
rect 11480 26800 11486 26812
rect 13725 26809 13737 26812
rect 13771 26809 13783 26843
rect 13725 26803 13783 26809
rect 14090 26800 14096 26852
rect 14148 26840 14154 26852
rect 14461 26843 14519 26849
rect 14461 26840 14473 26843
rect 14148 26812 14473 26840
rect 14148 26800 14154 26812
rect 14461 26809 14473 26812
rect 14507 26809 14519 26843
rect 14461 26803 14519 26809
rect 11330 26772 11336 26784
rect 10796 26744 11336 26772
rect 8205 26735 8263 26741
rect 11330 26732 11336 26744
rect 11388 26732 11394 26784
rect 12253 26775 12311 26781
rect 12253 26741 12265 26775
rect 12299 26772 12311 26775
rect 12618 26772 12624 26784
rect 12299 26744 12624 26772
rect 12299 26741 12311 26744
rect 12253 26735 12311 26741
rect 12618 26732 12624 26744
rect 12676 26732 12682 26784
rect 12986 26732 12992 26784
rect 13044 26772 13050 26784
rect 13446 26772 13452 26784
rect 13044 26744 13452 26772
rect 13044 26732 13050 26744
rect 13446 26732 13452 26744
rect 13504 26772 13510 26784
rect 14936 26772 14964 26871
rect 15580 26840 15608 26871
rect 15838 26868 15844 26880
rect 15896 26868 15902 26920
rect 16206 26908 16212 26920
rect 16167 26880 16212 26908
rect 16206 26868 16212 26880
rect 16264 26868 16270 26920
rect 17494 26908 17500 26920
rect 17455 26880 17500 26908
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 17586 26868 17592 26920
rect 17644 26908 17650 26920
rect 17644 26880 17689 26908
rect 17644 26868 17650 26880
rect 17862 26868 17868 26920
rect 17920 26908 17926 26920
rect 18340 26917 18368 26948
rect 21082 26936 21088 26988
rect 21140 26976 21146 26988
rect 21269 26979 21327 26985
rect 21269 26976 21281 26979
rect 21140 26948 21281 26976
rect 21140 26936 21146 26948
rect 21269 26945 21281 26948
rect 21315 26945 21327 26979
rect 21269 26939 21327 26945
rect 18325 26911 18383 26917
rect 17920 26880 17965 26908
rect 17920 26868 17926 26880
rect 18325 26877 18337 26911
rect 18371 26877 18383 26911
rect 18325 26871 18383 26877
rect 18690 26868 18696 26920
rect 18748 26908 18754 26920
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 18748 26880 18981 26908
rect 18748 26868 18754 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 20993 26911 21051 26917
rect 18969 26871 19027 26877
rect 19076 26880 19564 26908
rect 18414 26840 18420 26852
rect 15580 26812 18276 26840
rect 18375 26812 18420 26840
rect 13504 26744 14964 26772
rect 18248 26772 18276 26812
rect 18414 26800 18420 26812
rect 18472 26800 18478 26852
rect 19076 26772 19104 26880
rect 19236 26843 19294 26849
rect 19236 26809 19248 26843
rect 19282 26840 19294 26843
rect 19426 26840 19432 26852
rect 19282 26812 19432 26840
rect 19282 26809 19294 26812
rect 19236 26803 19294 26809
rect 19426 26800 19432 26812
rect 19484 26800 19490 26852
rect 19536 26840 19564 26880
rect 20993 26877 21005 26911
rect 21039 26908 21051 26911
rect 21358 26908 21364 26920
rect 21039 26880 21364 26908
rect 21039 26877 21051 26880
rect 20993 26871 21051 26877
rect 21358 26868 21364 26880
rect 21416 26868 21422 26920
rect 22646 26908 22652 26920
rect 22607 26880 22652 26908
rect 22646 26868 22652 26880
rect 22704 26868 22710 26920
rect 25332 26908 25360 27084
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 26050 27112 26056 27124
rect 26011 27084 26056 27112
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 26418 27072 26424 27124
rect 26476 27112 26482 27124
rect 27154 27112 27160 27124
rect 26476 27084 27160 27112
rect 26476 27072 26482 27084
rect 27154 27072 27160 27084
rect 27212 27072 27218 27124
rect 27706 27072 27712 27124
rect 27764 27112 27770 27124
rect 27801 27115 27859 27121
rect 27801 27112 27813 27115
rect 27764 27084 27813 27112
rect 27764 27072 27770 27084
rect 27801 27081 27813 27084
rect 27847 27081 27859 27115
rect 29362 27112 29368 27124
rect 27801 27075 27859 27081
rect 28184 27084 29368 27112
rect 26602 27044 26608 27056
rect 25516 27016 26608 27044
rect 22848 26880 25360 26908
rect 25409 26911 25467 26917
rect 22848 26840 22876 26880
rect 25409 26877 25421 26911
rect 25455 26908 25467 26911
rect 25516 26908 25544 27016
rect 26602 27004 26608 27016
rect 26660 27004 26666 27056
rect 28184 27053 28212 27084
rect 29362 27072 29368 27084
rect 29420 27112 29426 27124
rect 33042 27112 33048 27124
rect 29420 27084 32904 27112
rect 33003 27084 33048 27112
rect 29420 27072 29426 27084
rect 28169 27047 28227 27053
rect 28169 27044 28181 27047
rect 26712 27016 28181 27044
rect 25590 26936 25596 26988
rect 25648 26976 25654 26988
rect 26510 26976 26516 26988
rect 25648 26948 26372 26976
rect 26471 26948 26516 26976
rect 25648 26936 25654 26948
rect 25455 26880 25544 26908
rect 25455 26877 25467 26880
rect 25409 26871 25467 26877
rect 25774 26868 25780 26920
rect 25832 26908 25838 26920
rect 26344 26917 26372 26948
rect 26510 26936 26516 26948
rect 26568 26976 26574 26988
rect 26712 26976 26740 27016
rect 28169 27013 28181 27016
rect 28215 27013 28227 27047
rect 28169 27007 28227 27013
rect 29181 27047 29239 27053
rect 29181 27013 29193 27047
rect 29227 27044 29239 27047
rect 32214 27044 32220 27056
rect 29227 27016 32220 27044
rect 29227 27013 29239 27016
rect 29181 27007 29239 27013
rect 32214 27004 32220 27016
rect 32272 27004 32278 27056
rect 32876 27044 32904 27084
rect 33042 27072 33048 27084
rect 33100 27072 33106 27124
rect 35526 27112 35532 27124
rect 33152 27084 35532 27112
rect 33152 27044 33180 27084
rect 35526 27072 35532 27084
rect 35584 27072 35590 27124
rect 56778 27112 56784 27124
rect 56739 27084 56784 27112
rect 56778 27072 56784 27084
rect 56836 27072 56842 27124
rect 57241 27115 57299 27121
rect 57241 27081 57253 27115
rect 57287 27112 57299 27115
rect 57698 27112 57704 27124
rect 57287 27084 57704 27112
rect 57287 27081 57299 27084
rect 57241 27075 57299 27081
rect 57698 27072 57704 27084
rect 57756 27072 57762 27124
rect 32876 27016 33180 27044
rect 33410 27004 33416 27056
rect 33468 27044 33474 27056
rect 33468 27016 34836 27044
rect 33468 27004 33474 27016
rect 28261 26979 28319 26985
rect 28261 26976 28273 26979
rect 26568 26948 26740 26976
rect 26804 26948 28273 26976
rect 26568 26936 26574 26948
rect 26804 26920 26832 26948
rect 28261 26945 28273 26948
rect 28307 26945 28319 26979
rect 28261 26939 28319 26945
rect 29273 26979 29331 26985
rect 29273 26945 29285 26979
rect 29319 26976 29331 26979
rect 32122 26976 32128 26988
rect 29319 26948 32128 26976
rect 29319 26945 29331 26948
rect 29273 26939 29331 26945
rect 32122 26936 32128 26948
rect 32180 26936 32186 26988
rect 33778 26976 33784 26988
rect 33428 26948 33784 26976
rect 26237 26911 26295 26917
rect 26237 26908 26249 26911
rect 25832 26880 26249 26908
rect 25832 26868 25838 26880
rect 26237 26877 26249 26880
rect 26283 26877 26295 26911
rect 26237 26871 26295 26877
rect 26329 26911 26387 26917
rect 26329 26877 26341 26911
rect 26375 26877 26387 26911
rect 26329 26871 26387 26877
rect 26605 26911 26663 26917
rect 26605 26877 26617 26911
rect 26651 26908 26663 26911
rect 26786 26908 26792 26920
rect 26651 26880 26792 26908
rect 26651 26877 26663 26880
rect 26605 26871 26663 26877
rect 26786 26868 26792 26880
rect 26844 26868 26850 26920
rect 27982 26908 27988 26920
rect 27943 26880 27988 26908
rect 27982 26868 27988 26880
rect 28040 26868 28046 26920
rect 28994 26868 29000 26920
rect 29052 26908 29058 26920
rect 29089 26911 29147 26917
rect 29089 26908 29101 26911
rect 29052 26880 29101 26908
rect 29052 26868 29058 26880
rect 29089 26877 29101 26880
rect 29135 26877 29147 26911
rect 29089 26871 29147 26877
rect 29365 26911 29423 26917
rect 29365 26877 29377 26911
rect 29411 26877 29423 26911
rect 29365 26871 29423 26877
rect 19536 26812 20484 26840
rect 18248 26744 19104 26772
rect 13504 26732 13510 26744
rect 19334 26732 19340 26784
rect 19392 26772 19398 26784
rect 20349 26775 20407 26781
rect 20349 26772 20361 26775
rect 19392 26744 20361 26772
rect 19392 26732 19398 26744
rect 20349 26741 20361 26744
rect 20395 26741 20407 26775
rect 20456 26772 20484 26812
rect 22204 26812 22876 26840
rect 22916 26843 22974 26849
rect 20714 26772 20720 26784
rect 20456 26744 20720 26772
rect 20349 26735 20407 26741
rect 20714 26732 20720 26744
rect 20772 26772 20778 26784
rect 21269 26775 21327 26781
rect 21269 26772 21281 26775
rect 20772 26744 21281 26772
rect 20772 26732 20778 26744
rect 21269 26741 21281 26744
rect 21315 26741 21327 26775
rect 21269 26735 21327 26741
rect 21358 26732 21364 26784
rect 21416 26772 21422 26784
rect 22204 26772 22232 26812
rect 22916 26809 22928 26843
rect 22962 26840 22974 26843
rect 23014 26840 23020 26852
rect 22962 26812 23020 26840
rect 22962 26809 22974 26812
rect 22916 26803 22974 26809
rect 23014 26800 23020 26812
rect 23072 26800 23078 26852
rect 24578 26840 24584 26852
rect 24539 26812 24584 26840
rect 24578 26800 24584 26812
rect 24636 26800 24642 26852
rect 25222 26840 25228 26852
rect 25183 26812 25228 26840
rect 25222 26800 25228 26812
rect 25280 26800 25286 26852
rect 25593 26843 25651 26849
rect 25593 26809 25605 26843
rect 25639 26840 25651 26843
rect 28000 26840 28028 26868
rect 29380 26840 29408 26871
rect 29454 26868 29460 26920
rect 29512 26908 29518 26920
rect 29549 26911 29607 26917
rect 29549 26908 29561 26911
rect 29512 26880 29561 26908
rect 29512 26868 29518 26880
rect 29549 26877 29561 26880
rect 29595 26877 29607 26911
rect 30006 26908 30012 26920
rect 29967 26880 30012 26908
rect 29549 26871 29607 26877
rect 30006 26868 30012 26880
rect 30064 26868 30070 26920
rect 30190 26908 30196 26920
rect 30151 26880 30196 26908
rect 30190 26868 30196 26880
rect 30248 26868 30254 26920
rect 30374 26908 30380 26920
rect 30335 26880 30380 26908
rect 30374 26868 30380 26880
rect 30432 26868 30438 26920
rect 31386 26908 31392 26920
rect 30484 26880 31392 26908
rect 30208 26840 30236 26868
rect 25639 26812 28028 26840
rect 28092 26812 29040 26840
rect 29380 26812 30236 26840
rect 25639 26809 25651 26812
rect 25593 26803 25651 26809
rect 21416 26744 22232 26772
rect 21416 26732 21422 26744
rect 22278 26732 22284 26784
rect 22336 26772 22342 26784
rect 28092 26772 28120 26812
rect 22336 26744 28120 26772
rect 22336 26732 22342 26744
rect 28534 26732 28540 26784
rect 28592 26772 28598 26784
rect 28905 26775 28963 26781
rect 28905 26772 28917 26775
rect 28592 26744 28917 26772
rect 28592 26732 28598 26744
rect 28905 26741 28917 26744
rect 28951 26741 28963 26775
rect 29012 26772 29040 26812
rect 30282 26800 30288 26852
rect 30340 26840 30346 26852
rect 30340 26812 30385 26840
rect 30340 26800 30346 26812
rect 30484 26772 30512 26880
rect 31386 26868 31392 26880
rect 31444 26868 31450 26920
rect 31665 26911 31723 26917
rect 31665 26877 31677 26911
rect 31711 26908 31723 26911
rect 31938 26908 31944 26920
rect 31711 26880 31944 26908
rect 31711 26877 31723 26880
rect 31665 26871 31723 26877
rect 31938 26868 31944 26880
rect 31996 26868 32002 26920
rect 33318 26908 33324 26920
rect 33279 26880 33324 26908
rect 33318 26868 33324 26880
rect 33376 26868 33382 26920
rect 33428 26917 33456 26948
rect 33778 26936 33784 26948
rect 33836 26936 33842 26988
rect 34698 26936 34704 26988
rect 34756 26976 34762 26988
rect 34808 26985 34836 27016
rect 34793 26979 34851 26985
rect 34793 26976 34805 26979
rect 34756 26948 34805 26976
rect 34756 26936 34762 26948
rect 34793 26945 34805 26948
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 56045 26979 56103 26985
rect 56045 26945 56057 26979
rect 56091 26976 56103 26979
rect 56870 26976 56876 26988
rect 56091 26948 56876 26976
rect 56091 26945 56103 26948
rect 56045 26939 56103 26945
rect 56870 26936 56876 26948
rect 56928 26936 56934 26988
rect 33413 26911 33471 26917
rect 33413 26877 33425 26911
rect 33459 26877 33471 26911
rect 33413 26871 33471 26877
rect 33502 26868 33508 26920
rect 33560 26908 33566 26920
rect 33560 26880 33605 26908
rect 33560 26868 33566 26880
rect 33686 26868 33692 26920
rect 33744 26908 33750 26920
rect 34149 26911 34207 26917
rect 33744 26880 33789 26908
rect 33744 26868 33750 26880
rect 34149 26877 34161 26911
rect 34195 26877 34207 26911
rect 57422 26908 57428 26920
rect 57383 26880 57428 26908
rect 34149 26871 34207 26877
rect 31110 26840 31116 26852
rect 30576 26812 31116 26840
rect 30576 26781 30604 26812
rect 31110 26800 31116 26812
rect 31168 26840 31174 26852
rect 31481 26843 31539 26849
rect 31481 26840 31493 26843
rect 31168 26812 31493 26840
rect 31168 26800 31174 26812
rect 31481 26809 31493 26812
rect 31527 26809 31539 26843
rect 31481 26803 31539 26809
rect 33042 26800 33048 26852
rect 33100 26840 33106 26852
rect 34164 26840 34192 26871
rect 57422 26868 57428 26880
rect 57480 26868 57486 26920
rect 33100 26812 34192 26840
rect 35060 26843 35118 26849
rect 33100 26800 33106 26812
rect 35060 26809 35072 26843
rect 35106 26840 35118 26843
rect 37182 26840 37188 26852
rect 35106 26812 37188 26840
rect 35106 26809 35118 26812
rect 35060 26803 35118 26809
rect 37182 26800 37188 26812
rect 37240 26800 37246 26852
rect 55398 26840 55404 26852
rect 55359 26812 55404 26840
rect 55398 26800 55404 26812
rect 55456 26800 55462 26852
rect 55490 26800 55496 26852
rect 55548 26840 55554 26852
rect 57974 26840 57980 26852
rect 55548 26812 55593 26840
rect 57935 26812 57980 26840
rect 55548 26800 55554 26812
rect 57974 26800 57980 26812
rect 58032 26800 58038 26852
rect 29012 26744 30512 26772
rect 30561 26775 30619 26781
rect 28905 26735 28963 26741
rect 30561 26741 30573 26775
rect 30607 26741 30619 26775
rect 31846 26772 31852 26784
rect 31807 26744 31852 26772
rect 30561 26735 30619 26741
rect 31846 26732 31852 26744
rect 31904 26732 31910 26784
rect 32766 26732 32772 26784
rect 32824 26772 32830 26784
rect 34241 26775 34299 26781
rect 34241 26772 34253 26775
rect 32824 26744 34253 26772
rect 32824 26732 32830 26744
rect 34241 26741 34253 26744
rect 34287 26741 34299 26775
rect 34241 26735 34299 26741
rect 35618 26732 35624 26784
rect 35676 26772 35682 26784
rect 36173 26775 36231 26781
rect 36173 26772 36185 26775
rect 35676 26744 36185 26772
rect 35676 26732 35682 26744
rect 36173 26741 36185 26744
rect 36219 26741 36231 26775
rect 36173 26735 36231 26741
rect 58069 26775 58127 26781
rect 58069 26741 58081 26775
rect 58115 26772 58127 26775
rect 58342 26772 58348 26784
rect 58115 26744 58348 26772
rect 58115 26741 58127 26744
rect 58069 26735 58127 26741
rect 58342 26732 58348 26744
rect 58400 26732 58406 26784
rect 1104 26682 58880 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 50326 26682
rect 50378 26630 50390 26682
rect 50442 26630 50454 26682
rect 50506 26630 50518 26682
rect 50570 26630 58880 26682
rect 1104 26608 58880 26630
rect 2498 26568 2504 26580
rect 2459 26540 2504 26568
rect 2498 26528 2504 26540
rect 2556 26528 2562 26580
rect 4522 26528 4528 26580
rect 4580 26568 4586 26580
rect 7561 26571 7619 26577
rect 7561 26568 7573 26571
rect 4580 26540 7573 26568
rect 4580 26528 4586 26540
rect 7561 26537 7573 26540
rect 7607 26568 7619 26571
rect 7742 26568 7748 26580
rect 7607 26540 7748 26568
rect 7607 26537 7619 26540
rect 7561 26531 7619 26537
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8478 26568 8484 26580
rect 8439 26540 8484 26568
rect 8478 26528 8484 26540
rect 8536 26528 8542 26580
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 10870 26568 10876 26580
rect 9732 26540 10876 26568
rect 9732 26528 9738 26540
rect 10870 26528 10876 26540
rect 10928 26528 10934 26580
rect 11238 26528 11244 26580
rect 11296 26568 11302 26580
rect 12342 26568 12348 26580
rect 11296 26540 12348 26568
rect 11296 26528 11302 26540
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 12434 26528 12440 26580
rect 12492 26568 12498 26580
rect 12618 26568 12624 26580
rect 12492 26540 12624 26568
rect 12492 26528 12498 26540
rect 12618 26528 12624 26540
rect 12676 26528 12682 26580
rect 16117 26571 16175 26577
rect 16117 26537 16129 26571
rect 16163 26568 16175 26571
rect 16206 26568 16212 26580
rect 16163 26540 16212 26568
rect 16163 26537 16175 26540
rect 16117 26531 16175 26537
rect 16206 26528 16212 26540
rect 16264 26568 16270 26580
rect 16264 26540 16896 26568
rect 16264 26528 16270 26540
rect 4617 26503 4675 26509
rect 4617 26500 4629 26503
rect 1872 26472 4629 26500
rect 1872 26441 1900 26472
rect 4617 26469 4629 26472
rect 4663 26469 4675 26503
rect 9490 26500 9496 26512
rect 4617 26463 4675 26469
rect 8404 26472 9496 26500
rect 1857 26435 1915 26441
rect 1857 26401 1869 26435
rect 1903 26401 1915 26435
rect 2038 26432 2044 26444
rect 1999 26404 2044 26432
rect 1857 26395 1915 26401
rect 2038 26392 2044 26404
rect 2096 26392 2102 26444
rect 3050 26432 3056 26444
rect 3011 26404 3056 26432
rect 3050 26392 3056 26404
rect 3108 26392 3114 26444
rect 4525 26435 4583 26441
rect 4525 26401 4537 26435
rect 4571 26401 4583 26435
rect 4706 26432 4712 26444
rect 4667 26404 4712 26432
rect 4525 26395 4583 26401
rect 4540 26364 4568 26395
rect 4706 26392 4712 26404
rect 4764 26392 4770 26444
rect 5350 26432 5356 26444
rect 5311 26404 5356 26432
rect 5350 26392 5356 26404
rect 5408 26392 5414 26444
rect 6178 26432 6184 26444
rect 6139 26404 6184 26432
rect 6178 26392 6184 26404
rect 6236 26392 6242 26444
rect 6825 26435 6883 26441
rect 6825 26401 6837 26435
rect 6871 26432 6883 26435
rect 6914 26432 6920 26444
rect 6871 26404 6920 26432
rect 6871 26401 6883 26404
rect 6825 26395 6883 26401
rect 6914 26392 6920 26404
rect 6972 26392 6978 26444
rect 7006 26392 7012 26444
rect 7064 26432 7070 26444
rect 7466 26432 7472 26444
rect 7064 26404 7109 26432
rect 7427 26404 7472 26432
rect 7064 26392 7070 26404
rect 7466 26392 7472 26404
rect 7524 26392 7530 26444
rect 8404 26441 8432 26472
rect 9490 26460 9496 26472
rect 9548 26460 9554 26512
rect 15010 26509 15016 26512
rect 13817 26503 13875 26509
rect 13817 26500 13829 26503
rect 10060 26472 13829 26500
rect 8389 26435 8447 26441
rect 8389 26401 8401 26435
rect 8435 26401 8447 26435
rect 8389 26395 8447 26401
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26401 8631 26435
rect 8573 26395 8631 26401
rect 9769 26435 9827 26441
rect 9769 26401 9781 26435
rect 9815 26432 9827 26435
rect 9858 26432 9864 26444
rect 9815 26404 9864 26432
rect 9815 26401 9827 26404
rect 9769 26395 9827 26401
rect 4540 26336 8156 26364
rect 6825 26299 6883 26305
rect 6825 26265 6837 26299
rect 6871 26296 6883 26299
rect 7190 26296 7196 26308
rect 6871 26268 7196 26296
rect 6871 26265 6883 26268
rect 6825 26259 6883 26265
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 8128 26296 8156 26336
rect 8202 26324 8208 26376
rect 8260 26364 8266 26376
rect 8588 26364 8616 26395
rect 9858 26392 9864 26404
rect 9916 26392 9922 26444
rect 10060 26441 10088 26472
rect 13817 26469 13829 26472
rect 13863 26469 13875 26503
rect 13817 26463 13875 26469
rect 15004 26463 15016 26509
rect 15068 26500 15074 26512
rect 15068 26472 15104 26500
rect 15010 26460 15016 26463
rect 15068 26460 15074 26472
rect 9953 26435 10011 26441
rect 9953 26401 9965 26435
rect 9999 26401 10011 26435
rect 9953 26395 10011 26401
rect 10045 26435 10103 26441
rect 10045 26401 10057 26435
rect 10091 26401 10103 26435
rect 10318 26432 10324 26444
rect 10279 26404 10324 26432
rect 10045 26395 10103 26401
rect 8260 26336 8616 26364
rect 9968 26364 9996 26395
rect 10318 26392 10324 26404
rect 10376 26392 10382 26444
rect 10410 26392 10416 26444
rect 10468 26432 10474 26444
rect 10778 26432 10784 26444
rect 10468 26404 10784 26432
rect 10468 26392 10474 26404
rect 10778 26392 10784 26404
rect 10836 26432 10842 26444
rect 10965 26435 11023 26441
rect 10965 26432 10977 26435
rect 10836 26404 10977 26432
rect 10836 26392 10842 26404
rect 10965 26401 10977 26404
rect 11011 26401 11023 26435
rect 11146 26432 11152 26444
rect 11107 26404 11152 26432
rect 10965 26395 11023 26401
rect 11146 26392 11152 26404
rect 11204 26392 11210 26444
rect 11250 26435 11308 26441
rect 11250 26401 11262 26435
rect 11296 26432 11308 26435
rect 11422 26432 11428 26444
rect 11296 26404 11428 26432
rect 11296 26401 11308 26404
rect 11250 26395 11308 26401
rect 11422 26392 11428 26404
rect 11480 26392 11486 26444
rect 11514 26392 11520 26444
rect 11572 26432 11578 26444
rect 11572 26404 11617 26432
rect 11572 26392 11578 26404
rect 11974 26392 11980 26444
rect 12032 26432 12038 26444
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 12032 26404 12173 26432
rect 12032 26392 12038 26404
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 12342 26432 12348 26444
rect 12303 26404 12348 26432
rect 12161 26395 12219 26401
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 12434 26392 12440 26444
rect 12492 26432 12498 26444
rect 12710 26432 12716 26444
rect 12492 26404 12537 26432
rect 12671 26404 12716 26432
rect 12492 26392 12498 26404
rect 12710 26392 12716 26404
rect 12768 26392 12774 26444
rect 13541 26435 13599 26441
rect 13541 26401 13553 26435
rect 13587 26432 13599 26435
rect 15470 26432 15476 26444
rect 13587 26404 15476 26432
rect 13587 26401 13599 26404
rect 13541 26395 13599 26401
rect 15470 26392 15476 26404
rect 15528 26392 15534 26444
rect 16868 26441 16896 26540
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 21358 26568 21364 26580
rect 17000 26540 21364 26568
rect 17000 26528 17006 26540
rect 21358 26528 21364 26540
rect 21416 26528 21422 26580
rect 21818 26568 21824 26580
rect 21468 26540 21824 26568
rect 17034 26460 17040 26512
rect 17092 26500 17098 26512
rect 21468 26500 21496 26540
rect 21818 26528 21824 26540
rect 21876 26528 21882 26580
rect 23382 26528 23388 26580
rect 23440 26528 23446 26580
rect 25590 26528 25596 26580
rect 25648 26568 25654 26580
rect 25685 26571 25743 26577
rect 25685 26568 25697 26571
rect 25648 26540 25697 26568
rect 25648 26528 25654 26540
rect 25685 26537 25697 26540
rect 25731 26568 25743 26571
rect 27157 26571 27215 26577
rect 27157 26568 27169 26571
rect 25731 26540 27169 26568
rect 25731 26537 25743 26540
rect 25685 26531 25743 26537
rect 27157 26537 27169 26540
rect 27203 26537 27215 26571
rect 27157 26531 27215 26537
rect 29549 26571 29607 26577
rect 29549 26537 29561 26571
rect 29595 26568 29607 26571
rect 30282 26568 30288 26580
rect 29595 26540 30288 26568
rect 29595 26537 29607 26540
rect 29549 26531 29607 26537
rect 30282 26528 30288 26540
rect 30340 26528 30346 26580
rect 31297 26571 31355 26577
rect 31297 26537 31309 26571
rect 31343 26568 31355 26571
rect 31938 26568 31944 26580
rect 31343 26540 31944 26568
rect 31343 26537 31355 26540
rect 31297 26531 31355 26537
rect 31938 26528 31944 26540
rect 31996 26528 32002 26580
rect 32122 26568 32128 26580
rect 32083 26540 32128 26568
rect 32122 26528 32128 26540
rect 32180 26528 32186 26580
rect 33229 26571 33287 26577
rect 33229 26537 33241 26571
rect 33275 26568 33287 26571
rect 33686 26568 33692 26580
rect 33275 26540 33692 26568
rect 33275 26537 33287 26540
rect 33229 26531 33287 26537
rect 33686 26528 33692 26540
rect 33744 26528 33750 26580
rect 37182 26568 37188 26580
rect 37143 26540 37188 26568
rect 37182 26528 37188 26540
rect 37240 26528 37246 26580
rect 55769 26571 55827 26577
rect 41386 26540 45554 26568
rect 23400 26500 23428 26528
rect 17092 26472 21496 26500
rect 21744 26472 23428 26500
rect 23477 26503 23535 26509
rect 17092 26460 17098 26472
rect 16761 26435 16819 26441
rect 16761 26401 16773 26435
rect 16807 26401 16819 26435
rect 16761 26395 16819 26401
rect 16853 26435 16911 26441
rect 16853 26401 16865 26435
rect 16899 26401 16911 26435
rect 16853 26395 16911 26401
rect 10137 26367 10195 26373
rect 9968 26336 10088 26364
rect 8260 26324 8266 26336
rect 10060 26296 10088 26336
rect 10137 26333 10149 26367
rect 10183 26364 10195 26367
rect 10226 26364 10232 26376
rect 10183 26336 10232 26364
rect 10183 26333 10195 26336
rect 10137 26327 10195 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 11164 26296 11192 26392
rect 11330 26364 11336 26376
rect 11243 26336 11336 26364
rect 11330 26324 11336 26336
rect 11388 26364 11394 26376
rect 12529 26367 12587 26373
rect 12529 26364 12541 26367
rect 11388 26336 12541 26364
rect 11388 26324 11394 26336
rect 12529 26333 12541 26336
rect 12575 26333 12587 26367
rect 12529 26327 12587 26333
rect 13170 26324 13176 26376
rect 13228 26364 13234 26376
rect 13446 26364 13452 26376
rect 13228 26336 13452 26364
rect 13228 26324 13234 26336
rect 13446 26324 13452 26336
rect 13504 26324 13510 26376
rect 13814 26364 13820 26376
rect 13775 26336 13820 26364
rect 13814 26324 13820 26336
rect 13872 26324 13878 26376
rect 14366 26324 14372 26376
rect 14424 26364 14430 26376
rect 14737 26367 14795 26373
rect 14737 26364 14749 26367
rect 14424 26336 14749 26364
rect 14424 26324 14430 26336
rect 14737 26333 14749 26336
rect 14783 26333 14795 26367
rect 14737 26327 14795 26333
rect 16206 26324 16212 26376
rect 16264 26364 16270 26376
rect 16776 26364 16804 26395
rect 16942 26392 16948 26444
rect 17000 26432 17006 26444
rect 17129 26435 17187 26441
rect 17129 26432 17141 26435
rect 17000 26404 17141 26432
rect 17000 26392 17006 26404
rect 17129 26401 17141 26404
rect 17175 26432 17187 26435
rect 17494 26432 17500 26444
rect 17175 26404 17500 26432
rect 17175 26401 17187 26404
rect 17129 26395 17187 26401
rect 17494 26392 17500 26404
rect 17552 26392 17558 26444
rect 17586 26392 17592 26444
rect 17644 26432 17650 26444
rect 17681 26435 17739 26441
rect 17681 26432 17693 26435
rect 17644 26404 17693 26432
rect 17644 26392 17650 26404
rect 17681 26401 17693 26404
rect 17727 26401 17739 26435
rect 19334 26432 19340 26444
rect 17681 26395 17739 26401
rect 17788 26404 19340 26432
rect 17788 26364 17816 26404
rect 19334 26392 19340 26404
rect 19392 26392 19398 26444
rect 19886 26392 19892 26444
rect 19944 26432 19950 26444
rect 20806 26432 20812 26444
rect 19944 26404 20291 26432
rect 20767 26404 20812 26432
rect 19944 26392 19950 26404
rect 16264 26336 17816 26364
rect 16264 26324 16270 26336
rect 17862 26324 17868 26376
rect 17920 26364 17926 26376
rect 18322 26364 18328 26376
rect 17920 26336 17965 26364
rect 18283 26336 18328 26364
rect 17920 26324 17926 26336
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 19058 26324 19064 26376
rect 19116 26364 19122 26376
rect 20165 26367 20223 26373
rect 20165 26364 20177 26367
rect 19116 26336 20177 26364
rect 19116 26324 19122 26336
rect 20165 26333 20177 26336
rect 20211 26333 20223 26367
rect 20263 26364 20291 26404
rect 20806 26392 20812 26404
rect 20864 26392 20870 26444
rect 21082 26392 21088 26444
rect 21140 26432 21146 26444
rect 21450 26432 21456 26444
rect 21140 26404 21456 26432
rect 21140 26392 21146 26404
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 21646 26435 21704 26441
rect 21646 26401 21658 26435
rect 21692 26432 21704 26435
rect 21744 26432 21772 26472
rect 23477 26469 23489 26503
rect 23523 26500 23535 26503
rect 23658 26500 23664 26512
rect 23523 26472 23664 26500
rect 23523 26469 23535 26472
rect 23477 26463 23535 26469
rect 23658 26460 23664 26472
rect 23716 26460 23722 26512
rect 21692 26404 21772 26432
rect 21692 26401 21704 26404
rect 21646 26395 21704 26401
rect 21818 26392 21824 26444
rect 21876 26432 21882 26444
rect 21913 26435 21971 26441
rect 21913 26432 21925 26435
rect 21876 26404 21925 26432
rect 21876 26392 21882 26404
rect 21913 26401 21925 26404
rect 21959 26401 21971 26435
rect 21913 26395 21971 26401
rect 22186 26392 22192 26444
rect 22244 26432 22250 26444
rect 22465 26435 22523 26441
rect 22465 26432 22477 26435
rect 22244 26404 22477 26432
rect 22244 26392 22250 26404
rect 22465 26401 22477 26404
rect 22511 26401 22523 26435
rect 22465 26395 22523 26401
rect 23293 26435 23351 26441
rect 23293 26401 23305 26435
rect 23339 26432 23351 26435
rect 23382 26432 23388 26444
rect 23339 26404 23388 26432
rect 23339 26401 23351 26404
rect 23293 26395 23351 26401
rect 23382 26392 23388 26404
rect 23440 26432 23446 26444
rect 23937 26435 23995 26441
rect 23937 26432 23949 26435
rect 23440 26404 23949 26432
rect 23440 26392 23446 26404
rect 23937 26401 23949 26404
rect 23983 26401 23995 26435
rect 23937 26395 23995 26401
rect 25409 26435 25467 26441
rect 25409 26401 25421 26435
rect 25455 26432 25467 26435
rect 25608 26432 25636 26528
rect 25958 26460 25964 26512
rect 26016 26500 26022 26512
rect 30558 26500 30564 26512
rect 26016 26472 30564 26500
rect 26016 26460 26022 26472
rect 30558 26460 30564 26472
rect 30616 26460 30622 26512
rect 31110 26500 31116 26512
rect 31071 26472 31116 26500
rect 31110 26460 31116 26472
rect 31168 26500 31174 26512
rect 32950 26500 32956 26512
rect 31168 26472 31800 26500
rect 32911 26472 32956 26500
rect 31168 26460 31174 26472
rect 26602 26432 26608 26444
rect 25455 26404 25636 26432
rect 26563 26404 26608 26432
rect 25455 26401 25467 26404
rect 25409 26395 25467 26401
rect 26602 26392 26608 26404
rect 26660 26392 26666 26444
rect 26786 26432 26792 26444
rect 26699 26404 26792 26432
rect 26786 26392 26792 26404
rect 26844 26392 26850 26444
rect 26878 26392 26884 26444
rect 26936 26432 26942 26444
rect 27019 26435 27077 26441
rect 26936 26404 26981 26432
rect 26936 26392 26942 26404
rect 27019 26401 27031 26435
rect 27065 26432 27077 26435
rect 28258 26432 28264 26444
rect 27065 26404 28264 26432
rect 27065 26401 27077 26404
rect 27019 26395 27077 26401
rect 28258 26392 28264 26404
rect 28316 26392 28322 26444
rect 28436 26435 28494 26441
rect 28436 26401 28448 26435
rect 28482 26432 28494 26435
rect 29546 26432 29552 26444
rect 28482 26404 29552 26432
rect 28482 26401 28494 26404
rect 28436 26395 28494 26401
rect 29546 26392 29552 26404
rect 29604 26392 29610 26444
rect 31772 26441 31800 26472
rect 32950 26460 32956 26472
rect 33008 26500 33014 26512
rect 33008 26472 33732 26500
rect 33008 26460 33014 26472
rect 30929 26435 30987 26441
rect 30929 26401 30941 26435
rect 30975 26401 30987 26435
rect 30929 26395 30987 26401
rect 31757 26435 31815 26441
rect 31757 26401 31769 26435
rect 31803 26401 31815 26435
rect 31757 26395 31815 26401
rect 31941 26435 31999 26441
rect 31941 26401 31953 26435
rect 31987 26432 31999 26435
rect 32306 26432 32312 26444
rect 31987 26404 32312 26432
rect 31987 26401 31999 26404
rect 31941 26395 31999 26401
rect 21545 26367 21603 26373
rect 21545 26364 21557 26367
rect 20263 26336 21557 26364
rect 20165 26327 20223 26333
rect 21545 26333 21557 26336
rect 21591 26333 21603 26367
rect 21545 26327 21603 26333
rect 21729 26367 21787 26373
rect 21729 26333 21741 26367
rect 21775 26364 21787 26367
rect 22002 26364 22008 26376
rect 21775 26336 22008 26364
rect 21775 26333 21787 26336
rect 21729 26327 21787 26333
rect 22002 26324 22008 26336
rect 22060 26324 22066 26376
rect 25225 26367 25283 26373
rect 25225 26333 25237 26367
rect 25271 26364 25283 26367
rect 25774 26364 25780 26376
rect 25271 26336 25780 26364
rect 25271 26333 25283 26336
rect 25225 26327 25283 26333
rect 25774 26324 25780 26336
rect 25832 26324 25838 26376
rect 26804 26364 26832 26392
rect 27154 26364 27160 26376
rect 26804 26336 27160 26364
rect 27154 26324 27160 26336
rect 27212 26324 27218 26376
rect 27246 26324 27252 26376
rect 27304 26364 27310 26376
rect 28169 26367 28227 26373
rect 28169 26364 28181 26367
rect 27304 26336 28181 26364
rect 27304 26324 27310 26336
rect 28169 26333 28181 26336
rect 28215 26333 28227 26367
rect 30944 26364 30972 26395
rect 31956 26364 31984 26395
rect 32306 26392 32312 26404
rect 32364 26392 32370 26444
rect 32582 26432 32588 26444
rect 32543 26404 32588 26432
rect 32582 26392 32588 26404
rect 32640 26392 32646 26444
rect 32766 26441 32772 26444
rect 32733 26435 32772 26441
rect 32733 26401 32745 26435
rect 32733 26395 32772 26401
rect 32766 26392 32772 26395
rect 32824 26392 32830 26444
rect 32858 26392 32864 26444
rect 32916 26432 32922 26444
rect 32916 26404 32961 26432
rect 32916 26392 32922 26404
rect 33042 26392 33048 26444
rect 33100 26441 33106 26444
rect 33704 26441 33732 26472
rect 33778 26460 33784 26512
rect 33836 26500 33842 26512
rect 34790 26500 34796 26512
rect 33836 26472 34796 26500
rect 33836 26460 33842 26472
rect 33891 26441 33919 26472
rect 34790 26460 34796 26472
rect 34848 26460 34854 26512
rect 35802 26460 35808 26512
rect 35860 26500 35866 26512
rect 35860 26472 36492 26500
rect 35860 26460 35866 26472
rect 33100 26432 33108 26441
rect 33689 26435 33747 26441
rect 33100 26404 33145 26432
rect 33100 26395 33108 26404
rect 33689 26401 33701 26435
rect 33735 26401 33747 26435
rect 33689 26395 33747 26401
rect 33874 26435 33932 26441
rect 33874 26401 33886 26435
rect 33920 26401 33932 26435
rect 33874 26395 33932 26401
rect 33100 26392 33106 26395
rect 33962 26392 33968 26444
rect 34020 26432 34026 26444
rect 34241 26435 34299 26441
rect 34020 26404 34065 26432
rect 34020 26392 34026 26404
rect 34241 26401 34253 26435
rect 34287 26401 34299 26435
rect 36354 26432 36360 26444
rect 36315 26404 36360 26432
rect 34241 26395 34299 26401
rect 30944 26336 31984 26364
rect 28169 26327 28227 26333
rect 32398 26324 32404 26376
rect 32456 26364 32462 26376
rect 32876 26364 32904 26392
rect 32456 26336 32904 26364
rect 34256 26364 34284 26395
rect 36354 26392 36360 26404
rect 36412 26392 36418 26444
rect 36464 26441 36492 26472
rect 36630 26460 36636 26512
rect 36688 26500 36694 26512
rect 41386 26500 41414 26540
rect 36688 26472 41414 26500
rect 36688 26460 36694 26472
rect 36449 26435 36507 26441
rect 36449 26401 36461 26435
rect 36495 26401 36507 26435
rect 37090 26432 37096 26444
rect 37051 26404 37096 26432
rect 36449 26395 36507 26401
rect 37090 26392 37096 26404
rect 37148 26392 37154 26444
rect 37277 26435 37335 26441
rect 37277 26401 37289 26435
rect 37323 26401 37335 26435
rect 45526 26432 45554 26540
rect 55769 26537 55781 26571
rect 55815 26568 55827 26571
rect 56686 26568 56692 26580
rect 55815 26540 56692 26568
rect 55815 26537 55827 26540
rect 55769 26531 55827 26537
rect 56686 26528 56692 26540
rect 56744 26528 56750 26580
rect 57974 26528 57980 26580
rect 58032 26568 58038 26580
rect 58161 26571 58219 26577
rect 58161 26568 58173 26571
rect 58032 26540 58173 26568
rect 58032 26528 58038 26540
rect 58161 26537 58173 26540
rect 58207 26537 58219 26571
rect 58161 26531 58219 26537
rect 55125 26435 55183 26441
rect 55125 26432 55137 26435
rect 45526 26404 55137 26432
rect 37277 26395 37335 26401
rect 55125 26401 55137 26404
rect 55171 26401 55183 26435
rect 55125 26395 55183 26401
rect 35250 26364 35256 26376
rect 34256 26336 35256 26364
rect 32456 26324 32462 26336
rect 35250 26324 35256 26336
rect 35308 26364 35314 26376
rect 37292 26364 37320 26395
rect 35308 26336 37320 26364
rect 55309 26367 55367 26373
rect 35308 26324 35314 26336
rect 55309 26333 55321 26367
rect 55355 26364 55367 26367
rect 55950 26364 55956 26376
rect 55355 26336 55956 26364
rect 55355 26333 55367 26336
rect 55309 26327 55367 26333
rect 55950 26324 55956 26336
rect 56008 26324 56014 26376
rect 57057 26367 57115 26373
rect 57057 26333 57069 26367
rect 57103 26364 57115 26367
rect 57517 26367 57575 26373
rect 57517 26364 57529 26367
rect 57103 26336 57529 26364
rect 57103 26333 57115 26336
rect 57057 26327 57115 26333
rect 57517 26333 57529 26336
rect 57563 26333 57575 26367
rect 57517 26327 57575 26333
rect 57701 26367 57759 26373
rect 57701 26333 57713 26367
rect 57747 26364 57759 26367
rect 57974 26364 57980 26376
rect 57747 26336 57980 26364
rect 57747 26333 57759 26336
rect 57701 26327 57759 26333
rect 57974 26324 57980 26336
rect 58032 26324 58038 26376
rect 8128 26268 9904 26296
rect 10060 26268 11192 26296
rect 3142 26228 3148 26240
rect 3103 26200 3148 26228
rect 3142 26188 3148 26200
rect 3200 26188 3206 26240
rect 6270 26228 6276 26240
rect 6231 26200 6276 26228
rect 6270 26188 6276 26200
rect 6328 26188 6334 26240
rect 6730 26188 6736 26240
rect 6788 26228 6794 26240
rect 9674 26228 9680 26240
rect 6788 26200 9680 26228
rect 6788 26188 6794 26200
rect 9674 26188 9680 26200
rect 9732 26188 9738 26240
rect 9876 26228 9904 26268
rect 13538 26256 13544 26308
rect 13596 26296 13602 26308
rect 13633 26299 13691 26305
rect 13633 26296 13645 26299
rect 13596 26268 13645 26296
rect 13596 26256 13602 26268
rect 13633 26265 13645 26268
rect 13679 26265 13691 26299
rect 13633 26259 13691 26265
rect 16577 26299 16635 26305
rect 16577 26265 16589 26299
rect 16623 26296 16635 26299
rect 17310 26296 17316 26308
rect 16623 26268 17316 26296
rect 16623 26265 16635 26268
rect 16577 26259 16635 26265
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 18969 26299 19027 26305
rect 17420 26268 18920 26296
rect 10042 26228 10048 26240
rect 9876 26200 10048 26228
rect 10042 26188 10048 26200
rect 10100 26188 10106 26240
rect 10502 26228 10508 26240
rect 10463 26200 10508 26228
rect 10502 26188 10508 26200
rect 10560 26188 10566 26240
rect 11698 26228 11704 26240
rect 11659 26200 11704 26228
rect 11698 26188 11704 26200
rect 11756 26188 11762 26240
rect 12894 26228 12900 26240
rect 12855 26200 12900 26228
rect 12894 26188 12900 26200
rect 12952 26188 12958 26240
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 17037 26231 17095 26237
rect 17037 26228 17049 26231
rect 15528 26200 17049 26228
rect 15528 26188 15534 26200
rect 17037 26197 17049 26200
rect 17083 26197 17095 26231
rect 17037 26191 17095 26197
rect 17126 26188 17132 26240
rect 17184 26228 17190 26240
rect 17420 26228 17448 26268
rect 17184 26200 17448 26228
rect 18892 26228 18920 26268
rect 18969 26265 18981 26299
rect 19015 26296 19027 26299
rect 19015 26268 21496 26296
rect 19015 26265 19027 26268
rect 18969 26259 19027 26265
rect 21082 26228 21088 26240
rect 18892 26200 21088 26228
rect 17184 26188 17190 26200
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 21266 26228 21272 26240
rect 21227 26200 21272 26228
rect 21266 26188 21272 26200
rect 21324 26188 21330 26240
rect 21468 26228 21496 26268
rect 21818 26256 21824 26308
rect 21876 26296 21882 26308
rect 22649 26299 22707 26305
rect 22649 26296 22661 26299
rect 21876 26268 22661 26296
rect 21876 26256 21882 26268
rect 22649 26265 22661 26268
rect 22695 26265 22707 26299
rect 22649 26259 22707 26265
rect 25332 26268 25636 26296
rect 21634 26228 21640 26240
rect 21468 26200 21640 26228
rect 21634 26188 21640 26200
rect 21692 26188 21698 26240
rect 23658 26188 23664 26240
rect 23716 26228 23722 26240
rect 24121 26231 24179 26237
rect 24121 26228 24133 26231
rect 23716 26200 24133 26228
rect 23716 26188 23722 26200
rect 24121 26197 24133 26200
rect 24167 26228 24179 26231
rect 25332 26228 25360 26268
rect 25498 26228 25504 26240
rect 24167 26200 25360 26228
rect 25459 26200 25504 26228
rect 24167 26197 24179 26200
rect 24121 26191 24179 26197
rect 25498 26188 25504 26200
rect 25556 26188 25562 26240
rect 25608 26228 25636 26268
rect 25866 26256 25872 26308
rect 25924 26296 25930 26308
rect 27798 26296 27804 26308
rect 25924 26268 27804 26296
rect 25924 26256 25930 26268
rect 27798 26256 27804 26268
rect 27856 26256 27862 26308
rect 34149 26299 34207 26305
rect 34149 26265 34161 26299
rect 34195 26296 34207 26299
rect 34514 26296 34520 26308
rect 34195 26268 34520 26296
rect 34195 26265 34207 26268
rect 34149 26259 34207 26265
rect 34514 26256 34520 26268
rect 34572 26256 34578 26308
rect 36541 26299 36599 26305
rect 36541 26265 36553 26299
rect 36587 26296 36599 26299
rect 55398 26296 55404 26308
rect 36587 26268 55404 26296
rect 36587 26265 36599 26268
rect 36541 26259 36599 26265
rect 55398 26256 55404 26268
rect 55456 26256 55462 26308
rect 29178 26228 29184 26240
rect 25608 26200 29184 26228
rect 29178 26188 29184 26200
rect 29236 26188 29242 26240
rect 1104 26138 58880 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 58880 26138
rect 1104 26064 58880 26086
rect 2593 26027 2651 26033
rect 2593 25993 2605 26027
rect 2639 26024 2651 26027
rect 3050 26024 3056 26036
rect 2639 25996 3056 26024
rect 2639 25993 2651 25996
rect 2593 25987 2651 25993
rect 3050 25984 3056 25996
rect 3108 25984 3114 26036
rect 5905 26027 5963 26033
rect 4540 25996 5856 26024
rect 4062 25956 4068 25968
rect 1964 25928 4068 25956
rect 1964 25897 1992 25928
rect 4062 25916 4068 25928
rect 4120 25916 4126 25968
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25857 2007 25891
rect 1949 25851 2007 25857
rect 2133 25891 2191 25897
rect 2133 25857 2145 25891
rect 2179 25888 2191 25891
rect 3878 25888 3884 25900
rect 2179 25860 3884 25888
rect 2179 25857 2191 25860
rect 2133 25851 2191 25857
rect 3878 25848 3884 25860
rect 3936 25848 3942 25900
rect 3602 25820 3608 25832
rect 3563 25792 3608 25820
rect 3602 25780 3608 25792
rect 3660 25780 3666 25832
rect 3697 25823 3755 25829
rect 3697 25789 3709 25823
rect 3743 25789 3755 25823
rect 3697 25783 3755 25789
rect 3712 25752 3740 25783
rect 3970 25780 3976 25832
rect 4028 25820 4034 25832
rect 4540 25829 4568 25996
rect 5828 25888 5856 25996
rect 5905 25993 5917 26027
rect 5951 26024 5963 26027
rect 6178 26024 6184 26036
rect 5951 25996 6184 26024
rect 5951 25993 5963 25996
rect 5905 25987 5963 25993
rect 6178 25984 6184 25996
rect 6236 25984 6242 26036
rect 7558 25984 7564 26036
rect 7616 26024 7622 26036
rect 25222 26024 25228 26036
rect 7616 25996 25228 26024
rect 7616 25984 7622 25996
rect 25222 25984 25228 25996
rect 25280 25984 25286 26036
rect 25774 25984 25780 26036
rect 25832 26024 25838 26036
rect 29362 26024 29368 26036
rect 25832 25996 26464 26024
rect 29323 25996 29368 26024
rect 25832 25984 25838 25996
rect 8297 25959 8355 25965
rect 8297 25925 8309 25959
rect 8343 25956 8355 25959
rect 8478 25956 8484 25968
rect 8343 25928 8484 25956
rect 8343 25925 8355 25928
rect 8297 25919 8355 25925
rect 8478 25916 8484 25928
rect 8536 25916 8542 25968
rect 10042 25916 10048 25968
rect 10100 25956 10106 25968
rect 10689 25959 10747 25965
rect 10689 25956 10701 25959
rect 10100 25928 10701 25956
rect 10100 25916 10106 25928
rect 10689 25925 10701 25928
rect 10735 25925 10747 25959
rect 10689 25919 10747 25925
rect 15657 25959 15715 25965
rect 15657 25925 15669 25959
rect 15703 25956 15715 25959
rect 19058 25956 19064 25968
rect 15703 25928 19064 25956
rect 15703 25925 15715 25928
rect 15657 25919 15715 25925
rect 19058 25916 19064 25928
rect 19116 25916 19122 25968
rect 19426 25916 19432 25968
rect 19484 25956 19490 25968
rect 19613 25959 19671 25965
rect 19613 25956 19625 25959
rect 19484 25928 19625 25956
rect 19484 25916 19490 25928
rect 19613 25925 19625 25928
rect 19659 25925 19671 25959
rect 19613 25919 19671 25925
rect 21358 25916 21364 25968
rect 21416 25956 21422 25968
rect 23201 25959 23259 25965
rect 23201 25956 23213 25959
rect 21416 25928 23213 25956
rect 21416 25916 21422 25928
rect 23201 25925 23213 25928
rect 23247 25925 23259 25959
rect 23201 25919 23259 25925
rect 25501 25959 25559 25965
rect 25501 25925 25513 25959
rect 25547 25956 25559 25959
rect 26142 25956 26148 25968
rect 25547 25928 26148 25956
rect 25547 25925 25559 25928
rect 25501 25919 25559 25925
rect 26142 25916 26148 25928
rect 26200 25956 26206 25968
rect 26436 25956 26464 25996
rect 29362 25984 29368 25996
rect 29420 25984 29426 26036
rect 30101 26027 30159 26033
rect 30101 25993 30113 26027
rect 30147 26024 30159 26027
rect 30190 26024 30196 26036
rect 30147 25996 30196 26024
rect 30147 25993 30159 25996
rect 30101 25987 30159 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 31941 26027 31999 26033
rect 31941 25993 31953 26027
rect 31987 26024 31999 26027
rect 32582 26024 32588 26036
rect 31987 25996 32588 26024
rect 31987 25993 31999 25996
rect 31941 25987 31999 25993
rect 32582 25984 32588 25996
rect 32640 25984 32646 26036
rect 33042 26024 33048 26036
rect 33003 25996 33048 26024
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 34885 26027 34943 26033
rect 34885 25993 34897 26027
rect 34931 26024 34943 26027
rect 35250 26024 35256 26036
rect 34931 25996 35256 26024
rect 34931 25993 34943 25996
rect 34885 25987 34943 25993
rect 35250 25984 35256 25996
rect 35308 25984 35314 26036
rect 55309 26027 55367 26033
rect 55309 25993 55321 26027
rect 55355 26024 55367 26027
rect 55490 26024 55496 26036
rect 55355 25996 55496 26024
rect 55355 25993 55367 25996
rect 55309 25987 55367 25993
rect 55490 25984 55496 25996
rect 55548 25984 55554 26036
rect 55950 26024 55956 26036
rect 55911 25996 55956 26024
rect 55950 25984 55956 25996
rect 56008 25984 56014 26036
rect 30745 25959 30803 25965
rect 30745 25956 30757 25959
rect 26200 25928 26372 25956
rect 26436 25928 30757 25956
rect 26200 25916 26206 25928
rect 6917 25891 6975 25897
rect 6917 25888 6929 25891
rect 5828 25860 6929 25888
rect 6917 25857 6929 25860
rect 6963 25857 6975 25891
rect 6917 25851 6975 25857
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25888 15071 25891
rect 18322 25888 18328 25900
rect 15059 25860 18328 25888
rect 15059 25857 15071 25860
rect 15013 25851 15071 25857
rect 4525 25823 4583 25829
rect 4525 25820 4537 25823
rect 4028 25792 4537 25820
rect 4028 25780 4034 25792
rect 4525 25789 4537 25792
rect 4571 25789 4583 25823
rect 6730 25820 6736 25832
rect 4525 25783 4583 25789
rect 4724 25792 6736 25820
rect 4724 25752 4752 25792
rect 6730 25780 6736 25792
rect 6788 25780 6794 25832
rect 6932 25820 6960 25851
rect 18322 25848 18328 25860
rect 18380 25848 18386 25900
rect 19242 25888 19248 25900
rect 19203 25860 19248 25888
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 26344 25897 26372 25928
rect 30745 25925 30757 25928
rect 30791 25925 30803 25959
rect 30745 25919 30803 25925
rect 31110 25916 31116 25968
rect 31168 25956 31174 25968
rect 31168 25928 31213 25956
rect 31168 25916 31174 25928
rect 33318 25916 33324 25968
rect 33376 25956 33382 25968
rect 33505 25959 33563 25965
rect 33505 25956 33517 25959
rect 33376 25928 33517 25956
rect 33376 25916 33382 25928
rect 33505 25925 33517 25928
rect 33551 25925 33563 25959
rect 33505 25919 33563 25925
rect 33962 25916 33968 25968
rect 34020 25956 34026 25968
rect 34149 25959 34207 25965
rect 34149 25956 34161 25959
rect 34020 25928 34161 25956
rect 34020 25916 34026 25928
rect 34149 25925 34161 25928
rect 34195 25956 34207 25959
rect 34238 25956 34244 25968
rect 34195 25928 34244 25956
rect 34195 25925 34207 25928
rect 34149 25919 34207 25925
rect 34238 25916 34244 25928
rect 34296 25956 34302 25968
rect 35618 25956 35624 25968
rect 34296 25928 35624 25956
rect 34296 25916 34302 25928
rect 35618 25916 35624 25928
rect 35676 25916 35682 25968
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25888 20591 25891
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 20579 25860 22569 25888
rect 20579 25857 20591 25860
rect 20533 25851 20591 25857
rect 22557 25857 22569 25860
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 32122 25888 32128 25900
rect 26329 25851 26387 25857
rect 31036 25860 32128 25888
rect 7926 25820 7932 25832
rect 6932 25792 7932 25820
rect 7926 25780 7932 25792
rect 7984 25780 7990 25832
rect 8662 25780 8668 25832
rect 8720 25820 8726 25832
rect 8757 25823 8815 25829
rect 8757 25820 8769 25823
rect 8720 25792 8769 25820
rect 8720 25780 8726 25792
rect 8757 25789 8769 25792
rect 8803 25789 8815 25823
rect 8757 25783 8815 25789
rect 9024 25823 9082 25829
rect 9024 25789 9036 25823
rect 9070 25820 9082 25823
rect 10502 25820 10508 25832
rect 9070 25792 10508 25820
rect 9070 25789 9082 25792
rect 9024 25783 9082 25789
rect 10502 25780 10508 25792
rect 10560 25780 10566 25832
rect 10594 25780 10600 25832
rect 10652 25820 10658 25832
rect 10652 25792 10697 25820
rect 10652 25780 10658 25792
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 11112 25792 12081 25820
rect 11112 25780 11118 25792
rect 12069 25789 12081 25792
rect 12115 25789 12127 25823
rect 12069 25783 12127 25789
rect 12336 25823 12394 25829
rect 12336 25789 12348 25823
rect 12382 25820 12394 25823
rect 12894 25820 12900 25832
rect 12382 25792 12900 25820
rect 12382 25789 12394 25792
rect 12336 25783 12394 25789
rect 12894 25780 12900 25792
rect 12952 25780 12958 25832
rect 14921 25823 14979 25829
rect 14921 25789 14933 25823
rect 14967 25789 14979 25823
rect 15102 25820 15108 25832
rect 15063 25792 15108 25820
rect 14921 25783 14979 25789
rect 3712 25724 4752 25752
rect 4792 25755 4850 25761
rect 4792 25721 4804 25755
rect 4838 25752 4850 25755
rect 5166 25752 5172 25764
rect 4838 25724 5172 25752
rect 4838 25721 4850 25724
rect 4792 25715 4850 25721
rect 5166 25712 5172 25724
rect 5224 25712 5230 25764
rect 7190 25761 7196 25764
rect 7184 25715 7196 25761
rect 7248 25752 7254 25764
rect 7248 25724 7284 25752
rect 7190 25712 7196 25715
rect 7248 25712 7254 25724
rect 7650 25712 7656 25764
rect 7708 25752 7714 25764
rect 10318 25752 10324 25764
rect 7708 25724 10324 25752
rect 7708 25712 7714 25724
rect 2866 25644 2872 25696
rect 2924 25684 2930 25696
rect 3881 25687 3939 25693
rect 3881 25684 3893 25687
rect 2924 25656 3893 25684
rect 2924 25644 2930 25656
rect 3881 25653 3893 25656
rect 3927 25653 3939 25687
rect 3881 25647 3939 25653
rect 4062 25644 4068 25696
rect 4120 25684 4126 25696
rect 9858 25684 9864 25696
rect 4120 25656 9864 25684
rect 4120 25644 4126 25656
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 10152 25693 10180 25724
rect 10318 25712 10324 25724
rect 10376 25712 10382 25764
rect 13630 25712 13636 25764
rect 13688 25752 13694 25764
rect 14001 25755 14059 25761
rect 14001 25752 14013 25755
rect 13688 25724 14013 25752
rect 13688 25712 13694 25724
rect 14001 25721 14013 25724
rect 14047 25721 14059 25755
rect 14001 25715 14059 25721
rect 14185 25755 14243 25761
rect 14185 25721 14197 25755
rect 14231 25752 14243 25755
rect 14274 25752 14280 25764
rect 14231 25724 14280 25752
rect 14231 25721 14243 25724
rect 14185 25715 14243 25721
rect 14274 25712 14280 25724
rect 14332 25712 14338 25764
rect 14936 25752 14964 25783
rect 15102 25780 15108 25792
rect 15160 25780 15166 25832
rect 15562 25820 15568 25832
rect 15523 25792 15568 25820
rect 15562 25780 15568 25792
rect 15620 25780 15626 25832
rect 16206 25820 16212 25832
rect 16167 25792 16212 25820
rect 16206 25780 16212 25792
rect 16264 25780 16270 25832
rect 17865 25823 17923 25829
rect 17865 25789 17877 25823
rect 17911 25820 17923 25823
rect 17954 25820 17960 25832
rect 17911 25792 17960 25820
rect 17911 25789 17923 25792
rect 17865 25783 17923 25789
rect 17954 25780 17960 25792
rect 18012 25780 18018 25832
rect 18874 25829 18880 25832
rect 18865 25823 18880 25829
rect 18865 25789 18877 25823
rect 18865 25783 18880 25789
rect 18874 25780 18880 25783
rect 18932 25780 18938 25832
rect 19065 25823 19123 25829
rect 19065 25789 19077 25823
rect 19111 25789 19123 25823
rect 19065 25783 19123 25789
rect 19153 25823 19211 25829
rect 19153 25789 19165 25823
rect 19199 25789 19211 25823
rect 19153 25783 19211 25789
rect 19429 25823 19487 25829
rect 19429 25789 19441 25823
rect 19475 25820 19487 25823
rect 20162 25820 20168 25832
rect 19475 25792 20168 25820
rect 19475 25789 19487 25792
rect 19429 25783 19487 25789
rect 18506 25752 18512 25764
rect 14936 25724 18512 25752
rect 18506 25712 18512 25724
rect 18564 25712 18570 25764
rect 18966 25712 18972 25764
rect 19024 25752 19030 25764
rect 19076 25752 19104 25783
rect 19024 25724 19104 25752
rect 19024 25712 19030 25724
rect 10137 25687 10195 25693
rect 10137 25653 10149 25687
rect 10183 25653 10195 25687
rect 10137 25647 10195 25653
rect 12710 25644 12716 25696
rect 12768 25684 12774 25696
rect 13449 25687 13507 25693
rect 13449 25684 13461 25687
rect 12768 25656 13461 25684
rect 12768 25644 12774 25656
rect 13449 25653 13461 25656
rect 13495 25653 13507 25687
rect 13449 25647 13507 25653
rect 15378 25644 15384 25696
rect 15436 25684 15442 25696
rect 16301 25687 16359 25693
rect 16301 25684 16313 25687
rect 15436 25656 16313 25684
rect 15436 25644 15442 25656
rect 16301 25653 16313 25656
rect 16347 25684 16359 25687
rect 16942 25684 16948 25696
rect 16347 25656 16948 25684
rect 16347 25653 16359 25656
rect 16301 25647 16359 25653
rect 16942 25644 16948 25656
rect 17000 25644 17006 25696
rect 17310 25644 17316 25696
rect 17368 25684 17374 25696
rect 18230 25684 18236 25696
rect 17368 25656 18236 25684
rect 17368 25644 17374 25656
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 18417 25687 18475 25693
rect 18417 25653 18429 25687
rect 18463 25684 18475 25687
rect 18598 25684 18604 25696
rect 18463 25656 18604 25684
rect 18463 25653 18475 25656
rect 18417 25647 18475 25653
rect 18598 25644 18604 25656
rect 18656 25644 18662 25696
rect 18782 25644 18788 25696
rect 18840 25684 18846 25696
rect 19168 25684 19196 25783
rect 20162 25780 20168 25792
rect 20220 25780 20226 25832
rect 20349 25823 20407 25829
rect 20349 25789 20361 25823
rect 20395 25820 20407 25823
rect 20990 25820 20996 25832
rect 20395 25792 20996 25820
rect 20395 25789 20407 25792
rect 20349 25783 20407 25789
rect 20990 25780 20996 25792
rect 21048 25780 21054 25832
rect 21085 25823 21143 25829
rect 21085 25789 21097 25823
rect 21131 25820 21143 25823
rect 21358 25820 21364 25832
rect 21131 25792 21364 25820
rect 21131 25789 21143 25792
rect 21085 25783 21143 25789
rect 21358 25780 21364 25792
rect 21416 25780 21422 25832
rect 21450 25780 21456 25832
rect 21508 25820 21514 25832
rect 22278 25820 22284 25832
rect 21508 25792 22284 25820
rect 21508 25780 21514 25792
rect 22278 25780 22284 25792
rect 22336 25780 22342 25832
rect 22646 25780 22652 25832
rect 22704 25820 22710 25832
rect 23290 25820 23296 25832
rect 22704 25792 23296 25820
rect 22704 25780 22710 25792
rect 23290 25780 23296 25792
rect 23348 25820 23354 25832
rect 24121 25823 24179 25829
rect 24121 25820 24133 25823
rect 23348 25792 24133 25820
rect 23348 25780 23354 25792
rect 24121 25789 24133 25792
rect 24167 25789 24179 25823
rect 25958 25820 25964 25832
rect 25919 25792 25964 25820
rect 24121 25783 24179 25789
rect 25958 25780 25964 25792
rect 26016 25780 26022 25832
rect 26142 25820 26148 25832
rect 26103 25792 26148 25820
rect 26142 25780 26148 25792
rect 26200 25780 26206 25832
rect 26234 25780 26240 25832
rect 26292 25820 26298 25832
rect 26510 25820 26516 25832
rect 26292 25792 26337 25820
rect 26471 25792 26516 25820
rect 26292 25780 26298 25792
rect 26510 25780 26516 25792
rect 26568 25780 26574 25832
rect 28258 25780 28264 25832
rect 28316 25820 28322 25832
rect 29273 25823 29331 25829
rect 29273 25820 29285 25823
rect 28316 25792 29285 25820
rect 28316 25780 28322 25792
rect 29273 25789 29285 25792
rect 29319 25789 29331 25823
rect 29273 25783 29331 25789
rect 30009 25823 30067 25829
rect 30009 25789 30021 25823
rect 30055 25820 30067 25823
rect 30282 25820 30288 25832
rect 30055 25792 30288 25820
rect 30055 25789 30067 25792
rect 30009 25783 30067 25789
rect 30282 25780 30288 25792
rect 30340 25780 30346 25832
rect 31036 25829 31064 25860
rect 32122 25848 32128 25860
rect 32180 25848 32186 25900
rect 32582 25848 32588 25900
rect 32640 25888 32646 25900
rect 34330 25888 34336 25900
rect 32640 25860 33272 25888
rect 34291 25860 34336 25888
rect 32640 25848 32646 25860
rect 30929 25823 30987 25829
rect 30929 25789 30941 25823
rect 30975 25789 30987 25823
rect 30929 25783 30987 25789
rect 31021 25823 31079 25829
rect 31021 25789 31033 25823
rect 31067 25789 31079 25823
rect 31021 25783 31079 25789
rect 24388 25755 24446 25761
rect 24388 25721 24400 25755
rect 24434 25752 24446 25755
rect 26697 25755 26755 25761
rect 26697 25752 26709 25755
rect 24434 25724 26709 25752
rect 24434 25721 24446 25724
rect 24388 25715 24446 25721
rect 26697 25721 26709 25724
rect 26743 25721 26755 25755
rect 26697 25715 26755 25721
rect 27893 25755 27951 25761
rect 27893 25721 27905 25755
rect 27939 25752 27951 25755
rect 28629 25755 28687 25761
rect 28629 25752 28641 25755
rect 27939 25724 28641 25752
rect 27939 25721 27951 25724
rect 27893 25715 27951 25721
rect 28629 25721 28641 25724
rect 28675 25721 28687 25755
rect 28629 25715 28687 25721
rect 28813 25755 28871 25761
rect 28813 25721 28825 25755
rect 28859 25752 28871 25755
rect 29638 25752 29644 25764
rect 28859 25724 29644 25752
rect 28859 25721 28871 25724
rect 28813 25715 28871 25721
rect 18840 25656 19196 25684
rect 21637 25687 21695 25693
rect 18840 25644 18846 25656
rect 21637 25653 21649 25687
rect 21683 25684 21695 25687
rect 22186 25684 22192 25696
rect 21683 25656 22192 25684
rect 21683 25653 21695 25656
rect 21637 25647 21695 25653
rect 22186 25644 22192 25656
rect 22244 25644 22250 25696
rect 24578 25644 24584 25696
rect 24636 25684 24642 25696
rect 27908 25684 27936 25715
rect 29638 25712 29644 25724
rect 29696 25712 29702 25764
rect 24636 25656 27936 25684
rect 27985 25687 28043 25693
rect 24636 25644 24642 25656
rect 27985 25653 27997 25687
rect 28031 25684 28043 25687
rect 29822 25684 29828 25696
rect 28031 25656 29828 25684
rect 28031 25653 28043 25656
rect 27985 25647 28043 25653
rect 29822 25644 29828 25656
rect 29880 25684 29886 25696
rect 30466 25684 30472 25696
rect 29880 25656 30472 25684
rect 29880 25644 29886 25656
rect 30466 25644 30472 25656
rect 30524 25644 30530 25696
rect 30944 25684 30972 25783
rect 31202 25780 31208 25832
rect 31260 25820 31266 25832
rect 31757 25823 31815 25829
rect 31260 25792 31305 25820
rect 31260 25780 31266 25792
rect 31757 25789 31769 25823
rect 31803 25820 31815 25823
rect 31846 25820 31852 25832
rect 31803 25792 31852 25820
rect 31803 25789 31815 25792
rect 31757 25783 31815 25789
rect 31846 25780 31852 25792
rect 31904 25780 31910 25832
rect 31941 25823 31999 25829
rect 31941 25789 31953 25823
rect 31987 25820 31999 25823
rect 32398 25820 32404 25832
rect 31987 25792 32404 25820
rect 31987 25789 31999 25792
rect 31941 25783 31999 25789
rect 32398 25780 32404 25792
rect 32456 25780 32462 25832
rect 33244 25829 33272 25860
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 36630 25888 36636 25900
rect 36591 25860 36636 25888
rect 36630 25848 36636 25860
rect 36688 25848 36694 25900
rect 33229 25823 33287 25829
rect 33229 25789 33241 25823
rect 33275 25789 33287 25823
rect 33229 25783 33287 25789
rect 33321 25823 33379 25829
rect 33321 25789 33333 25823
rect 33367 25789 33379 25823
rect 33321 25783 33379 25789
rect 33597 25823 33655 25829
rect 33597 25789 33609 25823
rect 33643 25789 33655 25823
rect 34054 25820 34060 25832
rect 33967 25792 34060 25820
rect 33597 25783 33655 25789
rect 32674 25712 32680 25764
rect 32732 25752 32738 25764
rect 33336 25752 33364 25783
rect 32732 25724 33364 25752
rect 33612 25752 33640 25783
rect 34054 25780 34060 25792
rect 34112 25820 34118 25832
rect 34790 25820 34796 25832
rect 34112 25792 34796 25820
rect 34112 25780 34118 25792
rect 34790 25780 34796 25792
rect 34848 25780 34854 25832
rect 35618 25820 35624 25832
rect 35579 25792 35624 25820
rect 35618 25780 35624 25792
rect 35676 25780 35682 25832
rect 36354 25820 36360 25832
rect 36315 25792 36360 25820
rect 36354 25780 36360 25792
rect 36412 25780 36418 25832
rect 36449 25823 36507 25829
rect 36449 25789 36461 25823
rect 36495 25789 36507 25823
rect 36449 25783 36507 25789
rect 55493 25823 55551 25829
rect 55493 25789 55505 25823
rect 55539 25820 55551 25823
rect 55674 25820 55680 25832
rect 55539 25792 55680 25820
rect 55539 25789 55551 25792
rect 55493 25783 55551 25789
rect 33612 25724 34468 25752
rect 32732 25712 32738 25724
rect 34440 25696 34468 25724
rect 35986 25712 35992 25764
rect 36044 25752 36050 25764
rect 36464 25752 36492 25783
rect 55674 25780 55680 25792
rect 55732 25820 55738 25832
rect 56137 25823 56195 25829
rect 56137 25820 56149 25823
rect 55732 25792 56149 25820
rect 55732 25780 55738 25792
rect 56137 25789 56149 25792
rect 56183 25789 56195 25823
rect 56137 25783 56195 25789
rect 56502 25780 56508 25832
rect 56560 25820 56566 25832
rect 56597 25823 56655 25829
rect 56597 25820 56609 25823
rect 56560 25792 56609 25820
rect 56560 25780 56566 25792
rect 56597 25789 56609 25792
rect 56643 25789 56655 25823
rect 56597 25783 56655 25789
rect 56870 25780 56876 25832
rect 56928 25820 56934 25832
rect 57241 25823 57299 25829
rect 57241 25820 57253 25823
rect 56928 25792 57253 25820
rect 56928 25780 56934 25792
rect 57241 25789 57253 25792
rect 57287 25820 57299 25823
rect 57606 25820 57612 25832
rect 57287 25792 57612 25820
rect 57287 25789 57299 25792
rect 57241 25783 57299 25789
rect 57606 25780 57612 25792
rect 57664 25780 57670 25832
rect 57977 25823 58035 25829
rect 57977 25789 57989 25823
rect 58023 25820 58035 25823
rect 58250 25820 58256 25832
rect 58023 25792 58256 25820
rect 58023 25789 58035 25792
rect 57977 25783 58035 25789
rect 58250 25780 58256 25792
rect 58308 25780 58314 25832
rect 58158 25752 58164 25764
rect 36044 25724 36492 25752
rect 58119 25724 58164 25752
rect 36044 25712 36050 25724
rect 58158 25712 58164 25724
rect 58216 25712 58222 25764
rect 31294 25684 31300 25696
rect 30944 25656 31300 25684
rect 31294 25644 31300 25656
rect 31352 25684 31358 25696
rect 32125 25687 32183 25693
rect 32125 25684 32137 25687
rect 31352 25656 32137 25684
rect 31352 25644 31358 25656
rect 32125 25653 32137 25656
rect 32171 25653 32183 25687
rect 32125 25647 32183 25653
rect 33134 25644 33140 25696
rect 33192 25684 33198 25696
rect 34333 25687 34391 25693
rect 34333 25684 34345 25687
rect 33192 25656 34345 25684
rect 33192 25644 33198 25656
rect 34333 25653 34345 25656
rect 34379 25653 34391 25687
rect 34333 25647 34391 25653
rect 34422 25644 34428 25696
rect 34480 25644 34486 25696
rect 34514 25644 34520 25696
rect 34572 25684 34578 25696
rect 35713 25687 35771 25693
rect 35713 25684 35725 25687
rect 34572 25656 35725 25684
rect 34572 25644 34578 25656
rect 35713 25653 35725 25656
rect 35759 25684 35771 25687
rect 35802 25684 35808 25696
rect 35759 25656 35808 25684
rect 35759 25653 35771 25656
rect 35713 25647 35771 25653
rect 35802 25644 35808 25656
rect 35860 25644 35866 25696
rect 57054 25644 57060 25696
rect 57112 25684 57118 25696
rect 57422 25684 57428 25696
rect 57112 25656 57428 25684
rect 57112 25644 57118 25656
rect 57422 25644 57428 25656
rect 57480 25644 57486 25696
rect 1104 25594 58880 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 50326 25594
rect 50378 25542 50390 25594
rect 50442 25542 50454 25594
rect 50506 25542 50518 25594
rect 50570 25542 58880 25594
rect 1104 25520 58880 25542
rect 5166 25480 5172 25492
rect 5127 25452 5172 25480
rect 5166 25440 5172 25452
rect 5224 25440 5230 25492
rect 6822 25480 6828 25492
rect 5828 25452 6828 25480
rect 5828 25412 5856 25452
rect 6822 25440 6828 25452
rect 6880 25440 6886 25492
rect 6914 25440 6920 25492
rect 6972 25480 6978 25492
rect 7469 25483 7527 25489
rect 7469 25480 7481 25483
rect 6972 25452 7481 25480
rect 6972 25440 6978 25452
rect 7469 25449 7481 25452
rect 7515 25449 7527 25483
rect 17954 25480 17960 25492
rect 7469 25443 7527 25449
rect 7668 25452 15792 25480
rect 17915 25452 17960 25480
rect 7558 25412 7564 25424
rect 3160 25384 5856 25412
rect 5920 25384 7564 25412
rect 1854 25344 1860 25356
rect 1815 25316 1860 25344
rect 1854 25304 1860 25316
rect 1912 25304 1918 25356
rect 3160 25353 3188 25384
rect 3145 25347 3203 25353
rect 3145 25313 3157 25347
rect 3191 25313 3203 25347
rect 3145 25307 3203 25313
rect 3602 25304 3608 25356
rect 3660 25344 3666 25356
rect 4062 25344 4068 25356
rect 3660 25316 4068 25344
rect 3660 25304 3666 25316
rect 4062 25304 4068 25316
rect 4120 25344 4126 25356
rect 4249 25347 4307 25353
rect 4249 25344 4261 25347
rect 4120 25316 4261 25344
rect 4120 25304 4126 25316
rect 4249 25313 4261 25316
rect 4295 25313 4307 25347
rect 4249 25307 4307 25313
rect 4433 25347 4491 25353
rect 4433 25313 4445 25347
rect 4479 25313 4491 25347
rect 4433 25307 4491 25313
rect 5077 25347 5135 25353
rect 5077 25313 5089 25347
rect 5123 25313 5135 25347
rect 5258 25344 5264 25356
rect 5171 25316 5264 25344
rect 5077 25307 5135 25313
rect 2961 25279 3019 25285
rect 2961 25245 2973 25279
rect 3007 25276 3019 25279
rect 3620 25276 3648 25304
rect 3007 25248 3648 25276
rect 3007 25245 3019 25248
rect 2961 25239 3019 25245
rect 4448 25208 4476 25307
rect 5092 25276 5120 25307
rect 5258 25304 5264 25316
rect 5316 25344 5322 25356
rect 5920 25353 5948 25384
rect 7558 25372 7564 25384
rect 7616 25372 7622 25424
rect 5905 25347 5963 25353
rect 5316 25316 5856 25344
rect 5316 25304 5322 25316
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5092 25248 5733 25276
rect 5721 25245 5733 25248
rect 5767 25245 5779 25279
rect 5828 25276 5856 25316
rect 5905 25313 5917 25347
rect 5951 25313 5963 25347
rect 5905 25307 5963 25313
rect 5994 25304 6000 25356
rect 6052 25344 6058 25356
rect 6052 25316 6097 25344
rect 6052 25304 6058 25316
rect 6178 25304 6184 25356
rect 6236 25344 6242 25356
rect 7668 25353 7696 25452
rect 7834 25412 7840 25424
rect 7747 25384 7840 25412
rect 7760 25353 7788 25384
rect 7834 25372 7840 25384
rect 7892 25412 7898 25424
rect 9766 25412 9772 25424
rect 7892 25384 9772 25412
rect 7892 25372 7898 25384
rect 9766 25372 9772 25384
rect 9824 25372 9830 25424
rect 11048 25415 11106 25421
rect 11048 25381 11060 25415
rect 11094 25412 11106 25415
rect 11698 25412 11704 25424
rect 11094 25384 11704 25412
rect 11094 25381 11106 25384
rect 11048 25375 11106 25381
rect 11698 25372 11704 25384
rect 11756 25372 11762 25424
rect 13630 25412 13636 25424
rect 13591 25384 13636 25412
rect 13630 25372 13636 25384
rect 13688 25372 13694 25424
rect 6273 25347 6331 25353
rect 6273 25344 6285 25347
rect 6236 25316 6285 25344
rect 6236 25304 6242 25316
rect 6273 25313 6285 25316
rect 6319 25313 6331 25347
rect 6273 25307 6331 25313
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7653 25347 7711 25353
rect 6871 25316 7604 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 7006 25276 7012 25288
rect 5828 25248 7012 25276
rect 5721 25239 5779 25245
rect 7006 25236 7012 25248
rect 7064 25236 7070 25288
rect 7576 25276 7604 25316
rect 7653 25313 7665 25347
rect 7699 25313 7711 25347
rect 7653 25307 7711 25313
rect 7745 25347 7803 25353
rect 7745 25313 7757 25347
rect 7791 25313 7803 25347
rect 8018 25344 8024 25356
rect 7979 25316 8024 25344
rect 7745 25307 7803 25313
rect 8018 25304 8024 25316
rect 8076 25304 8082 25356
rect 9582 25344 9588 25356
rect 9543 25316 9588 25344
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 12710 25344 12716 25356
rect 9692 25316 12716 25344
rect 8386 25276 8392 25288
rect 7576 25248 8392 25276
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 9692 25208 9720 25316
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 12897 25347 12955 25353
rect 12897 25313 12909 25347
rect 12943 25344 12955 25347
rect 14642 25344 14648 25356
rect 12943 25316 14648 25344
rect 12943 25313 12955 25316
rect 12897 25307 12955 25313
rect 14642 25304 14648 25316
rect 14700 25304 14706 25356
rect 14826 25304 14832 25356
rect 14884 25344 14890 25356
rect 14921 25347 14979 25353
rect 14921 25344 14933 25347
rect 14884 25316 14933 25344
rect 14884 25304 14890 25316
rect 14921 25313 14933 25316
rect 14967 25313 14979 25347
rect 14921 25307 14979 25313
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25245 10839 25279
rect 12989 25279 13047 25285
rect 12989 25276 13001 25279
rect 10781 25239 10839 25245
rect 11808 25248 13001 25276
rect 4448 25180 9720 25208
rect 1946 25140 1952 25152
rect 1907 25112 1952 25140
rect 1946 25100 1952 25112
rect 2004 25100 2010 25152
rect 3326 25140 3332 25152
rect 3287 25112 3332 25140
rect 3326 25100 3332 25112
rect 3384 25100 3390 25152
rect 4614 25140 4620 25152
rect 4575 25112 4620 25140
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 6181 25143 6239 25149
rect 6181 25109 6193 25143
rect 6227 25140 6239 25143
rect 6546 25140 6552 25152
rect 6227 25112 6552 25140
rect 6227 25109 6239 25112
rect 6181 25103 6239 25109
rect 6546 25100 6552 25112
rect 6604 25100 6610 25152
rect 6822 25100 6828 25152
rect 6880 25140 6886 25152
rect 7650 25140 7656 25152
rect 6880 25112 7656 25140
rect 6880 25100 6886 25112
rect 7650 25100 7656 25112
rect 7708 25100 7714 25152
rect 7926 25140 7932 25152
rect 7887 25112 7932 25140
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 10796 25140 10824 25239
rect 11054 25140 11060 25152
rect 10796 25112 11060 25140
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11808 25140 11836 25248
rect 12989 25245 13001 25248
rect 13035 25276 13047 25279
rect 15654 25276 15660 25288
rect 13035 25248 15660 25276
rect 13035 25245 13047 25248
rect 12989 25239 13047 25245
rect 15654 25236 15660 25248
rect 15712 25236 15718 25288
rect 15764 25276 15792 25452
rect 17954 25440 17960 25452
rect 18012 25440 18018 25492
rect 18138 25440 18144 25492
rect 18196 25480 18202 25492
rect 21358 25480 21364 25492
rect 18196 25452 21220 25480
rect 21319 25452 21364 25480
rect 18196 25440 18202 25452
rect 16298 25372 16304 25424
rect 16356 25412 16362 25424
rect 16485 25415 16543 25421
rect 16485 25412 16497 25415
rect 16356 25384 16497 25412
rect 16356 25372 16362 25384
rect 16485 25381 16497 25384
rect 16531 25412 16543 25415
rect 18506 25412 18512 25424
rect 16531 25384 18267 25412
rect 16531 25381 16543 25384
rect 16485 25375 16543 25381
rect 15841 25347 15899 25353
rect 15841 25313 15853 25347
rect 15887 25344 15899 25347
rect 16206 25344 16212 25356
rect 15887 25316 16212 25344
rect 15887 25313 15899 25316
rect 15841 25307 15899 25313
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 16666 25344 16672 25356
rect 16627 25316 16672 25344
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 16761 25347 16819 25353
rect 16761 25313 16773 25347
rect 16807 25344 16819 25347
rect 16850 25344 16856 25356
rect 16807 25316 16856 25344
rect 16807 25313 16819 25316
rect 16761 25307 16819 25313
rect 16850 25304 16856 25316
rect 16908 25304 16914 25356
rect 17310 25344 17316 25356
rect 17271 25316 17316 25344
rect 17310 25304 17316 25316
rect 17368 25304 17374 25356
rect 18239 25353 18267 25384
rect 18340 25384 18512 25412
rect 18340 25353 18368 25384
rect 18506 25372 18512 25384
rect 18564 25372 18570 25424
rect 20248 25415 20306 25421
rect 20248 25381 20260 25415
rect 20294 25412 20306 25415
rect 20622 25412 20628 25424
rect 20294 25384 20628 25412
rect 20294 25381 20306 25384
rect 20248 25375 20306 25381
rect 20622 25372 20628 25384
rect 20680 25372 20686 25424
rect 21192 25412 21220 25452
rect 21358 25440 21364 25452
rect 21416 25440 21422 25492
rect 22186 25480 22192 25492
rect 21468 25452 22192 25480
rect 21468 25412 21496 25452
rect 22186 25440 22192 25452
rect 22244 25480 22250 25492
rect 22830 25480 22836 25492
rect 22244 25452 22836 25480
rect 22244 25440 22250 25452
rect 22830 25440 22836 25452
rect 22888 25440 22894 25492
rect 23201 25483 23259 25489
rect 23201 25449 23213 25483
rect 23247 25480 23259 25483
rect 23474 25480 23480 25492
rect 23247 25452 23480 25480
rect 23247 25449 23259 25452
rect 23201 25443 23259 25449
rect 23474 25440 23480 25452
rect 23532 25440 23538 25492
rect 28258 25480 28264 25492
rect 25516 25452 26648 25480
rect 28219 25452 28264 25480
rect 21192 25384 21496 25412
rect 21634 25372 21640 25424
rect 21692 25412 21698 25424
rect 22066 25415 22124 25421
rect 22066 25412 22078 25415
rect 21692 25384 22078 25412
rect 21692 25372 21698 25384
rect 22066 25381 22078 25384
rect 22112 25381 22124 25415
rect 22066 25375 22124 25381
rect 22370 25372 22376 25424
rect 22428 25412 22434 25424
rect 24121 25415 24179 25421
rect 24121 25412 24133 25415
rect 22428 25384 24133 25412
rect 22428 25372 22434 25384
rect 24121 25381 24133 25384
rect 24167 25381 24179 25415
rect 25516 25412 25544 25452
rect 26510 25412 26516 25424
rect 24121 25375 24179 25381
rect 25424 25384 25544 25412
rect 25792 25384 26516 25412
rect 18233 25347 18291 25353
rect 18233 25313 18245 25347
rect 18279 25313 18291 25347
rect 18233 25307 18291 25313
rect 18325 25347 18383 25353
rect 18325 25313 18337 25347
rect 18371 25313 18383 25347
rect 18325 25307 18383 25313
rect 18414 25304 18420 25356
rect 18472 25353 18478 25356
rect 18472 25344 18480 25353
rect 18601 25347 18659 25353
rect 18472 25316 18517 25344
rect 18472 25307 18480 25316
rect 18601 25313 18613 25347
rect 18647 25344 18659 25347
rect 18874 25344 18880 25356
rect 18647 25316 18880 25344
rect 18647 25313 18659 25316
rect 18601 25307 18659 25313
rect 18472 25304 18478 25307
rect 18874 25304 18880 25316
rect 18932 25344 18938 25356
rect 22388 25344 22416 25372
rect 18932 25316 22416 25344
rect 18932 25304 18938 25316
rect 23566 25304 23572 25356
rect 23624 25344 23630 25356
rect 25424 25353 25452 25384
rect 23937 25347 23995 25353
rect 23937 25344 23949 25347
rect 23624 25316 23949 25344
rect 23624 25304 23630 25316
rect 23937 25313 23949 25316
rect 23983 25313 23995 25347
rect 23937 25307 23995 25313
rect 25225 25347 25283 25353
rect 25225 25313 25237 25347
rect 25271 25313 25283 25347
rect 25225 25307 25283 25313
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25313 25467 25347
rect 25409 25307 25467 25313
rect 17494 25276 17500 25288
rect 15764 25248 17500 25276
rect 17494 25236 17500 25248
rect 17552 25236 17558 25288
rect 17586 25236 17592 25288
rect 17644 25276 17650 25288
rect 19981 25279 20039 25285
rect 19981 25276 19993 25279
rect 17644 25248 19993 25276
rect 17644 25236 17650 25248
rect 19981 25245 19993 25248
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 21542 25236 21548 25288
rect 21600 25276 21606 25288
rect 21821 25279 21879 25285
rect 21821 25276 21833 25279
rect 21600 25248 21833 25276
rect 21600 25236 21606 25248
rect 21821 25245 21833 25248
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 15562 25208 15568 25220
rect 13740 25180 15568 25208
rect 12158 25140 12164 25152
rect 11204 25112 11836 25140
rect 12119 25112 12164 25140
rect 11204 25100 11210 25112
rect 12158 25100 12164 25112
rect 12216 25100 12222 25152
rect 13446 25100 13452 25152
rect 13504 25140 13510 25152
rect 13740 25149 13768 25180
rect 15562 25168 15568 25180
rect 15620 25168 15626 25220
rect 15933 25211 15991 25217
rect 15933 25177 15945 25211
rect 15979 25208 15991 25211
rect 19886 25208 19892 25220
rect 15979 25180 19892 25208
rect 15979 25177 15991 25180
rect 15933 25171 15991 25177
rect 19886 25168 19892 25180
rect 19944 25168 19950 25220
rect 25240 25208 25268 25307
rect 25498 25304 25504 25356
rect 25556 25344 25562 25356
rect 25792 25353 25820 25384
rect 26510 25372 26516 25384
rect 26568 25372 26574 25424
rect 25777 25347 25835 25353
rect 25556 25316 25601 25344
rect 25556 25304 25562 25316
rect 25777 25313 25789 25347
rect 25823 25313 25835 25347
rect 26620 25344 26648 25452
rect 28258 25440 28264 25452
rect 28316 25440 28322 25492
rect 31202 25440 31208 25492
rect 31260 25480 31266 25492
rect 31849 25483 31907 25489
rect 31849 25480 31861 25483
rect 31260 25452 31861 25480
rect 31260 25440 31266 25452
rect 31849 25449 31861 25452
rect 31895 25449 31907 25483
rect 32306 25480 32312 25492
rect 32267 25452 32312 25480
rect 31849 25443 31907 25449
rect 32306 25440 32312 25452
rect 32364 25440 32370 25492
rect 34330 25480 34336 25492
rect 34291 25452 34336 25480
rect 34330 25440 34336 25452
rect 34388 25440 34394 25492
rect 34422 25440 34428 25492
rect 34480 25480 34486 25492
rect 34480 25452 37412 25480
rect 34480 25440 34486 25452
rect 27148 25415 27206 25421
rect 27148 25381 27160 25415
rect 27194 25412 27206 25415
rect 29914 25412 29920 25424
rect 27194 25384 29920 25412
rect 27194 25381 27206 25384
rect 27148 25375 27206 25381
rect 29914 25372 29920 25384
rect 29972 25372 29978 25424
rect 30558 25372 30564 25424
rect 30616 25412 30622 25424
rect 30616 25384 35756 25412
rect 30616 25372 30622 25384
rect 26620 25316 27936 25344
rect 25777 25307 25835 25313
rect 25593 25279 25651 25285
rect 25593 25245 25605 25279
rect 25639 25276 25651 25279
rect 26786 25276 26792 25288
rect 25639 25248 26792 25276
rect 25639 25245 25651 25248
rect 25593 25239 25651 25245
rect 26786 25236 26792 25248
rect 26844 25236 26850 25288
rect 26881 25279 26939 25285
rect 26881 25245 26893 25279
rect 26927 25245 26939 25279
rect 27908 25276 27936 25316
rect 27982 25304 27988 25356
rect 28040 25344 28046 25356
rect 28813 25347 28871 25353
rect 28813 25344 28825 25347
rect 28040 25316 28825 25344
rect 28040 25304 28046 25316
rect 28813 25313 28825 25316
rect 28859 25313 28871 25347
rect 28813 25307 28871 25313
rect 28997 25347 29055 25353
rect 28997 25313 29009 25347
rect 29043 25313 29055 25347
rect 28997 25307 29055 25313
rect 28718 25276 28724 25288
rect 27908 25248 28724 25276
rect 26881 25239 26939 25245
rect 25240 25180 26096 25208
rect 26068 25152 26096 25180
rect 26510 25168 26516 25220
rect 26568 25208 26574 25220
rect 26896 25208 26924 25239
rect 28718 25236 28724 25248
rect 28776 25276 28782 25288
rect 29012 25276 29040 25307
rect 29270 25304 29276 25356
rect 29328 25344 29334 25356
rect 29365 25347 29423 25353
rect 29365 25344 29377 25347
rect 29328 25316 29377 25344
rect 29328 25304 29334 25316
rect 29365 25313 29377 25316
rect 29411 25313 29423 25347
rect 30466 25344 30472 25356
rect 30427 25316 30472 25344
rect 29365 25307 29423 25313
rect 30466 25304 30472 25316
rect 30524 25304 30530 25356
rect 30926 25304 30932 25356
rect 30984 25344 30990 25356
rect 31113 25347 31171 25353
rect 31113 25344 31125 25347
rect 30984 25316 31125 25344
rect 30984 25304 30990 25316
rect 31113 25313 31125 25316
rect 31159 25313 31171 25347
rect 31294 25344 31300 25356
rect 31255 25316 31300 25344
rect 31113 25307 31171 25313
rect 31294 25304 31300 25316
rect 31352 25304 31358 25356
rect 31665 25347 31723 25353
rect 31665 25313 31677 25347
rect 31711 25344 31723 25347
rect 31846 25344 31852 25356
rect 31711 25316 31852 25344
rect 31711 25313 31723 25316
rect 31665 25307 31723 25313
rect 31846 25304 31852 25316
rect 31904 25304 31910 25356
rect 32398 25304 32404 25356
rect 32456 25344 32462 25356
rect 32493 25347 32551 25353
rect 32493 25344 32505 25347
rect 32456 25316 32505 25344
rect 32456 25304 32462 25316
rect 32493 25313 32505 25316
rect 32539 25313 32551 25347
rect 32493 25307 32551 25313
rect 32769 25347 32827 25353
rect 32769 25313 32781 25347
rect 32815 25344 32827 25347
rect 33134 25344 33140 25356
rect 32815 25316 33140 25344
rect 32815 25313 32827 25316
rect 32769 25307 32827 25313
rect 28776 25248 29040 25276
rect 29089 25279 29147 25285
rect 28776 25236 28782 25248
rect 29089 25245 29101 25279
rect 29135 25245 29147 25279
rect 29089 25239 29147 25245
rect 29181 25279 29239 25285
rect 29181 25245 29193 25279
rect 29227 25276 29239 25279
rect 30374 25276 30380 25288
rect 29227 25248 30380 25276
rect 29227 25245 29239 25248
rect 29181 25239 29239 25245
rect 26568 25180 26924 25208
rect 29104 25208 29132 25239
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 31389 25279 31447 25285
rect 31389 25245 31401 25279
rect 31435 25245 31447 25279
rect 31389 25239 31447 25245
rect 31481 25279 31539 25285
rect 31481 25245 31493 25279
rect 31527 25276 31539 25279
rect 32582 25276 32588 25288
rect 31527 25248 32444 25276
rect 32543 25248 32588 25276
rect 31527 25245 31539 25248
rect 31481 25239 31539 25245
rect 31294 25208 31300 25220
rect 29104 25180 31300 25208
rect 26568 25168 26574 25180
rect 31294 25168 31300 25180
rect 31352 25168 31358 25220
rect 31404 25208 31432 25239
rect 31754 25208 31760 25220
rect 31404 25180 31760 25208
rect 31754 25168 31760 25180
rect 31812 25168 31818 25220
rect 13725 25143 13783 25149
rect 13725 25140 13737 25143
rect 13504 25112 13737 25140
rect 13504 25100 13510 25112
rect 13725 25109 13737 25112
rect 13771 25109 13783 25143
rect 13725 25103 13783 25109
rect 15197 25143 15255 25149
rect 15197 25109 15209 25143
rect 15243 25140 15255 25143
rect 16114 25140 16120 25152
rect 15243 25112 16120 25140
rect 15243 25109 15255 25112
rect 15197 25103 15255 25109
rect 16114 25100 16120 25112
rect 16172 25100 16178 25152
rect 16485 25143 16543 25149
rect 16485 25109 16497 25143
rect 16531 25140 16543 25143
rect 16850 25140 16856 25152
rect 16531 25112 16856 25140
rect 16531 25109 16543 25112
rect 16485 25103 16543 25109
rect 16850 25100 16856 25112
rect 16908 25100 16914 25152
rect 17402 25140 17408 25152
rect 17363 25112 17408 25140
rect 17402 25100 17408 25112
rect 17460 25100 17466 25152
rect 17494 25100 17500 25152
rect 17552 25140 17558 25152
rect 22094 25140 22100 25152
rect 17552 25112 22100 25140
rect 17552 25100 17558 25112
rect 22094 25100 22100 25112
rect 22152 25100 22158 25152
rect 25774 25100 25780 25152
rect 25832 25140 25838 25152
rect 25961 25143 26019 25149
rect 25961 25140 25973 25143
rect 25832 25112 25973 25140
rect 25832 25100 25838 25112
rect 25961 25109 25973 25112
rect 26007 25109 26019 25143
rect 25961 25103 26019 25109
rect 26050 25100 26056 25152
rect 26108 25140 26114 25152
rect 27982 25140 27988 25152
rect 26108 25112 27988 25140
rect 26108 25100 26114 25112
rect 27982 25100 27988 25112
rect 28040 25100 28046 25152
rect 29362 25100 29368 25152
rect 29420 25140 29426 25152
rect 29549 25143 29607 25149
rect 29549 25140 29561 25143
rect 29420 25112 29561 25140
rect 29420 25100 29426 25112
rect 29549 25109 29561 25112
rect 29595 25109 29607 25143
rect 29549 25103 29607 25109
rect 30561 25143 30619 25149
rect 30561 25109 30573 25143
rect 30607 25140 30619 25143
rect 32030 25140 32036 25152
rect 30607 25112 32036 25140
rect 30607 25109 30619 25112
rect 30561 25103 30619 25109
rect 32030 25100 32036 25112
rect 32088 25100 32094 25152
rect 32416 25140 32444 25248
rect 32582 25236 32588 25248
rect 32640 25236 32646 25288
rect 32674 25236 32680 25288
rect 32732 25276 32738 25288
rect 32732 25248 32777 25276
rect 32732 25236 32738 25248
rect 32968 25140 32996 25316
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 33686 25304 33692 25356
rect 33744 25344 33750 25356
rect 33781 25347 33839 25353
rect 33781 25344 33793 25347
rect 33744 25316 33793 25344
rect 33744 25304 33750 25316
rect 33781 25313 33793 25316
rect 33827 25313 33839 25347
rect 33962 25344 33968 25356
rect 33923 25316 33968 25344
rect 33781 25307 33839 25313
rect 33962 25304 33968 25316
rect 34020 25304 34026 25356
rect 34054 25304 34060 25356
rect 34112 25344 34118 25356
rect 34238 25353 34244 25356
rect 34195 25347 34244 25353
rect 34112 25316 34157 25344
rect 34112 25304 34118 25316
rect 34195 25313 34207 25347
rect 34241 25313 34244 25347
rect 34195 25307 34244 25313
rect 34238 25304 34244 25307
rect 34296 25304 34302 25356
rect 35728 25353 35756 25384
rect 35713 25347 35771 25353
rect 35713 25313 35725 25347
rect 35759 25313 35771 25347
rect 36446 25344 36452 25356
rect 36407 25316 36452 25344
rect 35713 25307 35771 25313
rect 36446 25304 36452 25316
rect 36504 25304 36510 25356
rect 36538 25304 36544 25356
rect 36596 25344 36602 25356
rect 36596 25316 36641 25344
rect 36596 25304 36602 25316
rect 37090 25304 37096 25356
rect 37148 25344 37154 25356
rect 37384 25353 37412 25452
rect 55582 25440 55588 25492
rect 55640 25440 55646 25492
rect 57974 25480 57980 25492
rect 57935 25452 57980 25480
rect 57974 25440 57980 25452
rect 58032 25440 58038 25492
rect 55600 25412 55628 25440
rect 56318 25412 56324 25424
rect 55600 25384 56324 25412
rect 56318 25372 56324 25384
rect 56376 25412 56382 25424
rect 57149 25415 57207 25421
rect 57149 25412 57161 25415
rect 56376 25384 57161 25412
rect 56376 25372 56382 25384
rect 57149 25381 57161 25384
rect 57195 25381 57207 25415
rect 57149 25375 57207 25381
rect 37185 25347 37243 25353
rect 37185 25344 37197 25347
rect 37148 25316 37197 25344
rect 37148 25304 37154 25316
rect 37185 25313 37197 25316
rect 37231 25313 37243 25347
rect 37185 25307 37243 25313
rect 37369 25347 37427 25353
rect 37369 25313 37381 25347
rect 37415 25313 37427 25347
rect 37369 25307 37427 25313
rect 55585 25347 55643 25353
rect 55585 25313 55597 25347
rect 55631 25344 55643 25347
rect 55674 25344 55680 25356
rect 55631 25316 55680 25344
rect 55631 25313 55643 25316
rect 55585 25307 55643 25313
rect 36722 25276 36728 25288
rect 36683 25248 36728 25276
rect 36722 25236 36728 25248
rect 36780 25236 36786 25288
rect 36078 25168 36084 25220
rect 36136 25208 36142 25220
rect 37200 25208 37228 25307
rect 55674 25304 55680 25316
rect 55732 25304 55738 25356
rect 57422 25304 57428 25356
rect 57480 25344 57486 25356
rect 58161 25347 58219 25353
rect 58161 25344 58173 25347
rect 57480 25316 58173 25344
rect 57480 25304 57486 25316
rect 58161 25313 58173 25316
rect 58207 25313 58219 25347
rect 58161 25307 58219 25313
rect 36136 25180 37228 25208
rect 36136 25168 36142 25180
rect 32416 25112 32996 25140
rect 34606 25100 34612 25152
rect 34664 25140 34670 25152
rect 35805 25143 35863 25149
rect 35805 25140 35817 25143
rect 34664 25112 35817 25140
rect 34664 25100 34670 25112
rect 35805 25109 35817 25112
rect 35851 25109 35863 25143
rect 35805 25103 35863 25109
rect 35894 25100 35900 25152
rect 35952 25140 35958 25152
rect 37185 25143 37243 25149
rect 37185 25140 37197 25143
rect 35952 25112 37197 25140
rect 35952 25100 35958 25112
rect 37185 25109 37197 25112
rect 37231 25109 37243 25143
rect 55398 25140 55404 25152
rect 55359 25112 55404 25140
rect 37185 25103 37243 25109
rect 55398 25100 55404 25112
rect 55456 25100 55462 25152
rect 57238 25140 57244 25152
rect 57199 25112 57244 25140
rect 57238 25100 57244 25112
rect 57296 25100 57302 25152
rect 1104 25050 58880 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 58880 25050
rect 1104 24976 58880 24998
rect 1854 24896 1860 24948
rect 1912 24936 1918 24948
rect 2317 24939 2375 24945
rect 2317 24936 2329 24939
rect 1912 24908 2329 24936
rect 1912 24896 1918 24908
rect 2317 24905 2329 24908
rect 2363 24905 2375 24939
rect 2317 24899 2375 24905
rect 7300 24908 8432 24936
rect 4062 24868 4068 24880
rect 3528 24840 4068 24868
rect 1949 24803 2007 24809
rect 1949 24769 1961 24803
rect 1995 24800 2007 24803
rect 3326 24800 3332 24812
rect 1995 24772 3332 24800
rect 1995 24769 2007 24772
rect 1949 24763 2007 24769
rect 3326 24760 3332 24772
rect 3384 24760 3390 24812
rect 3528 24809 3556 24840
rect 4062 24828 4068 24840
rect 4120 24828 4126 24880
rect 3513 24803 3571 24809
rect 3513 24769 3525 24803
rect 3559 24769 3571 24803
rect 7300 24800 7328 24908
rect 8294 24828 8300 24880
rect 8352 24828 8358 24880
rect 8312 24800 8340 24828
rect 3513 24763 3571 24769
rect 3712 24772 7328 24800
rect 7392 24772 8340 24800
rect 8404 24800 8432 24908
rect 9582 24896 9588 24948
rect 9640 24936 9646 24948
rect 13446 24936 13452 24948
rect 9640 24908 13452 24936
rect 9640 24896 9646 24908
rect 13446 24896 13452 24908
rect 13504 24896 13510 24948
rect 13630 24936 13636 24948
rect 13591 24908 13636 24936
rect 13630 24896 13636 24908
rect 13688 24896 13694 24948
rect 14550 24896 14556 24948
rect 14608 24936 14614 24948
rect 14608 24908 15516 24936
rect 14608 24896 14614 24908
rect 11514 24868 11520 24880
rect 10428 24840 11520 24868
rect 10428 24800 10456 24840
rect 11514 24828 11520 24840
rect 11572 24868 11578 24880
rect 12158 24868 12164 24880
rect 11572 24840 12164 24868
rect 11572 24828 11578 24840
rect 12158 24828 12164 24840
rect 12216 24828 12222 24880
rect 15488 24868 15516 24908
rect 15654 24896 15660 24948
rect 15712 24936 15718 24948
rect 16758 24936 16764 24948
rect 15712 24908 16764 24936
rect 15712 24896 15718 24908
rect 16758 24896 16764 24908
rect 16816 24896 16822 24948
rect 17402 24896 17408 24948
rect 17460 24936 17466 24948
rect 21082 24936 21088 24948
rect 17460 24908 21088 24936
rect 17460 24896 17466 24908
rect 21082 24896 21088 24908
rect 21140 24936 21146 24948
rect 24578 24936 24584 24948
rect 21140 24908 24584 24936
rect 21140 24896 21146 24908
rect 24578 24896 24584 24908
rect 24636 24896 24642 24948
rect 26142 24936 26148 24948
rect 24872 24908 26148 24936
rect 17586 24868 17592 24880
rect 15488 24840 17592 24868
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 17681 24871 17739 24877
rect 17681 24837 17693 24871
rect 17727 24868 17739 24871
rect 17954 24868 17960 24880
rect 17727 24840 17960 24868
rect 17727 24837 17739 24840
rect 17681 24831 17739 24837
rect 17954 24828 17960 24840
rect 18012 24868 18018 24880
rect 18322 24868 18328 24880
rect 18012 24840 18328 24868
rect 18012 24828 18018 24840
rect 18322 24828 18328 24840
rect 18380 24828 18386 24880
rect 20162 24828 20168 24880
rect 20220 24868 20226 24880
rect 24121 24871 24179 24877
rect 24121 24868 24133 24871
rect 20220 24840 24133 24868
rect 20220 24828 20226 24840
rect 24121 24837 24133 24840
rect 24167 24868 24179 24871
rect 24486 24868 24492 24880
rect 24167 24840 24492 24868
rect 24167 24837 24179 24840
rect 24121 24831 24179 24837
rect 24486 24828 24492 24840
rect 24544 24828 24550 24880
rect 8404 24772 10456 24800
rect 10505 24803 10563 24809
rect 2133 24735 2191 24741
rect 2133 24701 2145 24735
rect 2179 24732 2191 24735
rect 3142 24732 3148 24744
rect 2179 24704 3148 24732
rect 2179 24701 2191 24704
rect 2133 24695 2191 24701
rect 3142 24692 3148 24704
rect 3200 24692 3206 24744
rect 3712 24741 3740 24772
rect 3697 24735 3755 24741
rect 3697 24701 3709 24735
rect 3743 24701 3755 24735
rect 3697 24695 3755 24701
rect 4709 24735 4767 24741
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 4893 24735 4951 24741
rect 4893 24701 4905 24735
rect 4939 24732 4951 24735
rect 4982 24732 4988 24744
rect 4939 24704 4988 24732
rect 4939 24701 4951 24704
rect 4893 24695 4951 24701
rect 4724 24664 4752 24695
rect 4982 24692 4988 24704
rect 5040 24732 5046 24744
rect 5258 24732 5264 24744
rect 5040 24704 5264 24732
rect 5040 24692 5046 24704
rect 5258 24692 5264 24704
rect 5316 24692 5322 24744
rect 5353 24735 5411 24741
rect 5353 24701 5365 24735
rect 5399 24732 5411 24735
rect 5626 24732 5632 24744
rect 5399 24704 5632 24732
rect 5399 24701 5411 24704
rect 5353 24695 5411 24701
rect 5626 24692 5632 24704
rect 5684 24692 5690 24744
rect 7392 24741 7420 24772
rect 10505 24769 10517 24803
rect 10551 24800 10563 24803
rect 10962 24800 10968 24812
rect 10551 24772 10968 24800
rect 10551 24769 10563 24772
rect 10505 24763 10563 24769
rect 10962 24760 10968 24772
rect 11020 24760 11026 24812
rect 12066 24760 12072 24812
rect 12124 24800 12130 24812
rect 14458 24800 14464 24812
rect 12124 24772 14464 24800
rect 12124 24760 12130 24772
rect 14458 24760 14464 24772
rect 14516 24760 14522 24812
rect 16666 24760 16672 24812
rect 16724 24800 16730 24812
rect 18138 24800 18144 24812
rect 16724 24772 18144 24800
rect 16724 24760 16730 24772
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 20530 24800 20536 24812
rect 20491 24772 20536 24800
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24800 21143 24803
rect 21818 24800 21824 24812
rect 21131 24772 21824 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 24872 24809 24900 24908
rect 26142 24896 26148 24908
rect 26200 24896 26206 24948
rect 26878 24936 26884 24948
rect 26839 24908 26884 24936
rect 26878 24896 26884 24908
rect 26936 24896 26942 24948
rect 30374 24896 30380 24948
rect 30432 24936 30438 24948
rect 30469 24939 30527 24945
rect 30469 24936 30481 24939
rect 30432 24908 30481 24936
rect 30432 24896 30438 24908
rect 30469 24905 30481 24908
rect 30515 24905 30527 24939
rect 32030 24936 32036 24948
rect 31943 24908 32036 24936
rect 30469 24899 30527 24905
rect 30484 24868 30512 24899
rect 32030 24896 32036 24908
rect 32088 24936 32094 24948
rect 32674 24936 32680 24948
rect 32088 24908 32680 24936
rect 32088 24896 32094 24908
rect 32674 24896 32680 24908
rect 32732 24896 32738 24948
rect 35986 24936 35992 24948
rect 33704 24908 35992 24936
rect 30484 24840 32720 24868
rect 24857 24803 24915 24809
rect 24857 24800 24869 24803
rect 22520 24772 24869 24800
rect 22520 24760 22526 24772
rect 24857 24769 24869 24772
rect 24903 24769 24915 24803
rect 24857 24763 24915 24769
rect 27798 24760 27804 24812
rect 27856 24800 27862 24812
rect 27856 24772 29040 24800
rect 27856 24760 27862 24772
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24701 7435 24735
rect 7377 24695 7435 24701
rect 8021 24735 8079 24741
rect 8021 24701 8033 24735
rect 8067 24732 8079 24735
rect 8202 24732 8208 24744
rect 8067 24704 8208 24732
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 8297 24735 8355 24741
rect 8297 24701 8309 24735
rect 8343 24701 8355 24735
rect 8297 24695 8355 24701
rect 6086 24664 6092 24676
rect 4724 24636 6092 24664
rect 6086 24624 6092 24636
rect 6144 24624 6150 24676
rect 7926 24624 7932 24676
rect 7984 24664 7990 24676
rect 8312 24664 8340 24695
rect 8478 24692 8484 24744
rect 8536 24732 8542 24744
rect 9309 24735 9367 24741
rect 9309 24732 9321 24735
rect 8536 24704 9321 24732
rect 8536 24692 8542 24704
rect 9309 24701 9321 24704
rect 9355 24701 9367 24735
rect 10134 24732 10140 24744
rect 10095 24704 10140 24732
rect 9309 24695 9367 24701
rect 10134 24692 10140 24704
rect 10192 24692 10198 24744
rect 10321 24735 10379 24741
rect 10321 24701 10333 24735
rect 10367 24701 10379 24735
rect 10321 24695 10379 24701
rect 7984 24636 8340 24664
rect 10336 24664 10364 24695
rect 10410 24692 10416 24744
rect 10468 24732 10474 24744
rect 10686 24732 10692 24744
rect 10468 24704 10513 24732
rect 10647 24704 10692 24732
rect 10468 24692 10474 24704
rect 10686 24692 10692 24704
rect 10744 24692 10750 24744
rect 12621 24735 12679 24741
rect 12621 24701 12633 24735
rect 12667 24732 12679 24735
rect 12802 24732 12808 24744
rect 12667 24704 12808 24732
rect 12667 24701 12679 24704
rect 12621 24695 12679 24701
rect 12802 24692 12808 24704
rect 12860 24692 12866 24744
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 12912 24704 13461 24732
rect 11146 24664 11152 24676
rect 10336 24636 11152 24664
rect 7984 24624 7990 24636
rect 11146 24624 11152 24636
rect 11204 24664 11210 24676
rect 11514 24664 11520 24676
rect 11204 24636 11520 24664
rect 11204 24624 11210 24636
rect 11514 24624 11520 24636
rect 11572 24624 11578 24676
rect 11790 24624 11796 24676
rect 11848 24664 11854 24676
rect 12912 24664 12940 24704
rect 13449 24701 13461 24704
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 14553 24735 14611 24741
rect 14553 24732 14565 24735
rect 14424 24704 14565 24732
rect 14424 24692 14430 24704
rect 14553 24701 14565 24704
rect 14599 24732 14611 24735
rect 15838 24732 15844 24744
rect 14599 24704 15844 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 15838 24692 15844 24704
rect 15896 24692 15902 24744
rect 16850 24692 16856 24744
rect 16908 24732 16914 24744
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16908 24704 17325 24732
rect 16908 24692 16914 24704
rect 17313 24701 17325 24704
rect 17359 24701 17371 24735
rect 17494 24732 17500 24744
rect 17455 24704 17500 24732
rect 17313 24695 17371 24701
rect 17494 24692 17500 24704
rect 17552 24692 17558 24744
rect 18598 24741 18604 24744
rect 18332 24735 18390 24741
rect 18332 24732 18344 24735
rect 17788 24704 18344 24732
rect 11848 24636 12940 24664
rect 11848 24624 11854 24636
rect 12986 24624 12992 24676
rect 13044 24664 13050 24676
rect 13265 24667 13323 24673
rect 13265 24664 13277 24667
rect 13044 24636 13277 24664
rect 13044 24624 13050 24636
rect 13265 24633 13277 24636
rect 13311 24633 13323 24667
rect 13265 24627 13323 24633
rect 14734 24624 14740 24676
rect 14792 24673 14798 24676
rect 14792 24667 14856 24673
rect 14792 24633 14810 24667
rect 14844 24633 14856 24667
rect 14792 24627 14856 24633
rect 14792 24624 14798 24627
rect 17126 24624 17132 24676
rect 17184 24664 17190 24676
rect 17512 24664 17540 24692
rect 17184 24636 17540 24664
rect 17184 24624 17190 24636
rect 17788 24608 17816 24704
rect 18332 24701 18344 24704
rect 18378 24732 18390 24735
rect 18592 24732 18604 24741
rect 18378 24704 18460 24732
rect 18559 24704 18604 24732
rect 18378 24701 18390 24704
rect 18332 24695 18390 24701
rect 3878 24596 3884 24608
rect 3839 24568 3884 24596
rect 3878 24556 3884 24568
rect 3936 24556 3942 24608
rect 4798 24596 4804 24608
rect 4759 24568 4804 24596
rect 4798 24556 4804 24568
rect 4856 24556 4862 24608
rect 5258 24556 5264 24608
rect 5316 24596 5322 24608
rect 5445 24599 5503 24605
rect 5445 24596 5457 24599
rect 5316 24568 5457 24596
rect 5316 24556 5322 24568
rect 5445 24565 5457 24568
rect 5491 24565 5503 24599
rect 5445 24559 5503 24565
rect 7098 24556 7104 24608
rect 7156 24596 7162 24608
rect 7469 24599 7527 24605
rect 7469 24596 7481 24599
rect 7156 24568 7481 24596
rect 7156 24556 7162 24568
rect 7469 24565 7481 24568
rect 7515 24596 7527 24599
rect 8018 24596 8024 24608
rect 7515 24568 8024 24596
rect 7515 24565 7527 24568
rect 7469 24559 7527 24565
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8570 24596 8576 24608
rect 8352 24568 8576 24596
rect 8352 24556 8358 24568
rect 8570 24556 8576 24568
rect 8628 24556 8634 24608
rect 9493 24599 9551 24605
rect 9493 24565 9505 24599
rect 9539 24596 9551 24599
rect 9674 24596 9680 24608
rect 9539 24568 9680 24596
rect 9539 24565 9551 24568
rect 9493 24559 9551 24565
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 10870 24596 10876 24608
rect 10831 24568 10876 24596
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 12805 24599 12863 24605
rect 12805 24565 12817 24599
rect 12851 24596 12863 24599
rect 13446 24596 13452 24608
rect 12851 24568 13452 24596
rect 12851 24565 12863 24568
rect 12805 24559 12863 24565
rect 13446 24556 13452 24568
rect 13504 24596 13510 24608
rect 13998 24596 14004 24608
rect 13504 24568 14004 24596
rect 13504 24556 13510 24568
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 15933 24599 15991 24605
rect 15933 24596 15945 24599
rect 14700 24568 15945 24596
rect 14700 24556 14706 24568
rect 15933 24565 15945 24568
rect 15979 24565 15991 24599
rect 15933 24559 15991 24565
rect 17770 24556 17776 24608
rect 17828 24556 17834 24608
rect 18432 24596 18460 24704
rect 18592 24695 18604 24704
rect 18598 24692 18604 24695
rect 18656 24692 18662 24744
rect 20349 24735 20407 24741
rect 20349 24701 20361 24735
rect 20395 24732 20407 24735
rect 20806 24732 20812 24744
rect 20395 24704 20812 24732
rect 20395 24701 20407 24704
rect 20349 24695 20407 24701
rect 20806 24692 20812 24704
rect 20864 24732 20870 24744
rect 21450 24732 21456 24744
rect 20864 24704 21456 24732
rect 20864 24692 20870 24704
rect 21450 24692 21456 24704
rect 21508 24692 21514 24744
rect 21637 24735 21695 24741
rect 21637 24701 21649 24735
rect 21683 24732 21695 24735
rect 21726 24732 21732 24744
rect 21683 24704 21732 24732
rect 21683 24701 21695 24704
rect 21637 24695 21695 24701
rect 21726 24692 21732 24704
rect 21784 24692 21790 24744
rect 22741 24735 22799 24741
rect 22741 24732 22753 24735
rect 22066 24704 22753 24732
rect 22066 24676 22094 24704
rect 22741 24701 22753 24704
rect 22787 24701 22799 24735
rect 25498 24732 25504 24744
rect 22741 24695 22799 24701
rect 23308 24704 24808 24732
rect 25459 24704 25504 24732
rect 18690 24624 18696 24676
rect 18748 24664 18754 24676
rect 18748 24636 20944 24664
rect 18748 24624 18754 24636
rect 18782 24596 18788 24608
rect 18432 24568 18788 24596
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 19705 24599 19763 24605
rect 19705 24565 19717 24599
rect 19751 24596 19763 24599
rect 20070 24596 20076 24608
rect 19751 24568 20076 24596
rect 19751 24565 19763 24568
rect 19705 24559 19763 24565
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20916 24596 20944 24636
rect 20990 24624 20996 24676
rect 21048 24664 21054 24676
rect 22002 24664 22008 24676
rect 21048 24636 22008 24664
rect 21048 24624 21054 24636
rect 22002 24624 22008 24636
rect 22060 24636 22094 24676
rect 22060 24624 22066 24636
rect 23308 24596 23336 24704
rect 23382 24624 23388 24676
rect 23440 24664 23446 24676
rect 23937 24667 23995 24673
rect 23937 24664 23949 24667
rect 23440 24636 23949 24664
rect 23440 24624 23446 24636
rect 23937 24633 23949 24636
rect 23983 24664 23995 24667
rect 24578 24664 24584 24676
rect 23983 24636 24584 24664
rect 23983 24633 23995 24636
rect 23937 24627 23995 24633
rect 24578 24624 24584 24636
rect 24636 24624 24642 24676
rect 24673 24667 24731 24673
rect 24673 24633 24685 24667
rect 24719 24633 24731 24667
rect 24780 24664 24808 24704
rect 25498 24692 25504 24704
rect 25556 24692 25562 24744
rect 25774 24741 25780 24744
rect 25768 24732 25780 24741
rect 25735 24704 25780 24732
rect 25768 24695 25780 24704
rect 25774 24692 25780 24695
rect 25832 24692 25838 24744
rect 29012 24741 29040 24772
rect 31294 24760 31300 24812
rect 31352 24800 31358 24812
rect 31573 24803 31631 24809
rect 31573 24800 31585 24803
rect 31352 24772 31585 24800
rect 31352 24760 31358 24772
rect 31573 24769 31585 24772
rect 31619 24769 31631 24803
rect 31573 24763 31631 24769
rect 31662 24760 31668 24812
rect 31720 24800 31726 24812
rect 31720 24772 31892 24800
rect 31720 24760 31726 24772
rect 29362 24741 29368 24744
rect 28997 24735 29055 24741
rect 25884 24704 28028 24732
rect 25884 24664 25912 24704
rect 24780 24636 25912 24664
rect 24673 24627 24731 24633
rect 20916 24568 23336 24596
rect 24394 24556 24400 24608
rect 24452 24596 24458 24608
rect 24688 24596 24716 24627
rect 26142 24624 26148 24676
rect 26200 24664 26206 24676
rect 27893 24667 27951 24673
rect 27893 24664 27905 24667
rect 26200 24636 27905 24664
rect 26200 24624 26206 24636
rect 27893 24633 27905 24636
rect 27939 24633 27951 24667
rect 28000 24664 28028 24704
rect 28997 24701 29009 24735
rect 29043 24732 29055 24735
rect 29089 24735 29147 24741
rect 29089 24732 29101 24735
rect 29043 24704 29101 24732
rect 29043 24701 29055 24704
rect 28997 24695 29055 24701
rect 29089 24701 29101 24704
rect 29135 24701 29147 24735
rect 29356 24732 29368 24741
rect 29323 24704 29368 24732
rect 29089 24695 29147 24701
rect 29356 24695 29368 24704
rect 29362 24692 29368 24695
rect 29420 24692 29426 24744
rect 29730 24692 29736 24744
rect 29788 24732 29794 24744
rect 31864 24741 31892 24772
rect 30929 24735 30987 24741
rect 30929 24732 30941 24735
rect 29788 24704 30941 24732
rect 29788 24692 29794 24704
rect 30929 24701 30941 24704
rect 30975 24701 30987 24735
rect 30929 24695 30987 24701
rect 31757 24735 31815 24741
rect 31757 24701 31769 24735
rect 31803 24701 31815 24735
rect 31757 24695 31815 24701
rect 31849 24735 31907 24741
rect 31849 24701 31861 24735
rect 31895 24701 31907 24735
rect 31849 24695 31907 24701
rect 32125 24735 32183 24741
rect 32125 24701 32137 24735
rect 32171 24732 32183 24735
rect 32582 24732 32588 24744
rect 32171 24704 32588 24732
rect 32171 24701 32183 24704
rect 32125 24695 32183 24701
rect 31772 24664 31800 24695
rect 32582 24692 32588 24704
rect 32640 24692 32646 24744
rect 32692 24732 32720 24840
rect 33318 24828 33324 24880
rect 33376 24868 33382 24880
rect 33704 24877 33732 24908
rect 35986 24896 35992 24908
rect 36044 24896 36050 24948
rect 33689 24871 33747 24877
rect 33689 24868 33701 24871
rect 33376 24840 33701 24868
rect 33376 24828 33382 24840
rect 33689 24837 33701 24840
rect 33735 24837 33747 24871
rect 33689 24831 33747 24837
rect 33962 24800 33968 24812
rect 33428 24772 33968 24800
rect 33428 24741 33456 24772
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 54665 24803 54723 24809
rect 54665 24769 54677 24803
rect 54711 24800 54723 24803
rect 55398 24800 55404 24812
rect 54711 24772 55404 24800
rect 54711 24769 54723 24772
rect 54665 24763 54723 24769
rect 55398 24760 55404 24772
rect 55456 24760 55462 24812
rect 56229 24803 56287 24809
rect 55508 24772 55904 24800
rect 33413 24735 33471 24741
rect 33413 24732 33425 24735
rect 32692 24704 33425 24732
rect 33413 24701 33425 24704
rect 33459 24701 33471 24735
rect 33413 24695 33471 24701
rect 33551 24735 33609 24741
rect 33551 24701 33563 24735
rect 33597 24732 33609 24735
rect 33686 24732 33692 24744
rect 33597 24704 33692 24732
rect 33597 24701 33609 24704
rect 33551 24695 33609 24701
rect 33686 24692 33692 24704
rect 33744 24692 33750 24744
rect 33781 24735 33839 24741
rect 33781 24701 33793 24735
rect 33827 24732 33839 24735
rect 34422 24732 34428 24744
rect 33827 24704 34428 24732
rect 33827 24701 33839 24704
rect 33781 24695 33839 24701
rect 34422 24692 34428 24704
rect 34480 24692 34486 24744
rect 34609 24735 34667 24741
rect 34609 24701 34621 24735
rect 34655 24732 34667 24735
rect 34698 24732 34704 24744
rect 34655 24704 34704 24732
rect 34655 24701 34667 24704
rect 34609 24695 34667 24701
rect 34698 24692 34704 24704
rect 34756 24692 34762 24744
rect 34876 24735 34934 24741
rect 34876 24701 34888 24735
rect 34922 24732 34934 24735
rect 35894 24732 35900 24744
rect 34922 24704 35900 24732
rect 34922 24701 34934 24704
rect 34876 24695 34934 24701
rect 35894 24692 35900 24704
rect 35952 24692 35958 24744
rect 36446 24732 36452 24744
rect 36407 24704 36452 24732
rect 36446 24692 36452 24704
rect 36504 24692 36510 24744
rect 36630 24732 36636 24744
rect 36591 24704 36636 24732
rect 36630 24692 36636 24704
rect 36688 24692 36694 24744
rect 36722 24692 36728 24744
rect 36780 24732 36786 24744
rect 54481 24735 54539 24741
rect 54481 24732 54493 24735
rect 36780 24704 54493 24732
rect 36780 24692 36786 24704
rect 54481 24701 54493 24704
rect 54527 24701 54539 24735
rect 54481 24695 54539 24701
rect 55125 24735 55183 24741
rect 55125 24701 55137 24735
rect 55171 24732 55183 24735
rect 55508 24732 55536 24772
rect 55171 24704 55536 24732
rect 55585 24735 55643 24741
rect 55171 24701 55183 24704
rect 55125 24695 55183 24701
rect 55585 24701 55597 24735
rect 55631 24701 55643 24735
rect 55766 24732 55772 24744
rect 55727 24704 55772 24732
rect 55585 24695 55643 24701
rect 32398 24664 32404 24676
rect 28000 24636 31524 24664
rect 31772 24636 32404 24664
rect 27893 24627 27951 24633
rect 27982 24596 27988 24608
rect 24452 24568 24716 24596
rect 27943 24568 27988 24596
rect 24452 24556 24458 24568
rect 27982 24556 27988 24568
rect 28040 24556 28046 24608
rect 28997 24599 29055 24605
rect 28997 24565 29009 24599
rect 29043 24596 29055 24599
rect 30834 24596 30840 24608
rect 29043 24568 30840 24596
rect 29043 24565 29055 24568
rect 28997 24559 29055 24565
rect 30834 24556 30840 24568
rect 30892 24556 30898 24608
rect 31021 24599 31079 24605
rect 31021 24565 31033 24599
rect 31067 24596 31079 24599
rect 31386 24596 31392 24608
rect 31067 24568 31392 24596
rect 31067 24565 31079 24568
rect 31021 24559 31079 24565
rect 31386 24556 31392 24568
rect 31444 24556 31450 24608
rect 31496 24596 31524 24636
rect 32398 24624 32404 24636
rect 32456 24624 32462 24676
rect 33318 24664 33324 24676
rect 32600 24636 33324 24664
rect 32600 24596 32628 24636
rect 33318 24624 33324 24636
rect 33376 24624 33382 24676
rect 31496 24568 32628 24596
rect 32674 24556 32680 24608
rect 32732 24596 32738 24608
rect 33229 24599 33287 24605
rect 33229 24596 33241 24599
rect 32732 24568 33241 24596
rect 32732 24556 32738 24568
rect 33229 24565 33241 24568
rect 33275 24565 33287 24599
rect 33704 24596 33732 24692
rect 55600 24664 55628 24695
rect 55766 24692 55772 24704
rect 55824 24692 55830 24744
rect 55876 24732 55904 24772
rect 56229 24769 56241 24803
rect 56275 24800 56287 24803
rect 58066 24800 58072 24812
rect 56275 24772 58072 24800
rect 56275 24769 56287 24772
rect 56229 24763 56287 24769
rect 58066 24760 58072 24772
rect 58124 24760 58130 24812
rect 57054 24732 57060 24744
rect 55876 24704 56272 24732
rect 57015 24704 57060 24732
rect 45526 24636 55628 24664
rect 56244 24664 56272 24704
rect 57054 24692 57060 24704
rect 57112 24692 57118 24744
rect 57422 24692 57428 24744
rect 57480 24732 57486 24744
rect 57517 24735 57575 24741
rect 57517 24732 57529 24735
rect 57480 24704 57529 24732
rect 57480 24692 57486 24704
rect 57517 24701 57529 24704
rect 57563 24701 57575 24735
rect 57517 24695 57575 24701
rect 57701 24735 57759 24741
rect 57701 24701 57713 24735
rect 57747 24701 57759 24735
rect 57701 24695 57759 24701
rect 57330 24664 57336 24676
rect 56244 24636 57336 24664
rect 35802 24596 35808 24608
rect 33704 24568 35808 24596
rect 33229 24559 33287 24565
rect 35802 24556 35808 24568
rect 35860 24596 35866 24608
rect 35989 24599 36047 24605
rect 35989 24596 36001 24599
rect 35860 24568 36001 24596
rect 35860 24556 35866 24568
rect 35989 24565 36001 24568
rect 36035 24565 36047 24599
rect 35989 24559 36047 24565
rect 36725 24599 36783 24605
rect 36725 24565 36737 24599
rect 36771 24596 36783 24599
rect 45526 24596 45554 24636
rect 57330 24624 57336 24636
rect 57388 24624 57394 24676
rect 36771 24568 45554 24596
rect 56873 24599 56931 24605
rect 36771 24565 36783 24568
rect 36725 24559 36783 24565
rect 56873 24565 56885 24599
rect 56919 24596 56931 24599
rect 57716 24596 57744 24695
rect 56919 24568 57744 24596
rect 56919 24565 56931 24568
rect 56873 24559 56931 24565
rect 57974 24556 57980 24608
rect 58032 24596 58038 24608
rect 58161 24599 58219 24605
rect 58161 24596 58173 24599
rect 58032 24568 58173 24596
rect 58032 24556 58038 24568
rect 58161 24565 58173 24568
rect 58207 24565 58219 24599
rect 58161 24559 58219 24565
rect 1104 24506 58880 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 50326 24506
rect 50378 24454 50390 24506
rect 50442 24454 50454 24506
rect 50506 24454 50518 24506
rect 50570 24454 58880 24506
rect 1104 24432 58880 24454
rect 5074 24392 5080 24404
rect 1412 24364 5080 24392
rect 1412 24265 1440 24364
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 5626 24392 5632 24404
rect 5587 24364 5632 24392
rect 5626 24352 5632 24364
rect 5684 24352 5690 24404
rect 6086 24392 6092 24404
rect 6047 24364 6092 24392
rect 6086 24352 6092 24364
rect 6144 24352 6150 24404
rect 6362 24352 6368 24404
rect 6420 24392 6426 24404
rect 8478 24392 8484 24404
rect 6420 24364 7604 24392
rect 8439 24364 8484 24392
rect 6420 24352 6426 24364
rect 4516 24327 4574 24333
rect 4516 24293 4528 24327
rect 4562 24324 4574 24327
rect 4798 24324 4804 24336
rect 4562 24296 4804 24324
rect 4562 24293 4574 24296
rect 4516 24287 4574 24293
rect 4798 24284 4804 24296
rect 4856 24284 4862 24336
rect 5258 24284 5264 24336
rect 5316 24324 5322 24336
rect 5316 24296 6684 24324
rect 5316 24284 5322 24296
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24225 1455 24259
rect 1397 24219 1455 24225
rect 2501 24259 2559 24265
rect 2501 24225 2513 24259
rect 2547 24256 2559 24259
rect 3878 24256 3884 24268
rect 2547 24228 3884 24256
rect 2547 24225 2559 24228
rect 2501 24219 2559 24225
rect 3878 24216 3884 24228
rect 3936 24216 3942 24268
rect 6273 24259 6331 24265
rect 6273 24225 6285 24259
rect 6319 24225 6331 24259
rect 6273 24219 6331 24225
rect 1581 24191 1639 24197
rect 1581 24157 1593 24191
rect 1627 24157 1639 24191
rect 2682 24188 2688 24200
rect 2643 24160 2688 24188
rect 1581 24151 1639 24157
rect 1596 24120 1624 24151
rect 2682 24148 2688 24160
rect 2740 24148 2746 24200
rect 4062 24148 4068 24200
rect 4120 24188 4126 24200
rect 4249 24191 4307 24197
rect 4249 24188 4261 24191
rect 4120 24160 4261 24188
rect 4120 24148 4126 24160
rect 4249 24157 4261 24160
rect 4295 24157 4307 24191
rect 6288 24188 6316 24219
rect 6362 24216 6368 24268
rect 6420 24256 6426 24268
rect 6656 24265 6684 24296
rect 7576 24268 7604 24364
rect 8478 24352 8484 24364
rect 8536 24352 8542 24404
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 13633 24395 13691 24401
rect 13633 24392 13645 24395
rect 10468 24364 13645 24392
rect 10468 24352 10474 24364
rect 13633 24361 13645 24364
rect 13679 24361 13691 24395
rect 13633 24355 13691 24361
rect 14458 24352 14464 24404
rect 14516 24392 14522 24404
rect 17221 24395 17279 24401
rect 17221 24392 17233 24395
rect 14516 24364 17233 24392
rect 14516 24352 14522 24364
rect 17221 24361 17233 24364
rect 17267 24361 17279 24395
rect 21729 24395 21787 24401
rect 21729 24392 21741 24395
rect 17221 24355 17279 24361
rect 17696 24364 21741 24392
rect 9582 24324 9588 24336
rect 8404 24296 9588 24324
rect 6641 24259 6699 24265
rect 6420 24228 6465 24256
rect 6420 24216 6426 24228
rect 6641 24225 6653 24259
rect 6687 24225 6699 24259
rect 7466 24256 7472 24268
rect 7427 24228 7472 24256
rect 6641 24219 6699 24225
rect 7466 24216 7472 24228
rect 7524 24216 7530 24268
rect 7558 24216 7564 24268
rect 7616 24256 7622 24268
rect 7837 24259 7895 24265
rect 7616 24228 7661 24256
rect 7616 24216 7622 24228
rect 7837 24225 7849 24259
rect 7883 24256 7895 24259
rect 8018 24256 8024 24268
rect 7883 24228 8024 24256
rect 7883 24225 7895 24228
rect 7837 24219 7895 24225
rect 8018 24216 8024 24228
rect 8076 24216 8082 24268
rect 8294 24216 8300 24268
rect 8352 24256 8358 24268
rect 8404 24265 8432 24296
rect 9582 24284 9588 24296
rect 9640 24284 9646 24336
rect 9760 24327 9818 24333
rect 9760 24293 9772 24327
rect 9806 24324 9818 24327
rect 10870 24324 10876 24336
rect 9806 24296 10876 24324
rect 9806 24293 9818 24296
rect 9760 24287 9818 24293
rect 10870 24284 10876 24296
rect 10928 24284 10934 24336
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 11020 24296 11744 24324
rect 11020 24284 11026 24296
rect 8389 24259 8447 24265
rect 8389 24256 8401 24259
rect 8352 24228 8401 24256
rect 8352 24216 8358 24228
rect 8389 24225 8401 24228
rect 8435 24225 8447 24259
rect 10778 24256 10784 24268
rect 8389 24219 8447 24225
rect 9324 24228 10784 24256
rect 9324 24188 9352 24228
rect 10778 24216 10784 24228
rect 10836 24216 10842 24268
rect 11330 24256 11336 24268
rect 11291 24228 11336 24256
rect 11330 24216 11336 24228
rect 11388 24216 11394 24268
rect 11514 24256 11520 24268
rect 11475 24228 11520 24256
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 11716 24265 11744 24296
rect 12434 24284 12440 24336
rect 12492 24324 12498 24336
rect 16108 24327 16166 24333
rect 12492 24296 14872 24324
rect 12492 24284 12498 24296
rect 14844 24268 14872 24296
rect 16108 24293 16120 24327
rect 16154 24324 16166 24327
rect 16758 24324 16764 24336
rect 16154 24296 16764 24324
rect 16154 24293 16166 24296
rect 16108 24287 16166 24293
rect 16758 24284 16764 24296
rect 16816 24284 16822 24336
rect 11701 24259 11759 24265
rect 11701 24225 11713 24259
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 11885 24259 11943 24265
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 11974 24256 11980 24268
rect 11931 24228 11980 24256
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 11974 24216 11980 24228
rect 12032 24216 12038 24268
rect 12618 24216 12624 24268
rect 12676 24256 12682 24268
rect 12713 24259 12771 24265
rect 12713 24256 12725 24259
rect 12676 24228 12725 24256
rect 12676 24216 12682 24228
rect 12713 24225 12725 24228
rect 12759 24225 12771 24259
rect 12713 24219 12771 24225
rect 13357 24259 13415 24265
rect 13357 24225 13369 24259
rect 13403 24256 13415 24259
rect 14458 24256 14464 24268
rect 13403 24228 14464 24256
rect 13403 24225 13415 24228
rect 13357 24219 13415 24225
rect 14458 24216 14464 24228
rect 14516 24216 14522 24268
rect 14826 24256 14832 24268
rect 14787 24228 14832 24256
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 14918 24216 14924 24268
rect 14976 24256 14982 24268
rect 17696 24256 17724 24364
rect 21729 24361 21741 24364
rect 21775 24361 21787 24395
rect 21729 24355 21787 24361
rect 22833 24395 22891 24401
rect 22833 24361 22845 24395
rect 22879 24392 22891 24395
rect 24394 24392 24400 24404
rect 22879 24364 24400 24392
rect 22879 24361 22891 24364
rect 22833 24355 22891 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 29546 24392 29552 24404
rect 29507 24364 29552 24392
rect 29546 24352 29552 24364
rect 29604 24352 29610 24404
rect 30466 24352 30472 24404
rect 30524 24392 30530 24404
rect 31573 24395 31631 24401
rect 31573 24392 31585 24395
rect 30524 24364 31585 24392
rect 30524 24352 30530 24364
rect 31573 24361 31585 24364
rect 31619 24392 31631 24395
rect 31662 24392 31668 24404
rect 31619 24364 31668 24392
rect 31619 24361 31631 24364
rect 31573 24355 31631 24361
rect 31662 24352 31668 24364
rect 31720 24352 31726 24404
rect 32493 24395 32551 24401
rect 32493 24361 32505 24395
rect 32539 24392 32551 24395
rect 32582 24392 32588 24404
rect 32539 24364 32588 24392
rect 32539 24361 32551 24364
rect 32493 24355 32551 24361
rect 32582 24352 32588 24364
rect 32640 24352 32646 24404
rect 35897 24395 35955 24401
rect 35897 24361 35909 24395
rect 35943 24392 35955 24395
rect 35986 24392 35992 24404
rect 35943 24364 35992 24392
rect 35943 24361 35955 24364
rect 35897 24355 35955 24361
rect 35986 24352 35992 24364
rect 36044 24352 36050 24404
rect 55493 24395 55551 24401
rect 55493 24361 55505 24395
rect 55539 24392 55551 24395
rect 55766 24392 55772 24404
rect 55539 24364 55772 24392
rect 55539 24361 55551 24364
rect 55493 24355 55551 24361
rect 55766 24352 55772 24364
rect 55824 24352 55830 24404
rect 19058 24324 19064 24336
rect 19019 24296 19064 24324
rect 19058 24284 19064 24296
rect 19116 24284 19122 24336
rect 20901 24327 20959 24333
rect 20901 24324 20913 24327
rect 19720 24296 20913 24324
rect 14976 24228 17724 24256
rect 17865 24259 17923 24265
rect 14976 24216 14982 24228
rect 17865 24225 17877 24259
rect 17911 24225 17923 24259
rect 17865 24219 17923 24225
rect 6288 24160 9352 24188
rect 9493 24191 9551 24197
rect 4249 24151 4307 24157
rect 9493 24157 9505 24191
rect 9539 24157 9551 24191
rect 11606 24188 11612 24200
rect 11567 24160 11612 24188
rect 9493 24151 9551 24157
rect 3050 24120 3056 24132
rect 1596 24092 3056 24120
rect 3050 24080 3056 24092
rect 3108 24080 3114 24132
rect 7745 24123 7803 24129
rect 7745 24120 7757 24123
rect 6564 24092 7757 24120
rect 6564 24064 6592 24092
rect 7745 24089 7757 24092
rect 7791 24120 7803 24123
rect 7926 24120 7932 24132
rect 7791 24092 7932 24120
rect 7791 24089 7803 24092
rect 7745 24083 7803 24089
rect 7926 24080 7932 24092
rect 7984 24080 7990 24132
rect 8662 24080 8668 24132
rect 8720 24120 8726 24132
rect 9508 24120 9536 24151
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 12069 24191 12127 24197
rect 12069 24157 12081 24191
rect 12115 24188 12127 24191
rect 12342 24188 12348 24200
rect 12115 24160 12348 24188
rect 12115 24157 12127 24160
rect 12069 24151 12127 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 13633 24191 13691 24197
rect 13633 24188 13645 24191
rect 12912 24160 13645 24188
rect 12912 24129 12940 24160
rect 13633 24157 13645 24160
rect 13679 24188 13691 24191
rect 14182 24188 14188 24200
rect 13679 24160 14188 24188
rect 13679 24157 13691 24160
rect 13633 24151 13691 24157
rect 14182 24148 14188 24160
rect 14240 24148 14246 24200
rect 15838 24188 15844 24200
rect 15751 24160 15844 24188
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 17880 24188 17908 24219
rect 17954 24216 17960 24268
rect 18012 24256 18018 24268
rect 18012 24228 18057 24256
rect 18012 24216 18018 24228
rect 18230 24216 18236 24268
rect 18288 24256 18294 24268
rect 18325 24259 18383 24265
rect 18325 24256 18337 24259
rect 18288 24228 18337 24256
rect 18288 24216 18294 24228
rect 18325 24225 18337 24228
rect 18371 24225 18383 24259
rect 18325 24219 18383 24225
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 18877 24259 18935 24265
rect 18877 24256 18889 24259
rect 18656 24228 18889 24256
rect 18656 24216 18662 24228
rect 18877 24225 18889 24228
rect 18923 24256 18935 24259
rect 19720 24256 19748 24296
rect 20901 24293 20913 24296
rect 20947 24324 20959 24327
rect 21174 24324 21180 24336
rect 20947 24296 21180 24324
rect 20947 24293 20959 24296
rect 20901 24287 20959 24293
rect 21174 24284 21180 24296
rect 21232 24324 21238 24336
rect 21818 24324 21824 24336
rect 21232 24296 21824 24324
rect 21232 24284 21238 24296
rect 21818 24284 21824 24296
rect 21876 24284 21882 24336
rect 21910 24284 21916 24336
rect 21968 24324 21974 24336
rect 22005 24327 22063 24333
rect 22005 24324 22017 24327
rect 21968 24296 22017 24324
rect 21968 24284 21974 24296
rect 22005 24293 22017 24296
rect 22051 24324 22063 24327
rect 23477 24327 23535 24333
rect 23477 24324 23489 24327
rect 22051 24296 23489 24324
rect 22051 24293 22063 24296
rect 22005 24287 22063 24293
rect 23477 24293 23489 24296
rect 23523 24324 23535 24327
rect 26605 24327 26663 24333
rect 26605 24324 26617 24327
rect 23523 24296 26617 24324
rect 23523 24293 23535 24296
rect 23477 24287 23535 24293
rect 26605 24293 26617 24296
rect 26651 24293 26663 24327
rect 26605 24287 26663 24293
rect 26789 24327 26847 24333
rect 26789 24293 26801 24327
rect 26835 24324 26847 24327
rect 29086 24324 29092 24336
rect 26835 24296 29092 24324
rect 26835 24293 26847 24296
rect 26789 24287 26847 24293
rect 29086 24284 29092 24296
rect 29144 24284 29150 24336
rect 57974 24324 57980 24336
rect 57935 24296 57980 24324
rect 57974 24284 57980 24296
rect 58032 24284 58038 24336
rect 58158 24324 58164 24336
rect 58119 24296 58164 24324
rect 58158 24284 58164 24296
rect 58216 24284 58222 24336
rect 20622 24256 20628 24268
rect 18923 24228 19748 24256
rect 20180 24228 20628 24256
rect 18923 24225 18935 24228
rect 18877 24219 18935 24225
rect 18046 24188 18052 24200
rect 17788 24160 17908 24188
rect 18007 24160 18052 24188
rect 8720 24092 9536 24120
rect 12897 24123 12955 24129
rect 8720 24080 8726 24092
rect 12897 24089 12909 24123
rect 12943 24089 12955 24123
rect 12897 24083 12955 24089
rect 1854 24052 1860 24064
rect 1815 24024 1860 24052
rect 1854 24012 1860 24024
rect 1912 24012 1918 24064
rect 1946 24012 1952 24064
rect 2004 24052 2010 24064
rect 2869 24055 2927 24061
rect 2869 24052 2881 24055
rect 2004 24024 2881 24052
rect 2004 24012 2010 24024
rect 2869 24021 2881 24024
rect 2915 24021 2927 24055
rect 6546 24052 6552 24064
rect 6507 24024 6552 24052
rect 2869 24015 2927 24021
rect 6546 24012 6552 24024
rect 6604 24012 6610 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7285 24055 7343 24061
rect 7285 24052 7297 24055
rect 6972 24024 7297 24052
rect 6972 24012 6978 24024
rect 7285 24021 7297 24024
rect 7331 24021 7343 24055
rect 7285 24015 7343 24021
rect 8386 24012 8392 24064
rect 8444 24052 8450 24064
rect 10686 24052 10692 24064
rect 8444 24024 10692 24052
rect 8444 24012 8450 24024
rect 10686 24012 10692 24024
rect 10744 24052 10750 24064
rect 10873 24055 10931 24061
rect 10873 24052 10885 24055
rect 10744 24024 10885 24052
rect 10744 24012 10750 24024
rect 10873 24021 10885 24024
rect 10919 24021 10931 24055
rect 13446 24052 13452 24064
rect 13407 24024 13452 24052
rect 10873 24015 10931 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 13538 24012 13544 24064
rect 13596 24052 13602 24064
rect 15013 24055 15071 24061
rect 15013 24052 15025 24055
rect 13596 24024 15025 24052
rect 13596 24012 13602 24024
rect 15013 24021 15025 24024
rect 15059 24021 15071 24055
rect 15856 24052 15884 24148
rect 17586 24120 17592 24132
rect 16776 24092 17592 24120
rect 16776 24052 16804 24092
rect 17586 24080 17592 24092
rect 17644 24080 17650 24132
rect 15856 24024 16804 24052
rect 15013 24015 15071 24021
rect 17310 24012 17316 24064
rect 17368 24052 17374 24064
rect 17681 24055 17739 24061
rect 17681 24052 17693 24055
rect 17368 24024 17693 24052
rect 17368 24012 17374 24024
rect 17681 24021 17693 24024
rect 17727 24021 17739 24055
rect 17788 24052 17816 24160
rect 18046 24148 18052 24160
rect 18104 24148 18110 24200
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 20180 24188 20208 24228
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 22646 24216 22652 24268
rect 22704 24256 22710 24268
rect 22741 24259 22799 24265
rect 22741 24256 22753 24259
rect 22704 24228 22753 24256
rect 22704 24216 22710 24228
rect 22741 24225 22753 24228
rect 22787 24225 22799 24259
rect 22741 24219 22799 24225
rect 22830 24216 22836 24268
rect 22888 24256 22894 24268
rect 24121 24259 24179 24265
rect 24121 24256 24133 24259
rect 22888 24228 24133 24256
rect 22888 24216 22894 24228
rect 24121 24225 24133 24228
rect 24167 24225 24179 24259
rect 24121 24219 24179 24225
rect 25406 24216 25412 24268
rect 25464 24256 25470 24268
rect 25501 24259 25559 24265
rect 25501 24256 25513 24259
rect 25464 24228 25513 24256
rect 25464 24216 25470 24228
rect 25501 24225 25513 24228
rect 25547 24225 25559 24259
rect 25682 24256 25688 24268
rect 25643 24228 25688 24256
rect 25501 24219 25559 24225
rect 25682 24216 25688 24228
rect 25740 24216 25746 24268
rect 25777 24259 25835 24265
rect 25777 24225 25789 24259
rect 25823 24225 25835 24259
rect 25777 24219 25835 24225
rect 25869 24259 25927 24265
rect 25869 24225 25881 24259
rect 25915 24256 25927 24259
rect 27338 24256 27344 24268
rect 25915 24228 27344 24256
rect 25915 24225 25927 24228
rect 25869 24219 25927 24225
rect 20346 24188 20352 24200
rect 18187 24160 20208 24188
rect 20307 24160 20352 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 21729 24191 21787 24197
rect 21729 24157 21741 24191
rect 21775 24188 21787 24191
rect 25792 24188 25820 24219
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 30653 24259 30711 24265
rect 30653 24225 30665 24259
rect 30699 24256 30711 24259
rect 30742 24256 30748 24268
rect 30699 24228 30748 24256
rect 30699 24225 30711 24228
rect 30653 24219 30711 24225
rect 30742 24216 30748 24228
rect 30800 24216 30806 24268
rect 31297 24259 31355 24265
rect 31297 24225 31309 24259
rect 31343 24225 31355 24259
rect 31297 24219 31355 24225
rect 31389 24259 31447 24265
rect 31389 24225 31401 24259
rect 31435 24256 31447 24259
rect 32030 24256 32036 24268
rect 31435 24228 32036 24256
rect 31435 24225 31447 24228
rect 31389 24219 31447 24225
rect 26510 24188 26516 24200
rect 21775 24160 24431 24188
rect 25792 24160 26516 24188
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 21910 24120 21916 24132
rect 18012 24092 21916 24120
rect 18012 24080 18018 24092
rect 21910 24080 21916 24092
rect 21968 24080 21974 24132
rect 22002 24080 22008 24132
rect 22060 24120 22066 24132
rect 24305 24123 24363 24129
rect 24305 24120 24317 24123
rect 22060 24092 24317 24120
rect 22060 24080 22066 24092
rect 24305 24089 24317 24092
rect 24351 24089 24363 24123
rect 24403 24120 24431 24160
rect 26510 24148 26516 24160
rect 26568 24148 26574 24200
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24188 27951 24191
rect 28350 24188 28356 24200
rect 27939 24160 28356 24188
rect 27939 24157 27951 24160
rect 27893 24151 27951 24157
rect 28350 24148 28356 24160
rect 28408 24148 28414 24200
rect 28902 24188 28908 24200
rect 28863 24160 28908 24188
rect 28902 24148 28908 24160
rect 28960 24148 28966 24200
rect 30282 24148 30288 24200
rect 30340 24188 30346 24200
rect 30469 24191 30527 24197
rect 30469 24188 30481 24191
rect 30340 24160 30481 24188
rect 30340 24148 30346 24160
rect 30469 24157 30481 24160
rect 30515 24157 30527 24191
rect 30469 24151 30527 24157
rect 30834 24148 30840 24200
rect 30892 24188 30898 24200
rect 31312 24188 31340 24219
rect 32030 24216 32036 24228
rect 32088 24216 32094 24268
rect 32398 24256 32404 24268
rect 32311 24228 32404 24256
rect 32398 24216 32404 24228
rect 32456 24256 32462 24268
rect 32674 24256 32680 24268
rect 32456 24228 32680 24256
rect 32456 24216 32462 24228
rect 32674 24216 32680 24228
rect 32732 24216 32738 24268
rect 33134 24216 33140 24268
rect 33192 24256 33198 24268
rect 33301 24259 33359 24265
rect 33301 24256 33313 24259
rect 33192 24228 33313 24256
rect 33192 24216 33198 24228
rect 33301 24225 33313 24228
rect 33347 24225 33359 24259
rect 35802 24256 35808 24268
rect 35763 24228 35808 24256
rect 33301 24219 33359 24225
rect 35802 24216 35808 24228
rect 35860 24216 35866 24268
rect 55674 24256 55680 24268
rect 55635 24228 55680 24256
rect 55674 24216 55680 24228
rect 55732 24216 55738 24268
rect 57422 24256 57428 24268
rect 57383 24228 57428 24256
rect 57422 24216 57428 24228
rect 57480 24216 57486 24268
rect 31478 24188 31484 24200
rect 30892 24160 31156 24188
rect 31312 24160 31484 24188
rect 30892 24148 30898 24160
rect 31018 24120 31024 24132
rect 24403 24092 31024 24120
rect 24305 24083 24363 24089
rect 31018 24080 31024 24092
rect 31076 24080 31082 24132
rect 31128 24120 31156 24160
rect 31478 24148 31484 24160
rect 31536 24148 31542 24200
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24188 31631 24191
rect 31754 24188 31760 24200
rect 31619 24160 31760 24188
rect 31619 24157 31631 24160
rect 31573 24151 31631 24157
rect 31754 24148 31760 24160
rect 31812 24148 31818 24200
rect 33045 24191 33103 24197
rect 33045 24157 33057 24191
rect 33091 24157 33103 24191
rect 33045 24151 33103 24157
rect 33060 24120 33088 24151
rect 34698 24120 34704 24132
rect 31128 24092 33088 24120
rect 20162 24052 20168 24064
rect 17788 24024 20168 24052
rect 17681 24015 17739 24021
rect 20162 24012 20168 24024
rect 20220 24052 20226 24064
rect 20530 24052 20536 24064
rect 20220 24024 20536 24052
rect 20220 24012 20226 24024
rect 20530 24012 20536 24024
rect 20588 24012 20594 24064
rect 20898 24012 20904 24064
rect 20956 24052 20962 24064
rect 22097 24055 22155 24061
rect 22097 24052 22109 24055
rect 20956 24024 22109 24052
rect 20956 24012 20962 24024
rect 22097 24021 22109 24024
rect 22143 24021 22155 24055
rect 22097 24015 22155 24021
rect 23106 24012 23112 24064
rect 23164 24052 23170 24064
rect 23566 24052 23572 24064
rect 23164 24024 23572 24052
rect 23164 24012 23170 24024
rect 23566 24012 23572 24024
rect 23624 24012 23630 24064
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 26053 24055 26111 24061
rect 26053 24052 26065 24055
rect 25188 24024 26065 24052
rect 25188 24012 25194 24024
rect 26053 24021 26065 24024
rect 26099 24021 26111 24055
rect 28442 24052 28448 24064
rect 28403 24024 28448 24052
rect 26053 24015 26111 24021
rect 28442 24012 28448 24024
rect 28500 24012 28506 24064
rect 30834 24052 30840 24064
rect 30795 24024 30840 24052
rect 30834 24012 30840 24024
rect 30892 24012 30898 24064
rect 33060 24052 33088 24092
rect 33980 24092 34704 24120
rect 33980 24052 34008 24092
rect 34698 24080 34704 24092
rect 34756 24080 34762 24132
rect 33060 24024 34008 24052
rect 34146 24012 34152 24064
rect 34204 24052 34210 24064
rect 34425 24055 34483 24061
rect 34425 24052 34437 24055
rect 34204 24024 34437 24052
rect 34204 24012 34210 24024
rect 34425 24021 34437 24024
rect 34471 24021 34483 24055
rect 34425 24015 34483 24021
rect 1104 23962 58880 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 58880 23962
rect 1104 23888 58880 23910
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 6546 23848 6552 23860
rect 5859 23820 6552 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 6822 23808 6828 23860
rect 6880 23848 6886 23860
rect 8662 23848 8668 23860
rect 6880 23820 8668 23848
rect 6880 23808 6886 23820
rect 8662 23808 8668 23820
rect 8720 23808 8726 23860
rect 8846 23848 8852 23860
rect 8807 23820 8852 23848
rect 8846 23808 8852 23820
rect 8904 23848 8910 23860
rect 9122 23848 9128 23860
rect 8904 23820 9128 23848
rect 8904 23808 8910 23820
rect 9122 23808 9128 23820
rect 9180 23808 9186 23860
rect 9769 23851 9827 23857
rect 9769 23817 9781 23851
rect 9815 23848 9827 23851
rect 9858 23848 9864 23860
rect 9815 23820 9864 23848
rect 9815 23817 9827 23820
rect 9769 23811 9827 23817
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 11974 23848 11980 23860
rect 10428 23820 11980 23848
rect 2958 23740 2964 23792
rect 3016 23780 3022 23792
rect 3605 23783 3663 23789
rect 3605 23780 3617 23783
rect 3016 23752 3617 23780
rect 3016 23740 3022 23752
rect 3605 23749 3617 23752
rect 3651 23749 3663 23783
rect 3605 23743 3663 23749
rect 5552 23752 6888 23780
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23712 2191 23715
rect 2866 23712 2872 23724
rect 2179 23684 2872 23712
rect 2179 23681 2191 23684
rect 2133 23675 2191 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 3237 23715 3295 23721
rect 3237 23681 3249 23715
rect 3283 23712 3295 23715
rect 4614 23712 4620 23724
rect 3283 23684 4620 23712
rect 3283 23681 3295 23684
rect 3237 23675 3295 23681
rect 4614 23672 4620 23684
rect 4672 23672 4678 23724
rect 5353 23715 5411 23721
rect 5353 23712 5365 23715
rect 4724 23684 5365 23712
rect 1489 23647 1547 23653
rect 1489 23613 1501 23647
rect 1535 23644 1547 23647
rect 1946 23644 1952 23656
rect 1535 23616 1952 23644
rect 1535 23613 1547 23616
rect 1489 23607 1547 23613
rect 1946 23604 1952 23616
rect 2004 23604 2010 23656
rect 2317 23647 2375 23653
rect 2317 23613 2329 23647
rect 2363 23644 2375 23647
rect 3421 23647 3479 23653
rect 2363 23616 2774 23644
rect 2363 23613 2375 23616
rect 2317 23607 2375 23613
rect 2746 23576 2774 23616
rect 3421 23613 3433 23647
rect 3467 23644 3479 23647
rect 4430 23644 4436 23656
rect 3467 23616 4436 23644
rect 3467 23613 3479 23616
rect 3421 23607 3479 23613
rect 4430 23604 4436 23616
rect 4488 23604 4494 23656
rect 4724 23653 4752 23684
rect 5353 23681 5365 23684
rect 5399 23681 5411 23715
rect 5353 23675 5411 23681
rect 4709 23647 4767 23653
rect 4709 23613 4721 23647
rect 4755 23613 4767 23647
rect 4709 23607 4767 23613
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23644 4951 23647
rect 4982 23644 4988 23656
rect 4939 23616 4988 23644
rect 4939 23613 4951 23616
rect 4893 23607 4951 23613
rect 4982 23604 4988 23616
rect 5040 23604 5046 23656
rect 5552 23653 5580 23752
rect 5994 23712 6000 23724
rect 5644 23684 6000 23712
rect 5644 23653 5672 23684
rect 5994 23672 6000 23684
rect 6052 23712 6058 23724
rect 6362 23712 6368 23724
rect 6052 23684 6368 23712
rect 6052 23672 6058 23684
rect 6362 23672 6368 23684
rect 6420 23672 6426 23724
rect 6860 23712 6888 23752
rect 8202 23740 8208 23792
rect 8260 23780 8266 23792
rect 10428 23780 10456 23820
rect 11974 23808 11980 23820
rect 12032 23848 12038 23860
rect 13449 23851 13507 23857
rect 13449 23848 13461 23851
rect 12032 23820 13461 23848
rect 12032 23808 12038 23820
rect 13449 23817 13461 23820
rect 13495 23817 13507 23851
rect 13998 23848 14004 23860
rect 13959 23820 14004 23848
rect 13449 23811 13507 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14826 23808 14832 23860
rect 14884 23848 14890 23860
rect 17034 23848 17040 23860
rect 14884 23820 17040 23848
rect 14884 23808 14890 23820
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 20346 23848 20352 23860
rect 20307 23820 20352 23848
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 23382 23848 23388 23860
rect 20456 23820 23388 23848
rect 8260 23752 10456 23780
rect 10873 23783 10931 23789
rect 8260 23740 8266 23752
rect 10873 23749 10885 23783
rect 10919 23780 10931 23783
rect 11238 23780 11244 23792
rect 10919 23752 11244 23780
rect 10919 23749 10931 23752
rect 10873 23743 10931 23749
rect 11238 23740 11244 23752
rect 11296 23780 11302 23792
rect 11882 23780 11888 23792
rect 11296 23752 11888 23780
rect 11296 23740 11302 23752
rect 11882 23740 11888 23752
rect 11940 23740 11946 23792
rect 20456 23780 20484 23820
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 23566 23808 23572 23860
rect 23624 23848 23630 23860
rect 26142 23848 26148 23860
rect 23624 23820 26148 23848
rect 23624 23808 23630 23820
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 29181 23851 29239 23857
rect 29181 23817 29193 23851
rect 29227 23848 29239 23851
rect 29362 23848 29368 23860
rect 29227 23820 29368 23848
rect 29227 23817 29239 23820
rect 29181 23811 29239 23817
rect 29362 23808 29368 23820
rect 29420 23848 29426 23860
rect 29730 23848 29736 23860
rect 29420 23820 29736 23848
rect 29420 23808 29426 23820
rect 29730 23808 29736 23820
rect 29788 23808 29794 23860
rect 30469 23851 30527 23857
rect 30469 23817 30481 23851
rect 30515 23848 30527 23851
rect 30558 23848 30564 23860
rect 30515 23820 30564 23848
rect 30515 23817 30527 23820
rect 30469 23811 30527 23817
rect 30558 23808 30564 23820
rect 30616 23808 30622 23860
rect 32033 23851 32091 23857
rect 32033 23817 32045 23851
rect 32079 23848 32091 23851
rect 32214 23848 32220 23860
rect 32079 23820 32220 23848
rect 32079 23817 32091 23820
rect 32033 23811 32091 23817
rect 32214 23808 32220 23820
rect 32272 23808 32278 23860
rect 33045 23851 33103 23857
rect 33045 23817 33057 23851
rect 33091 23848 33103 23851
rect 33134 23848 33140 23860
rect 33091 23820 33140 23848
rect 33091 23817 33103 23820
rect 33045 23811 33103 23817
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 36630 23848 36636 23860
rect 34164 23820 36636 23848
rect 14016 23752 20484 23780
rect 11974 23712 11980 23724
rect 6860 23684 6960 23712
rect 5537 23647 5595 23653
rect 5537 23613 5549 23647
rect 5583 23613 5595 23647
rect 5537 23607 5595 23613
rect 5629 23647 5687 23653
rect 5629 23613 5641 23647
rect 5675 23613 5687 23647
rect 5902 23644 5908 23656
rect 5863 23616 5908 23644
rect 5629 23607 5687 23613
rect 5902 23604 5908 23616
rect 5960 23604 5966 23656
rect 6822 23644 6828 23656
rect 6783 23616 6828 23644
rect 6822 23604 6828 23616
rect 6880 23604 6886 23656
rect 6932 23644 6960 23684
rect 8404 23684 11980 23712
rect 8404 23644 8432 23684
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 14016 23712 14044 23752
rect 21542 23740 21548 23792
rect 21600 23780 21606 23792
rect 23290 23780 23296 23792
rect 21600 23752 23296 23780
rect 21600 23740 21606 23752
rect 23290 23740 23296 23752
rect 23348 23740 23354 23792
rect 25041 23783 25099 23789
rect 25041 23749 25053 23783
rect 25087 23780 25099 23783
rect 26510 23780 26516 23792
rect 25087 23752 26516 23780
rect 25087 23749 25099 23752
rect 25041 23743 25099 23749
rect 26510 23740 26516 23752
rect 26568 23740 26574 23792
rect 30926 23740 30932 23792
rect 30984 23780 30990 23792
rect 34164 23780 34192 23820
rect 36630 23808 36636 23820
rect 36688 23808 36694 23860
rect 56042 23848 56048 23860
rect 56003 23820 56048 23848
rect 56042 23808 56048 23820
rect 56100 23808 56106 23860
rect 30984 23752 34192 23780
rect 34241 23783 34299 23789
rect 30984 23740 30990 23752
rect 14182 23712 14188 23724
rect 13924 23684 14044 23712
rect 14143 23684 14188 23712
rect 6932 23616 8432 23644
rect 8478 23604 8484 23656
rect 8536 23644 8542 23656
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8536 23616 8769 23644
rect 8536 23604 8542 23616
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 8757 23607 8815 23613
rect 9585 23647 9643 23653
rect 9585 23613 9597 23647
rect 9631 23644 9643 23647
rect 9674 23644 9680 23656
rect 9631 23616 9680 23644
rect 9631 23613 9643 23616
rect 9585 23607 9643 23613
rect 9674 23604 9680 23616
rect 9732 23644 9738 23656
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 9732 23616 10609 23644
rect 9732 23604 9738 23616
rect 10597 23613 10609 23616
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12342 23653 12348 23656
rect 12336 23644 12348 23653
rect 12124 23616 12169 23644
rect 12303 23616 12348 23644
rect 12124 23604 12130 23616
rect 12336 23607 12348 23616
rect 12342 23604 12348 23607
rect 12400 23604 12406 23656
rect 13924 23653 13952 23684
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 15194 23712 15200 23724
rect 14752 23684 15056 23712
rect 15155 23684 15200 23712
rect 13910 23647 13968 23653
rect 13910 23613 13922 23647
rect 13956 23613 13968 23647
rect 14274 23644 14280 23656
rect 13910 23607 13968 23613
rect 14016 23616 14280 23644
rect 4522 23576 4528 23588
rect 2746 23548 4528 23576
rect 4522 23536 4528 23548
rect 4580 23536 4586 23588
rect 7006 23536 7012 23588
rect 7064 23585 7070 23588
rect 7064 23579 7128 23585
rect 7064 23545 7082 23579
rect 7116 23545 7128 23579
rect 7064 23539 7128 23545
rect 7064 23536 7070 23539
rect 7558 23536 7564 23588
rect 7616 23576 7622 23588
rect 7616 23548 9904 23576
rect 7616 23536 7622 23548
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 4798 23508 4804 23520
rect 2832 23480 2877 23508
rect 4759 23480 4804 23508
rect 2832 23468 2838 23480
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 7834 23468 7840 23520
rect 7892 23508 7898 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 7892 23480 8217 23508
rect 7892 23468 7898 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 9876 23508 9904 23548
rect 14016 23508 14044 23616
rect 14274 23604 14280 23616
rect 14332 23644 14338 23656
rect 14752 23644 14780 23684
rect 14918 23644 14924 23656
rect 14332 23616 14780 23644
rect 14879 23616 14924 23644
rect 14332 23604 14338 23616
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 15028 23653 15056 23684
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 16301 23715 16359 23721
rect 16301 23681 16313 23715
rect 16347 23712 16359 23715
rect 18969 23715 19027 23721
rect 18969 23712 18981 23715
rect 16347 23684 18981 23712
rect 16347 23681 16359 23684
rect 16301 23675 16359 23681
rect 18969 23681 18981 23684
rect 19015 23681 19027 23715
rect 18969 23675 19027 23681
rect 19613 23715 19671 23721
rect 19613 23681 19625 23715
rect 19659 23712 19671 23715
rect 26602 23712 26608 23724
rect 19659 23684 23796 23712
rect 19659 23681 19671 23684
rect 19613 23675 19671 23681
rect 15013 23647 15071 23653
rect 15013 23613 15025 23647
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 15289 23647 15347 23653
rect 15289 23613 15301 23647
rect 15335 23644 15347 23647
rect 15654 23644 15660 23656
rect 15335 23616 15660 23644
rect 15335 23613 15347 23616
rect 15289 23607 15347 23613
rect 15654 23604 15660 23616
rect 15712 23604 15718 23656
rect 16206 23644 16212 23656
rect 16167 23616 16212 23644
rect 16206 23604 16212 23616
rect 16264 23604 16270 23656
rect 16390 23644 16396 23656
rect 16351 23616 16396 23644
rect 16390 23604 16396 23616
rect 16448 23604 16454 23656
rect 17862 23644 17868 23656
rect 17823 23616 17868 23644
rect 17862 23604 17868 23616
rect 17920 23604 17926 23656
rect 20070 23644 20076 23656
rect 20031 23616 20076 23644
rect 20070 23604 20076 23616
rect 20128 23604 20134 23656
rect 22186 23644 22192 23656
rect 21376 23616 22192 23644
rect 14458 23536 14464 23588
rect 14516 23576 14522 23588
rect 14516 23548 18644 23576
rect 14516 23536 14522 23548
rect 14182 23508 14188 23520
rect 9876 23480 14044 23508
rect 14143 23480 14188 23508
rect 8205 23471 8263 23477
rect 14182 23468 14188 23480
rect 14240 23468 14246 23520
rect 14737 23511 14795 23517
rect 14737 23477 14749 23511
rect 14783 23508 14795 23511
rect 15378 23508 15384 23520
rect 14783 23480 15384 23508
rect 14783 23477 14795 23480
rect 14737 23471 14795 23477
rect 15378 23468 15384 23480
rect 15436 23468 15442 23520
rect 18506 23508 18512 23520
rect 18467 23480 18512 23508
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 18616 23508 18644 23548
rect 19426 23536 19432 23588
rect 19484 23576 19490 23588
rect 20257 23579 20315 23585
rect 20257 23576 20269 23579
rect 19484 23548 20269 23576
rect 19484 23536 19490 23548
rect 20257 23545 20269 23548
rect 20303 23545 20315 23579
rect 20257 23539 20315 23545
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 21269 23579 21327 23585
rect 21269 23576 21281 23579
rect 20404 23548 21281 23576
rect 20404 23536 20410 23548
rect 21269 23545 21281 23548
rect 21315 23545 21327 23579
rect 21269 23539 21327 23545
rect 21376 23508 21404 23616
rect 22186 23604 22192 23616
rect 22244 23604 22250 23656
rect 22278 23604 22284 23656
rect 22336 23644 22342 23656
rect 22830 23644 22836 23656
rect 22336 23616 22836 23644
rect 22336 23604 22342 23616
rect 22830 23604 22836 23616
rect 22888 23604 22894 23656
rect 23290 23604 23296 23656
rect 23348 23644 23354 23656
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23348 23616 23673 23644
rect 23348 23604 23354 23616
rect 23661 23613 23673 23616
rect 23707 23613 23719 23647
rect 23768 23644 23796 23684
rect 25332 23684 26608 23712
rect 23917 23647 23975 23653
rect 23917 23644 23929 23647
rect 23768 23616 23929 23644
rect 23661 23607 23719 23613
rect 23917 23613 23929 23616
rect 23963 23613 23975 23647
rect 23917 23607 23975 23613
rect 24210 23604 24216 23656
rect 24268 23644 24274 23656
rect 25332 23644 25360 23684
rect 26602 23672 26608 23684
rect 26660 23672 26666 23724
rect 27798 23712 27804 23724
rect 27759 23684 27804 23712
rect 27798 23672 27804 23684
rect 27856 23672 27862 23724
rect 30374 23672 30380 23724
rect 30432 23712 30438 23724
rect 30432 23684 31432 23712
rect 30432 23672 30438 23684
rect 31404 23656 31432 23684
rect 25498 23644 25504 23656
rect 24268 23616 25360 23644
rect 25459 23616 25504 23644
rect 24268 23604 24274 23616
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 26697 23647 26755 23653
rect 26697 23613 26709 23647
rect 26743 23644 26755 23647
rect 26878 23644 26884 23656
rect 26743 23616 26884 23644
rect 26743 23613 26755 23616
rect 26697 23607 26755 23613
rect 26878 23604 26884 23616
rect 26936 23604 26942 23656
rect 28068 23647 28126 23653
rect 28068 23613 28080 23647
rect 28114 23644 28126 23647
rect 28442 23644 28448 23656
rect 28114 23616 28448 23644
rect 28114 23613 28126 23616
rect 28068 23607 28126 23613
rect 28442 23604 28448 23616
rect 28500 23604 28506 23656
rect 30101 23647 30159 23653
rect 30101 23613 30113 23647
rect 30147 23644 30159 23647
rect 30742 23644 30748 23656
rect 30147 23616 30748 23644
rect 30147 23613 30159 23616
rect 30101 23607 30159 23613
rect 30742 23604 30748 23616
rect 30800 23604 30806 23656
rect 31018 23604 31024 23656
rect 31076 23644 31082 23656
rect 31113 23647 31171 23653
rect 31113 23644 31125 23647
rect 31076 23616 31125 23644
rect 31076 23604 31082 23616
rect 31113 23613 31125 23616
rect 31159 23613 31171 23647
rect 31113 23607 31171 23613
rect 31205 23647 31263 23653
rect 31205 23613 31217 23647
rect 31251 23613 31263 23647
rect 31386 23644 31392 23656
rect 31347 23616 31392 23644
rect 31205 23607 31263 23613
rect 21450 23536 21456 23588
rect 21508 23576 21514 23588
rect 22646 23576 22652 23588
rect 21508 23548 22652 23576
rect 21508 23536 21514 23548
rect 22646 23536 22652 23548
rect 22704 23536 22710 23588
rect 25314 23576 25320 23588
rect 23584 23548 25320 23576
rect 21634 23508 21640 23520
rect 18616 23480 21404 23508
rect 21595 23480 21640 23508
rect 21634 23468 21640 23480
rect 21692 23468 21698 23520
rect 21818 23468 21824 23520
rect 21876 23508 21882 23520
rect 23584 23508 23612 23548
rect 25314 23536 25320 23548
rect 25372 23536 25378 23588
rect 30006 23576 30012 23588
rect 25884 23548 30012 23576
rect 21876 23480 23612 23508
rect 21876 23468 21882 23480
rect 25038 23468 25044 23520
rect 25096 23508 25102 23520
rect 25884 23508 25912 23548
rect 30006 23536 30012 23548
rect 30064 23536 30070 23588
rect 30282 23576 30288 23588
rect 30243 23548 30288 23576
rect 30282 23536 30288 23548
rect 30340 23536 30346 23588
rect 25096 23480 25912 23508
rect 25096 23468 25102 23480
rect 25958 23468 25964 23520
rect 26016 23508 26022 23520
rect 26145 23511 26203 23517
rect 26145 23508 26157 23511
rect 26016 23480 26157 23508
rect 26016 23468 26022 23480
rect 26145 23477 26157 23480
rect 26191 23477 26203 23511
rect 26145 23471 26203 23477
rect 26789 23511 26847 23517
rect 26789 23477 26801 23511
rect 26835 23508 26847 23511
rect 27154 23508 27160 23520
rect 26835 23480 27160 23508
rect 26835 23477 26847 23480
rect 26789 23471 26847 23477
rect 27154 23468 27160 23480
rect 27212 23468 27218 23520
rect 30929 23511 30987 23517
rect 30929 23477 30941 23511
rect 30975 23508 30987 23511
rect 31018 23508 31024 23520
rect 30975 23480 31024 23508
rect 30975 23477 30987 23480
rect 30929 23471 30987 23477
rect 31018 23468 31024 23480
rect 31076 23468 31082 23520
rect 31128 23508 31156 23607
rect 31220 23576 31248 23607
rect 31386 23604 31392 23616
rect 31444 23604 31450 23656
rect 31496 23653 31524 23752
rect 34241 23749 34253 23783
rect 34287 23780 34299 23783
rect 34422 23780 34428 23792
rect 34287 23752 34428 23780
rect 34287 23749 34299 23752
rect 34241 23743 34299 23749
rect 34422 23740 34428 23752
rect 34480 23740 34486 23792
rect 58158 23780 58164 23792
rect 58119 23752 58164 23780
rect 58158 23740 58164 23752
rect 58216 23740 58222 23792
rect 34698 23672 34704 23724
rect 34756 23712 34762 23724
rect 34793 23715 34851 23721
rect 34793 23712 34805 23715
rect 34756 23684 34805 23712
rect 34756 23672 34762 23684
rect 34793 23681 34805 23684
rect 34839 23681 34851 23715
rect 34793 23675 34851 23681
rect 31481 23647 31539 23653
rect 31481 23613 31493 23647
rect 31527 23613 31539 23647
rect 31938 23644 31944 23656
rect 31899 23616 31944 23644
rect 31481 23607 31539 23613
rect 31938 23604 31944 23616
rect 31996 23604 32002 23656
rect 33226 23604 33232 23656
rect 33284 23644 33290 23656
rect 33321 23647 33379 23653
rect 33321 23644 33333 23647
rect 33284 23616 33333 23644
rect 33284 23604 33290 23616
rect 33321 23613 33333 23616
rect 33367 23613 33379 23647
rect 33321 23607 33379 23613
rect 33413 23647 33471 23653
rect 33413 23613 33425 23647
rect 33459 23613 33471 23647
rect 33413 23607 33471 23613
rect 31570 23576 31576 23588
rect 31220 23548 31576 23576
rect 31570 23536 31576 23548
rect 31628 23536 31634 23588
rect 33428 23576 33456 23607
rect 33502 23604 33508 23656
rect 33560 23644 33566 23656
rect 33686 23644 33692 23656
rect 33560 23616 33605 23644
rect 33647 23616 33692 23644
rect 33560 23604 33566 23616
rect 33686 23604 33692 23616
rect 33744 23604 33750 23656
rect 33962 23604 33968 23656
rect 34020 23644 34026 23656
rect 34149 23647 34207 23653
rect 34149 23644 34161 23647
rect 34020 23616 34161 23644
rect 34020 23604 34026 23616
rect 34149 23613 34161 23616
rect 34195 23613 34207 23647
rect 34149 23607 34207 23613
rect 34238 23604 34244 23656
rect 34296 23644 34302 23656
rect 34716 23644 34744 23672
rect 34296 23616 34744 23644
rect 34296 23604 34302 23616
rect 35342 23604 35348 23656
rect 35400 23644 35406 23656
rect 36633 23647 36691 23653
rect 36633 23644 36645 23647
rect 35400 23616 36645 23644
rect 35400 23604 35406 23616
rect 36633 23613 36645 23616
rect 36679 23613 36691 23647
rect 55401 23647 55459 23653
rect 55401 23644 55413 23647
rect 36633 23607 36691 23613
rect 55232 23616 55413 23644
rect 34054 23576 34060 23588
rect 33428 23548 34060 23576
rect 34054 23536 34060 23548
rect 34112 23536 34118 23588
rect 35060 23579 35118 23585
rect 35060 23545 35072 23579
rect 35106 23576 35118 23579
rect 35986 23576 35992 23588
rect 35106 23548 35992 23576
rect 35106 23545 35118 23548
rect 35060 23539 35118 23545
rect 35986 23536 35992 23548
rect 36044 23536 36050 23588
rect 55232 23520 55260 23616
rect 55401 23613 55413 23616
rect 55447 23613 55459 23647
rect 55582 23644 55588 23656
rect 55543 23616 55588 23644
rect 55401 23607 55459 23613
rect 55582 23604 55588 23616
rect 55640 23604 55646 23656
rect 56502 23604 56508 23656
rect 56560 23644 56566 23656
rect 56597 23647 56655 23653
rect 56597 23644 56609 23647
rect 56560 23616 56609 23644
rect 56560 23604 56566 23616
rect 56597 23613 56609 23616
rect 56643 23613 56655 23647
rect 56597 23607 56655 23613
rect 57241 23647 57299 23653
rect 57241 23613 57253 23647
rect 57287 23644 57299 23647
rect 57330 23644 57336 23656
rect 57287 23616 57336 23644
rect 57287 23613 57299 23616
rect 57241 23607 57299 23613
rect 57330 23604 57336 23616
rect 57388 23604 57394 23656
rect 57977 23579 58035 23585
rect 57977 23545 57989 23579
rect 58023 23576 58035 23579
rect 58066 23576 58072 23588
rect 58023 23548 58072 23576
rect 58023 23545 58035 23548
rect 57977 23539 58035 23545
rect 58066 23536 58072 23548
rect 58124 23536 58130 23588
rect 31386 23508 31392 23520
rect 31128 23480 31392 23508
rect 31386 23468 31392 23480
rect 31444 23468 31450 23520
rect 31938 23468 31944 23520
rect 31996 23508 32002 23520
rect 34514 23508 34520 23520
rect 31996 23480 34520 23508
rect 31996 23468 32002 23480
rect 34514 23468 34520 23480
rect 34572 23468 34578 23520
rect 36170 23508 36176 23520
rect 36131 23480 36176 23508
rect 36170 23468 36176 23480
rect 36228 23468 36234 23520
rect 36722 23508 36728 23520
rect 36683 23480 36728 23508
rect 36722 23468 36728 23480
rect 36780 23468 36786 23520
rect 55214 23468 55220 23520
rect 55272 23508 55278 23520
rect 55272 23480 55317 23508
rect 55272 23468 55278 23480
rect 1104 23418 58880 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 50326 23418
rect 50378 23366 50390 23418
rect 50442 23366 50454 23418
rect 50506 23366 50518 23418
rect 50570 23366 58880 23418
rect 1104 23344 58880 23366
rect 3142 23304 3148 23316
rect 3103 23276 3148 23304
rect 3142 23264 3148 23276
rect 3200 23264 3206 23316
rect 7006 23304 7012 23316
rect 6967 23276 7012 23304
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 10321 23307 10379 23313
rect 10321 23304 10333 23307
rect 10192 23276 10333 23304
rect 10192 23264 10198 23276
rect 10321 23273 10333 23276
rect 10367 23273 10379 23307
rect 10321 23267 10379 23273
rect 10962 23264 10968 23316
rect 11020 23264 11026 23316
rect 11146 23264 11152 23316
rect 11204 23304 11210 23316
rect 12345 23307 12403 23313
rect 12345 23304 12357 23307
rect 11204 23276 12357 23304
rect 11204 23264 11210 23276
rect 12345 23273 12357 23276
rect 12391 23273 12403 23307
rect 12345 23267 12403 23273
rect 13173 23307 13231 23313
rect 13173 23273 13185 23307
rect 13219 23304 13231 23307
rect 54294 23304 54300 23316
rect 13219 23276 54300 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 54294 23264 54300 23276
rect 54352 23264 54358 23316
rect 54665 23307 54723 23313
rect 54665 23273 54677 23307
rect 54711 23304 54723 23307
rect 55582 23304 55588 23316
rect 54711 23276 55588 23304
rect 54711 23273 54723 23276
rect 54665 23267 54723 23273
rect 55582 23264 55588 23276
rect 55640 23264 55646 23316
rect 1854 23236 1860 23248
rect 1815 23208 1860 23236
rect 1854 23196 1860 23208
rect 1912 23196 1918 23248
rect 4798 23196 4804 23248
rect 4856 23245 4862 23248
rect 4856 23239 4920 23245
rect 4856 23205 4874 23239
rect 4908 23205 4920 23239
rect 10980 23236 11008 23264
rect 10980 23208 11376 23236
rect 4856 23199 4920 23205
rect 4856 23196 4862 23199
rect 2501 23171 2559 23177
rect 2501 23137 2513 23171
rect 2547 23168 2559 23171
rect 2590 23168 2596 23180
rect 2547 23140 2596 23168
rect 2547 23137 2559 23140
rect 2501 23131 2559 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 3329 23171 3387 23177
rect 3329 23137 3341 23171
rect 3375 23168 3387 23171
rect 3418 23168 3424 23180
rect 3375 23140 3424 23168
rect 3375 23137 3387 23140
rect 3329 23131 3387 23137
rect 2685 23035 2743 23041
rect 2685 23001 2697 23035
rect 2731 23032 2743 23035
rect 3344 23032 3372 23131
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 4062 23128 4068 23180
rect 4120 23168 4126 23180
rect 4617 23171 4675 23177
rect 4617 23168 4629 23171
rect 4120 23140 4629 23168
rect 4120 23128 4126 23140
rect 4617 23137 4629 23140
rect 4663 23168 4675 23171
rect 6914 23168 6920 23180
rect 4663 23140 6776 23168
rect 6875 23140 6920 23168
rect 4663 23137 4675 23140
rect 4617 23131 4675 23137
rect 6748 23100 6776 23140
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7101 23171 7159 23177
rect 7101 23137 7113 23171
rect 7147 23168 7159 23171
rect 7190 23168 7196 23180
rect 7147 23140 7196 23168
rect 7147 23137 7159 23140
rect 7101 23131 7159 23137
rect 7190 23128 7196 23140
rect 7248 23128 7254 23180
rect 7834 23168 7840 23180
rect 7795 23140 7840 23168
rect 7834 23128 7840 23140
rect 7892 23128 7898 23180
rect 9493 23171 9551 23177
rect 9493 23137 9505 23171
rect 9539 23168 9551 23171
rect 9674 23168 9680 23180
rect 9539 23140 9680 23168
rect 9539 23137 9551 23140
rect 9493 23131 9551 23137
rect 9674 23128 9680 23140
rect 9732 23168 9738 23180
rect 10137 23171 10195 23177
rect 10137 23168 10149 23171
rect 9732 23140 10149 23168
rect 9732 23128 9738 23140
rect 10137 23137 10149 23140
rect 10183 23137 10195 23171
rect 10137 23131 10195 23137
rect 10318 23128 10324 23180
rect 10376 23168 10382 23180
rect 10965 23171 11023 23177
rect 10965 23168 10977 23171
rect 10376 23140 10977 23168
rect 10376 23128 10382 23140
rect 10965 23137 10977 23140
rect 11011 23137 11023 23171
rect 11146 23168 11152 23180
rect 11107 23140 11152 23168
rect 10965 23131 11023 23137
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 11348 23177 11376 23208
rect 12066 23196 12072 23248
rect 12124 23236 12130 23248
rect 14550 23236 14556 23248
rect 12124 23208 14556 23236
rect 12124 23196 12130 23208
rect 14550 23196 14556 23208
rect 14608 23236 14614 23248
rect 14608 23208 14780 23236
rect 14608 23196 14614 23208
rect 11333 23171 11391 23177
rect 11333 23137 11345 23171
rect 11379 23137 11391 23171
rect 11514 23168 11520 23180
rect 11475 23140 11520 23168
rect 11333 23131 11391 23137
rect 11514 23128 11520 23140
rect 11572 23128 11578 23180
rect 11790 23128 11796 23180
rect 11848 23168 11854 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11848 23140 12173 23168
rect 11848 23128 11854 23140
rect 12161 23137 12173 23140
rect 12207 23168 12219 23171
rect 12342 23168 12348 23180
rect 12207 23140 12348 23168
rect 12207 23137 12219 23140
rect 12161 23131 12219 23137
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 14752 23177 14780 23208
rect 16206 23196 16212 23248
rect 16264 23236 16270 23248
rect 17948 23239 18006 23245
rect 16264 23208 17908 23236
rect 16264 23196 16270 23208
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 14737 23171 14795 23177
rect 13311 23140 14688 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 7926 23100 7932 23112
rect 6748 23072 7932 23100
rect 7926 23060 7932 23072
rect 7984 23060 7990 23112
rect 2731 23004 3372 23032
rect 9677 23035 9735 23041
rect 2731 23001 2743 23004
rect 2685 22995 2743 23001
rect 9677 23001 9689 23035
rect 9723 23032 9735 23035
rect 10336 23032 10364 23128
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23069 11299 23103
rect 11241 23063 11299 23069
rect 9723 23004 10364 23032
rect 11256 23032 11284 23063
rect 11698 23060 11704 23112
rect 11756 23100 11762 23112
rect 13173 23103 13231 23109
rect 13173 23100 13185 23103
rect 11756 23072 13185 23100
rect 11756 23060 11762 23072
rect 13173 23069 13185 23072
rect 13219 23069 13231 23103
rect 13173 23063 13231 23069
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 14090 23100 14096 23112
rect 13587 23072 14096 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 14090 23060 14096 23072
rect 14148 23060 14154 23112
rect 13449 23035 13507 23041
rect 13449 23032 13461 23035
rect 11256 23004 13461 23032
rect 9723 23001 9735 23004
rect 9677 22995 9735 23001
rect 13449 23001 13461 23004
rect 13495 23001 13507 23035
rect 13449 22995 13507 23001
rect 1946 22964 1952 22976
rect 1907 22936 1952 22964
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 5718 22924 5724 22976
rect 5776 22964 5782 22976
rect 5997 22967 6055 22973
rect 5997 22964 6009 22967
rect 5776 22936 6009 22964
rect 5776 22924 5782 22936
rect 5997 22933 6009 22936
rect 6043 22933 6055 22967
rect 5997 22927 6055 22933
rect 7929 22967 7987 22973
rect 7929 22933 7941 22967
rect 7975 22964 7987 22967
rect 8018 22964 8024 22976
rect 7975 22936 8024 22964
rect 7975 22933 7987 22936
rect 7929 22927 7987 22933
rect 8018 22924 8024 22936
rect 8076 22924 8082 22976
rect 8570 22924 8576 22976
rect 8628 22964 8634 22976
rect 11238 22964 11244 22976
rect 8628 22936 11244 22964
rect 8628 22924 8634 22936
rect 11238 22924 11244 22936
rect 11296 22924 11302 22976
rect 11701 22967 11759 22973
rect 11701 22933 11713 22967
rect 11747 22964 11759 22967
rect 12158 22964 12164 22976
rect 11747 22936 12164 22964
rect 11747 22933 11759 22936
rect 11701 22927 11759 22933
rect 12158 22924 12164 22936
rect 12216 22924 12222 22976
rect 13357 22967 13415 22973
rect 13357 22933 13369 22967
rect 13403 22964 13415 22967
rect 13998 22964 14004 22976
rect 13403 22936 14004 22964
rect 13403 22933 13415 22936
rect 13357 22927 13415 22933
rect 13998 22924 14004 22936
rect 14056 22924 14062 22976
rect 14660 22964 14688 23140
rect 14737 23137 14749 23171
rect 14783 23137 14795 23171
rect 14737 23131 14795 23137
rect 15004 23171 15062 23177
rect 15004 23137 15016 23171
rect 15050 23168 15062 23171
rect 15286 23168 15292 23180
rect 15050 23140 15292 23168
rect 15050 23137 15062 23140
rect 15004 23131 15062 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 17034 23168 17040 23180
rect 16995 23140 17040 23168
rect 17034 23128 17040 23140
rect 17092 23128 17098 23180
rect 17681 23171 17739 23177
rect 17681 23137 17693 23171
rect 17727 23168 17739 23171
rect 17770 23168 17776 23180
rect 17727 23140 17776 23168
rect 17727 23137 17739 23140
rect 17681 23131 17739 23137
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 17880 23168 17908 23208
rect 17948 23205 17960 23239
rect 17994 23236 18006 23239
rect 18506 23236 18512 23248
rect 17994 23208 18512 23236
rect 17994 23205 18006 23208
rect 17948 23199 18006 23205
rect 18506 23196 18512 23208
rect 18564 23196 18570 23248
rect 19168 23208 22692 23236
rect 19168 23168 19196 23208
rect 20070 23168 20076 23180
rect 17880 23140 19196 23168
rect 19260 23140 20076 23168
rect 19260 23100 19288 23140
rect 20070 23128 20076 23140
rect 20128 23128 20134 23180
rect 20162 23128 20168 23180
rect 20220 23168 20226 23180
rect 20625 23171 20683 23177
rect 20220 23140 20265 23168
rect 20220 23128 20226 23140
rect 20625 23137 20637 23171
rect 20671 23168 20683 23171
rect 20714 23168 20720 23180
rect 20671 23140 20720 23168
rect 20671 23137 20683 23140
rect 20625 23131 20683 23137
rect 20714 23128 20720 23140
rect 20772 23128 20778 23180
rect 21726 23128 21732 23180
rect 21784 23168 21790 23180
rect 21893 23171 21951 23177
rect 21893 23168 21905 23171
rect 21784 23140 21905 23168
rect 21784 23128 21790 23140
rect 21893 23137 21905 23140
rect 21939 23137 21951 23171
rect 21893 23131 21951 23137
rect 18708 23072 19288 23100
rect 15672 23004 17264 23032
rect 15672 22964 15700 23004
rect 16114 22964 16120 22976
rect 14660 22936 15700 22964
rect 16075 22936 16120 22964
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 17034 22924 17040 22976
rect 17092 22964 17098 22976
rect 17129 22967 17187 22973
rect 17129 22964 17141 22967
rect 17092 22936 17141 22964
rect 17092 22924 17098 22936
rect 17129 22933 17141 22936
rect 17175 22933 17187 22967
rect 17236 22964 17264 23004
rect 18708 22964 18736 23072
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20349 23103 20407 23109
rect 20349 23100 20361 23103
rect 20036 23072 20361 23100
rect 20036 23060 20042 23072
rect 20349 23069 20361 23072
rect 20395 23069 20407 23103
rect 20349 23063 20407 23069
rect 20438 23060 20444 23112
rect 20496 23109 20502 23112
rect 20496 23103 20516 23109
rect 20504 23069 20516 23103
rect 20496 23063 20516 23069
rect 20496 23060 20502 23063
rect 21542 23060 21548 23112
rect 21600 23100 21606 23112
rect 21637 23103 21695 23109
rect 21637 23100 21649 23103
rect 21600 23072 21649 23100
rect 21600 23060 21606 23072
rect 21637 23069 21649 23072
rect 21683 23069 21695 23103
rect 22664 23100 22692 23208
rect 24854 23196 24860 23248
rect 24912 23236 24918 23248
rect 25317 23239 25375 23245
rect 25317 23236 25329 23239
rect 24912 23208 25329 23236
rect 24912 23196 24918 23208
rect 25317 23205 25329 23208
rect 25363 23205 25375 23239
rect 25317 23199 25375 23205
rect 25501 23239 25559 23245
rect 25501 23205 25513 23239
rect 25547 23236 25559 23239
rect 25866 23236 25872 23248
rect 25547 23208 25872 23236
rect 25547 23205 25559 23208
rect 25501 23199 25559 23205
rect 25866 23196 25872 23208
rect 25924 23196 25930 23248
rect 26228 23239 26286 23245
rect 26228 23205 26240 23239
rect 26274 23236 26286 23239
rect 26326 23236 26332 23248
rect 26274 23208 26332 23236
rect 26274 23205 26286 23208
rect 26228 23199 26286 23205
rect 26326 23196 26332 23208
rect 26384 23196 26390 23248
rect 30834 23236 30840 23248
rect 26436 23208 29040 23236
rect 22830 23128 22836 23180
rect 22888 23168 22894 23180
rect 23842 23168 23848 23180
rect 22888 23140 23848 23168
rect 22888 23128 22894 23140
rect 23842 23128 23848 23140
rect 23900 23128 23906 23180
rect 24121 23171 24179 23177
rect 24121 23137 24133 23171
rect 24167 23168 24179 23171
rect 24210 23168 24216 23180
rect 24167 23140 24216 23168
rect 24167 23137 24179 23140
rect 24121 23131 24179 23137
rect 24210 23128 24216 23140
rect 24268 23128 24274 23180
rect 24302 23128 24308 23180
rect 24360 23168 24366 23180
rect 26436 23168 26464 23208
rect 24360 23140 24405 23168
rect 25516 23140 26464 23168
rect 24360 23128 24366 23140
rect 23661 23103 23719 23109
rect 23661 23100 23673 23103
rect 22664 23072 23673 23100
rect 21637 23063 21695 23069
rect 23661 23069 23673 23072
rect 23707 23069 23719 23103
rect 24026 23100 24032 23112
rect 23987 23072 24032 23100
rect 23661 23063 23719 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 18782 22992 18788 23044
rect 18840 23032 18846 23044
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 18840 23004 20269 23032
rect 18840 22992 18846 23004
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 23937 23035 23995 23041
rect 23937 23001 23949 23035
rect 23983 23032 23995 23035
rect 25516 23032 25544 23140
rect 26510 23128 26516 23180
rect 26568 23168 26574 23180
rect 27801 23171 27859 23177
rect 27801 23168 27813 23171
rect 26568 23140 27813 23168
rect 26568 23128 26574 23140
rect 27801 23137 27813 23140
rect 27847 23137 27859 23171
rect 27801 23131 27859 23137
rect 28810 23128 28816 23180
rect 28868 23168 28874 23180
rect 28905 23171 28963 23177
rect 28905 23168 28917 23171
rect 28868 23140 28917 23168
rect 28868 23128 28874 23140
rect 28905 23137 28917 23140
rect 28951 23137 28963 23171
rect 28905 23131 28963 23137
rect 25590 23060 25596 23112
rect 25648 23100 25654 23112
rect 25961 23103 26019 23109
rect 25961 23100 25973 23103
rect 25648 23072 25973 23100
rect 25648 23060 25654 23072
rect 25961 23069 25973 23072
rect 26007 23069 26019 23103
rect 29012 23100 29040 23208
rect 29104 23208 30840 23236
rect 29104 23177 29132 23208
rect 30834 23196 30840 23208
rect 30892 23196 30898 23248
rect 31754 23196 31760 23248
rect 31812 23236 31818 23248
rect 32585 23239 32643 23245
rect 31812 23208 31857 23236
rect 31812 23196 31818 23208
rect 32585 23205 32597 23239
rect 32631 23236 32643 23239
rect 36170 23236 36176 23248
rect 32631 23208 33364 23236
rect 32631 23205 32643 23208
rect 32585 23199 32643 23205
rect 29089 23171 29147 23177
rect 29089 23137 29101 23171
rect 29135 23137 29147 23171
rect 29089 23131 29147 23137
rect 29365 23171 29423 23177
rect 29365 23137 29377 23171
rect 29411 23168 29423 23171
rect 29454 23168 29460 23180
rect 29411 23140 29460 23168
rect 29411 23137 29423 23140
rect 29365 23131 29423 23137
rect 29454 23128 29460 23140
rect 29512 23128 29518 23180
rect 31018 23168 31024 23180
rect 30979 23140 31024 23168
rect 31018 23128 31024 23140
rect 31076 23128 31082 23180
rect 31202 23168 31208 23180
rect 31163 23140 31208 23168
rect 31202 23128 31208 23140
rect 31260 23128 31266 23180
rect 31570 23168 31576 23180
rect 31531 23140 31576 23168
rect 31570 23128 31576 23140
rect 31628 23128 31634 23180
rect 32214 23168 32220 23180
rect 32175 23140 32220 23168
rect 32214 23128 32220 23140
rect 32272 23128 32278 23180
rect 32398 23177 32404 23180
rect 32365 23171 32404 23177
rect 32365 23137 32377 23171
rect 32365 23131 32404 23137
rect 32398 23128 32404 23131
rect 32456 23128 32462 23180
rect 33336 23177 33364 23208
rect 34256 23208 36176 23236
rect 32493 23171 32551 23177
rect 32493 23137 32505 23171
rect 32539 23137 32551 23171
rect 32493 23131 32551 23137
rect 32723 23171 32781 23177
rect 32723 23137 32735 23171
rect 32769 23168 32781 23171
rect 33321 23171 33379 23177
rect 32769 23140 33272 23168
rect 32769 23137 32781 23140
rect 32723 23131 32781 23137
rect 29181 23103 29239 23109
rect 29012 23072 29132 23100
rect 25961 23063 26019 23069
rect 27338 23032 27344 23044
rect 23983 23004 25544 23032
rect 27299 23004 27344 23032
rect 23983 23001 23995 23004
rect 23937 22995 23995 23001
rect 27338 22992 27344 23004
rect 27396 22992 27402 23044
rect 28997 23035 29055 23041
rect 28997 23001 29009 23035
rect 29043 23001 29055 23035
rect 29104 23032 29132 23072
rect 29181 23069 29193 23103
rect 29227 23100 29239 23103
rect 29270 23100 29276 23112
rect 29227 23072 29276 23100
rect 29227 23069 29239 23072
rect 29181 23063 29239 23069
rect 29270 23060 29276 23072
rect 29328 23100 29334 23112
rect 30374 23100 30380 23112
rect 29328 23072 30380 23100
rect 29328 23060 29334 23072
rect 30374 23060 30380 23072
rect 30432 23060 30438 23112
rect 31294 23100 31300 23112
rect 31255 23072 31300 23100
rect 31294 23060 31300 23072
rect 31352 23060 31358 23112
rect 31386 23060 31392 23112
rect 31444 23100 31450 23112
rect 31444 23072 31489 23100
rect 31444 23060 31450 23072
rect 31754 23060 31760 23112
rect 31812 23100 31818 23112
rect 32508 23100 32536 23131
rect 31812 23072 32536 23100
rect 33244 23100 33272 23140
rect 33321 23137 33333 23171
rect 33367 23168 33379 23171
rect 33965 23171 34023 23177
rect 33965 23168 33977 23171
rect 33367 23140 33977 23168
rect 33367 23137 33379 23140
rect 33321 23131 33379 23137
rect 33965 23137 33977 23140
rect 34011 23137 34023 23171
rect 34146 23168 34152 23180
rect 34107 23140 34152 23168
rect 33965 23131 34023 23137
rect 34146 23128 34152 23140
rect 34204 23128 34210 23180
rect 34256 23177 34284 23208
rect 34241 23171 34299 23177
rect 34241 23137 34253 23171
rect 34287 23137 34299 23171
rect 34514 23168 34520 23180
rect 34475 23140 34520 23168
rect 34241 23131 34299 23137
rect 34514 23128 34520 23140
rect 34572 23128 34578 23180
rect 36004 23177 36032 23208
rect 36170 23196 36176 23208
rect 36228 23196 36234 23248
rect 35989 23171 36047 23177
rect 35989 23137 36001 23171
rect 36035 23137 36047 23171
rect 35989 23131 36047 23137
rect 36081 23171 36139 23177
rect 36081 23137 36093 23171
rect 36127 23168 36139 23171
rect 36538 23168 36544 23180
rect 36127 23140 36544 23168
rect 36127 23137 36139 23140
rect 36081 23131 36139 23137
rect 36538 23128 36544 23140
rect 36596 23128 36602 23180
rect 54849 23171 54907 23177
rect 54849 23137 54861 23171
rect 54895 23168 54907 23171
rect 55309 23171 55367 23177
rect 54895 23140 55214 23168
rect 54895 23137 54907 23140
rect 54849 23131 54907 23137
rect 36722 23100 36728 23112
rect 33244 23072 36728 23100
rect 31812 23060 31818 23072
rect 29546 23032 29552 23044
rect 29104 23004 29552 23032
rect 28997 22995 29055 23001
rect 19058 22964 19064 22976
rect 17236 22936 18736 22964
rect 19019 22936 19064 22964
rect 17129 22927 17187 22933
rect 19058 22924 19064 22936
rect 19116 22924 19122 22976
rect 19150 22924 19156 22976
rect 19208 22964 19214 22976
rect 19981 22967 20039 22973
rect 19981 22964 19993 22967
rect 19208 22936 19993 22964
rect 19208 22924 19214 22936
rect 19981 22933 19993 22936
rect 20027 22933 20039 22967
rect 19981 22927 20039 22933
rect 21358 22924 21364 22976
rect 21416 22964 21422 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 21416 22936 23029 22964
rect 21416 22924 21422 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 23017 22927 23075 22933
rect 24210 22924 24216 22976
rect 24268 22964 24274 22976
rect 25682 22964 25688 22976
rect 24268 22936 25688 22964
rect 24268 22924 24274 22936
rect 25682 22924 25688 22936
rect 25740 22964 25746 22976
rect 26878 22964 26884 22976
rect 25740 22936 26884 22964
rect 25740 22924 25746 22936
rect 26878 22924 26884 22936
rect 26936 22964 26942 22976
rect 27893 22967 27951 22973
rect 27893 22964 27905 22967
rect 26936 22936 27905 22964
rect 26936 22924 26942 22936
rect 27893 22933 27905 22936
rect 27939 22933 27951 22967
rect 27893 22927 27951 22933
rect 28258 22924 28264 22976
rect 28316 22964 28322 22976
rect 28721 22967 28779 22973
rect 28721 22964 28733 22967
rect 28316 22936 28733 22964
rect 28316 22924 28322 22936
rect 28721 22933 28733 22936
rect 28767 22933 28779 22967
rect 29012 22964 29040 22995
rect 29546 22992 29552 23004
rect 29604 22992 29610 23044
rect 32306 22964 32312 22976
rect 29012 22936 32312 22964
rect 28721 22927 28779 22933
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 32508 22964 32536 23072
rect 36722 23060 36728 23072
rect 36780 23060 36786 23112
rect 32861 23035 32919 23041
rect 32861 23001 32873 23035
rect 32907 23032 32919 23035
rect 33686 23032 33692 23044
rect 32907 23004 33692 23032
rect 32907 23001 32919 23004
rect 32861 22995 32919 23001
rect 33686 22992 33692 23004
rect 33744 22992 33750 23044
rect 34422 23032 34428 23044
rect 34335 23004 34428 23032
rect 34422 22992 34428 23004
rect 34480 23032 34486 23044
rect 36538 23032 36544 23044
rect 34480 23004 36544 23032
rect 34480 22992 34486 23004
rect 36538 22992 36544 23004
rect 36596 22992 36602 23044
rect 55186 23032 55214 23140
rect 55309 23137 55321 23171
rect 55355 23168 55367 23171
rect 55398 23168 55404 23180
rect 55355 23140 55404 23168
rect 55355 23137 55367 23140
rect 55309 23131 55367 23137
rect 55398 23128 55404 23140
rect 55456 23128 55462 23180
rect 57974 23168 57980 23180
rect 57935 23140 57980 23168
rect 57974 23128 57980 23140
rect 58032 23128 58038 23180
rect 55493 23035 55551 23041
rect 55493 23032 55505 23035
rect 55186 23004 55505 23032
rect 55493 23001 55505 23004
rect 55539 23032 55551 23035
rect 55674 23032 55680 23044
rect 55539 23004 55680 23032
rect 55539 23001 55551 23004
rect 55493 22995 55551 23001
rect 55674 22992 55680 23004
rect 55732 22992 55738 23044
rect 58158 23032 58164 23044
rect 58119 23004 58164 23032
rect 58158 22992 58164 23004
rect 58216 22992 58222 23044
rect 33413 22967 33471 22973
rect 33413 22964 33425 22967
rect 32508 22936 33425 22964
rect 33413 22933 33425 22936
rect 33459 22933 33471 22967
rect 33413 22927 33471 22933
rect 57425 22967 57483 22973
rect 57425 22933 57437 22967
rect 57471 22964 57483 22967
rect 57514 22964 57520 22976
rect 57471 22936 57520 22964
rect 57471 22933 57483 22936
rect 57425 22927 57483 22933
rect 57514 22924 57520 22936
rect 57572 22924 57578 22976
rect 1104 22874 58880 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 58880 22874
rect 1104 22800 58880 22822
rect 6914 22760 6920 22772
rect 2746 22732 6920 22760
rect 2130 22692 2136 22704
rect 2091 22664 2136 22692
rect 2130 22652 2136 22664
rect 2188 22652 2194 22704
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2746 22624 2774 22732
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 14182 22760 14188 22772
rect 10612 22732 14188 22760
rect 2866 22652 2872 22704
rect 2924 22692 2930 22704
rect 3697 22695 3755 22701
rect 3697 22692 3709 22695
rect 2924 22664 3709 22692
rect 2924 22652 2930 22664
rect 3697 22661 3709 22664
rect 3743 22661 3755 22695
rect 9861 22695 9919 22701
rect 9861 22692 9873 22695
rect 3697 22655 3755 22661
rect 9646 22664 9873 22692
rect 1811 22596 2774 22624
rect 3329 22627 3387 22633
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 3329 22593 3341 22627
rect 3375 22624 3387 22627
rect 4890 22624 4896 22636
rect 3375 22596 4896 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 8478 22624 8484 22636
rect 8439 22596 8484 22624
rect 8478 22584 8484 22596
rect 8536 22584 8542 22636
rect 1949 22559 2007 22565
rect 1949 22525 1961 22559
rect 1995 22556 2007 22559
rect 2038 22556 2044 22568
rect 1995 22528 2044 22556
rect 1995 22525 2007 22528
rect 1949 22519 2007 22525
rect 2038 22516 2044 22528
rect 2096 22516 2102 22568
rect 3510 22556 3516 22568
rect 3471 22528 3516 22556
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 5718 22556 5724 22568
rect 5679 22528 5724 22556
rect 5718 22516 5724 22528
rect 5776 22516 5782 22568
rect 7466 22556 7472 22568
rect 7427 22528 7472 22556
rect 7466 22516 7472 22528
rect 7524 22516 7530 22568
rect 7561 22559 7619 22565
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 9646 22556 9674 22664
rect 9861 22661 9873 22664
rect 9907 22692 9919 22695
rect 10502 22692 10508 22704
rect 9907 22664 10508 22692
rect 9907 22661 9919 22664
rect 9861 22655 9919 22661
rect 10502 22652 10508 22664
rect 10560 22652 10566 22704
rect 10612 22633 10640 22732
rect 14182 22720 14188 22732
rect 14240 22720 14246 22772
rect 14737 22763 14795 22769
rect 14737 22760 14749 22763
rect 14292 22732 14749 22760
rect 13998 22692 14004 22704
rect 13959 22664 14004 22692
rect 13998 22652 14004 22664
rect 14056 22692 14062 22704
rect 14292 22692 14320 22732
rect 14737 22729 14749 22732
rect 14783 22729 14795 22763
rect 15654 22760 15660 22772
rect 15615 22732 15660 22760
rect 14737 22723 14795 22729
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 19794 22760 19800 22772
rect 15764 22732 19800 22760
rect 15764 22692 15792 22732
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 19978 22760 19984 22772
rect 19939 22732 19984 22760
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20162 22720 20168 22772
rect 20220 22760 20226 22772
rect 20346 22760 20352 22772
rect 20220 22732 20352 22760
rect 20220 22720 20226 22732
rect 20346 22720 20352 22732
rect 20404 22720 20410 22772
rect 21637 22763 21695 22769
rect 21637 22729 21649 22763
rect 21683 22760 21695 22763
rect 21726 22760 21732 22772
rect 21683 22732 21732 22760
rect 21683 22729 21695 22732
rect 21637 22723 21695 22729
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 24026 22720 24032 22772
rect 24084 22760 24090 22772
rect 24121 22763 24179 22769
rect 24121 22760 24133 22763
rect 24084 22732 24133 22760
rect 24084 22720 24090 22732
rect 24121 22729 24133 22732
rect 24167 22729 24179 22763
rect 24121 22723 24179 22729
rect 24486 22720 24492 22772
rect 24544 22760 24550 22772
rect 25866 22760 25872 22772
rect 24544 22732 25872 22760
rect 24544 22720 24550 22732
rect 25866 22720 25872 22732
rect 25924 22720 25930 22772
rect 28445 22763 28503 22769
rect 28445 22729 28457 22763
rect 28491 22760 28503 22763
rect 28902 22760 28908 22772
rect 28491 22732 28908 22760
rect 28491 22729 28503 22732
rect 28445 22723 28503 22729
rect 28902 22720 28908 22732
rect 28960 22720 28966 22772
rect 28994 22720 29000 22772
rect 29052 22760 29058 22772
rect 30926 22760 30932 22772
rect 29052 22732 30932 22760
rect 29052 22720 29058 22732
rect 14056 22664 14320 22692
rect 14752 22664 15792 22692
rect 16301 22695 16359 22701
rect 14056 22652 14062 22664
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 10962 22624 10968 22636
rect 10735 22596 10968 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 10962 22584 10968 22596
rect 11020 22584 11026 22636
rect 11054 22584 11060 22636
rect 11112 22624 11118 22636
rect 11606 22624 11612 22636
rect 11112 22596 11612 22624
rect 11112 22584 11118 22596
rect 11606 22584 11612 22596
rect 11664 22624 11670 22636
rect 12069 22627 12127 22633
rect 12069 22624 12081 22627
rect 11664 22596 12081 22624
rect 11664 22584 11670 22596
rect 12069 22593 12081 22596
rect 12115 22593 12127 22627
rect 12069 22587 12127 22593
rect 14090 22584 14096 22636
rect 14148 22624 14154 22636
rect 14185 22627 14243 22633
rect 14185 22624 14197 22627
rect 14148 22596 14197 22624
rect 14148 22584 14154 22596
rect 14185 22593 14197 22596
rect 14231 22593 14243 22627
rect 14752 22624 14780 22664
rect 16301 22661 16313 22695
rect 16347 22692 16359 22695
rect 18690 22692 18696 22704
rect 16347 22664 18696 22692
rect 16347 22661 16359 22664
rect 16301 22655 16359 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 18782 22652 18788 22704
rect 18840 22692 18846 22704
rect 19334 22692 19340 22704
rect 18840 22664 19340 22692
rect 18840 22652 18846 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 19518 22692 19524 22704
rect 19479 22664 19524 22692
rect 19518 22652 19524 22664
rect 19576 22652 19582 22704
rect 30208 22701 30236 22732
rect 30926 22720 30932 22732
rect 30984 22720 30990 22772
rect 31202 22760 31208 22772
rect 31163 22732 31208 22760
rect 31202 22720 31208 22732
rect 31260 22720 31266 22772
rect 31386 22720 31392 22772
rect 31444 22760 31450 22772
rect 31665 22763 31723 22769
rect 31665 22760 31677 22763
rect 31444 22732 31677 22760
rect 31444 22720 31450 22732
rect 31665 22729 31677 22732
rect 31711 22729 31723 22763
rect 32398 22760 32404 22772
rect 31665 22723 31723 22729
rect 32048 22732 32404 22760
rect 25225 22695 25283 22701
rect 25225 22661 25237 22695
rect 25271 22661 25283 22695
rect 25225 22655 25283 22661
rect 29641 22695 29699 22701
rect 29641 22661 29653 22695
rect 29687 22661 29699 22695
rect 29641 22655 29699 22661
rect 30193 22695 30251 22701
rect 30193 22661 30205 22695
rect 30239 22661 30251 22695
rect 30193 22655 30251 22661
rect 30285 22695 30343 22701
rect 30285 22661 30297 22695
rect 30331 22692 30343 22695
rect 32048 22692 32076 22732
rect 32398 22720 32404 22732
rect 32456 22760 32462 22772
rect 35342 22760 35348 22772
rect 32456 22732 35348 22760
rect 32456 22720 32462 22732
rect 35342 22720 35348 22732
rect 35400 22720 35406 22772
rect 35986 22760 35992 22772
rect 35947 22732 35992 22760
rect 35986 22720 35992 22732
rect 36044 22720 36050 22772
rect 57974 22760 57980 22772
rect 57935 22732 57980 22760
rect 57974 22720 57980 22732
rect 58032 22720 58038 22772
rect 34241 22695 34299 22701
rect 34241 22692 34253 22695
rect 30331 22664 32076 22692
rect 32140 22664 34253 22692
rect 30331 22661 30343 22664
rect 30285 22655 30343 22661
rect 14185 22587 14243 22593
rect 14660 22596 14780 22624
rect 14921 22627 14979 22633
rect 7607 22528 9674 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 10042 22516 10048 22568
rect 10100 22556 10106 22568
rect 10318 22556 10324 22568
rect 10100 22528 10324 22556
rect 10100 22516 10106 22528
rect 10318 22516 10324 22528
rect 10376 22516 10382 22568
rect 10410 22516 10416 22568
rect 10468 22556 10474 22568
rect 10505 22559 10563 22565
rect 10505 22556 10517 22559
rect 10468 22528 10517 22556
rect 10468 22516 10474 22528
rect 10505 22525 10517 22528
rect 10551 22525 10563 22559
rect 10505 22519 10563 22525
rect 10778 22516 10784 22568
rect 10836 22556 10842 22568
rect 10873 22559 10931 22565
rect 10873 22556 10885 22559
rect 10836 22528 10885 22556
rect 10836 22516 10842 22528
rect 10873 22525 10885 22528
rect 10919 22525 10931 22559
rect 10980 22556 11008 22584
rect 11422 22556 11428 22568
rect 10980 22528 11428 22556
rect 10873 22519 10931 22525
rect 11422 22516 11428 22528
rect 11480 22516 11486 22568
rect 12158 22516 12164 22568
rect 12216 22556 12222 22568
rect 12325 22559 12383 22565
rect 12325 22556 12337 22559
rect 12216 22528 12337 22556
rect 12216 22516 12222 22528
rect 12325 22525 12337 22528
rect 12371 22525 12383 22559
rect 13906 22556 13912 22568
rect 13867 22528 13912 22556
rect 12325 22519 12383 22525
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 4617 22491 4675 22497
rect 4617 22488 4629 22491
rect 2746 22460 4629 22488
rect 2590 22380 2596 22432
rect 2648 22420 2654 22432
rect 2746 22420 2774 22460
rect 4617 22457 4629 22460
rect 4663 22488 4675 22491
rect 4798 22488 4804 22500
rect 4663 22460 4804 22488
rect 4663 22457 4675 22460
rect 4617 22451 4675 22457
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 4982 22488 4988 22500
rect 4943 22460 4988 22488
rect 4982 22448 4988 22460
rect 5040 22488 5046 22500
rect 5442 22488 5448 22500
rect 5040 22460 5448 22488
rect 5040 22448 5046 22460
rect 5442 22448 5448 22460
rect 5500 22448 5506 22500
rect 8748 22491 8806 22497
rect 8748 22457 8760 22491
rect 8794 22488 8806 22491
rect 11057 22491 11115 22497
rect 11057 22488 11069 22491
rect 8794 22460 11069 22488
rect 8794 22457 8806 22460
rect 8748 22451 8806 22457
rect 11057 22457 11069 22460
rect 11103 22457 11115 22491
rect 11698 22488 11704 22500
rect 11057 22451 11115 22457
rect 11440 22460 11704 22488
rect 2648 22392 2774 22420
rect 5813 22423 5871 22429
rect 2648 22380 2654 22392
rect 5813 22389 5825 22423
rect 5859 22420 5871 22423
rect 5902 22420 5908 22432
rect 5859 22392 5908 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 5902 22380 5908 22392
rect 5960 22420 5966 22432
rect 6270 22420 6276 22432
rect 5960 22392 6276 22420
rect 5960 22380 5966 22392
rect 6270 22380 6276 22392
rect 6328 22380 6334 22432
rect 7282 22380 7288 22432
rect 7340 22420 7346 22432
rect 7745 22423 7803 22429
rect 7745 22420 7757 22423
rect 7340 22392 7757 22420
rect 7340 22380 7346 22392
rect 7745 22389 7757 22392
rect 7791 22389 7803 22423
rect 7745 22383 7803 22389
rect 8110 22380 8116 22432
rect 8168 22420 8174 22432
rect 11440 22420 11468 22460
rect 11698 22448 11704 22460
rect 11756 22448 11762 22500
rect 14200 22488 14228 22587
rect 14660 22565 14688 22596
rect 14921 22593 14933 22627
rect 14967 22593 14979 22627
rect 19058 22624 19064 22636
rect 14921 22587 14979 22593
rect 17604 22596 19064 22624
rect 14645 22559 14703 22565
rect 14645 22525 14657 22559
rect 14691 22525 14703 22559
rect 14645 22519 14703 22525
rect 14936 22488 14964 22587
rect 15565 22559 15623 22565
rect 15565 22525 15577 22559
rect 15611 22556 15623 22559
rect 16114 22556 16120 22568
rect 15611 22528 16120 22556
rect 15611 22525 15623 22528
rect 15565 22519 15623 22525
rect 16114 22516 16120 22528
rect 16172 22516 16178 22568
rect 16209 22559 16267 22565
rect 16209 22525 16221 22559
rect 16255 22556 16267 22559
rect 17402 22556 17408 22568
rect 16255 22528 17408 22556
rect 16255 22525 16267 22528
rect 16209 22519 16267 22525
rect 17402 22516 17408 22528
rect 17460 22516 17466 22568
rect 17604 22565 17632 22596
rect 19058 22584 19064 22596
rect 19116 22624 19122 22636
rect 25240 22624 25268 22655
rect 19116 22596 19288 22624
rect 25240 22596 26372 22624
rect 19116 22584 19122 22596
rect 17589 22559 17647 22565
rect 17589 22525 17601 22559
rect 17635 22525 17647 22559
rect 18966 22556 18972 22568
rect 17589 22519 17647 22525
rect 18064 22528 18736 22556
rect 18927 22528 18972 22556
rect 14200 22460 14964 22488
rect 16390 22448 16396 22500
rect 16448 22488 16454 22500
rect 17954 22488 17960 22500
rect 16448 22460 17960 22488
rect 16448 22448 16454 22460
rect 17954 22448 17960 22460
rect 18012 22448 18018 22500
rect 8168 22392 11468 22420
rect 8168 22380 8174 22392
rect 11514 22380 11520 22432
rect 11572 22420 11578 22432
rect 13449 22423 13507 22429
rect 13449 22420 13461 22423
rect 11572 22392 13461 22420
rect 11572 22380 11578 22392
rect 13449 22389 13461 22392
rect 13495 22389 13507 22423
rect 14182 22420 14188 22432
rect 14143 22392 14188 22420
rect 13449 22383 13507 22389
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 14274 22380 14280 22432
rect 14332 22420 14338 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 14332 22392 14933 22420
rect 14332 22380 14338 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 17678 22420 17684 22432
rect 17639 22392 17684 22420
rect 14921 22383 14979 22389
rect 17678 22380 17684 22392
rect 17736 22420 17742 22432
rect 18064 22420 18092 22528
rect 18325 22491 18383 22497
rect 18325 22457 18337 22491
rect 18371 22488 18383 22491
rect 18598 22488 18604 22500
rect 18371 22460 18604 22488
rect 18371 22457 18383 22460
rect 18325 22451 18383 22457
rect 18598 22448 18604 22460
rect 18656 22448 18662 22500
rect 18708 22488 18736 22528
rect 18966 22516 18972 22528
rect 19024 22516 19030 22568
rect 19260 22565 19288 22596
rect 19245 22559 19303 22565
rect 19245 22525 19257 22559
rect 19291 22525 19303 22559
rect 19245 22519 19303 22525
rect 19334 22516 19340 22568
rect 19392 22556 19398 22568
rect 19392 22528 19437 22556
rect 19392 22516 19398 22528
rect 19518 22516 19524 22568
rect 19576 22556 19582 22568
rect 20070 22556 20076 22568
rect 19576 22528 20076 22556
rect 19576 22516 19582 22528
rect 20070 22516 20076 22528
rect 20128 22556 20134 22568
rect 20165 22559 20223 22565
rect 20165 22556 20177 22559
rect 20128 22528 20177 22556
rect 20128 22516 20134 22528
rect 20165 22525 20177 22528
rect 20211 22525 20223 22559
rect 20438 22556 20444 22568
rect 20399 22528 20444 22556
rect 20165 22519 20223 22525
rect 20438 22516 20444 22528
rect 20496 22516 20502 22568
rect 20990 22556 20996 22568
rect 20951 22528 20996 22556
rect 20990 22516 20996 22528
rect 21048 22516 21054 22568
rect 21082 22516 21088 22568
rect 21140 22556 21146 22568
rect 21450 22556 21456 22568
rect 21140 22528 21185 22556
rect 21409 22528 21456 22556
rect 21140 22516 21146 22528
rect 21450 22516 21456 22528
rect 21508 22565 21514 22568
rect 21508 22559 21557 22565
rect 21508 22525 21511 22559
rect 21545 22556 21557 22559
rect 21634 22556 21640 22568
rect 21545 22528 21640 22556
rect 21545 22525 21557 22528
rect 21508 22519 21557 22525
rect 21508 22516 21514 22519
rect 21634 22516 21640 22528
rect 21692 22516 21698 22568
rect 22646 22556 22652 22568
rect 22607 22528 22652 22556
rect 22646 22516 22652 22528
rect 22704 22516 22710 22568
rect 23753 22559 23811 22565
rect 23753 22525 23765 22559
rect 23799 22525 23811 22559
rect 23934 22556 23940 22568
rect 23895 22528 23940 22556
rect 23753 22519 23811 22525
rect 19153 22491 19211 22497
rect 19153 22488 19165 22491
rect 18708 22460 19165 22488
rect 19153 22457 19165 22460
rect 19199 22488 19211 22491
rect 20346 22488 20352 22500
rect 19199 22460 20352 22488
rect 19199 22457 19211 22460
rect 19153 22451 19211 22457
rect 20346 22448 20352 22460
rect 20404 22448 20410 22500
rect 20456 22488 20484 22516
rect 21269 22491 21327 22497
rect 21269 22488 21281 22491
rect 20456 22460 21281 22488
rect 21269 22457 21281 22460
rect 21315 22457 21327 22491
rect 21269 22451 21327 22457
rect 21358 22448 21364 22500
rect 21416 22488 21422 22500
rect 23768 22488 23796 22519
rect 23934 22516 23940 22528
rect 23992 22516 23998 22568
rect 24394 22516 24400 22568
rect 24452 22556 24458 22568
rect 24578 22556 24584 22568
rect 24452 22528 24584 22556
rect 24452 22516 24458 22528
rect 24578 22516 24584 22528
rect 24636 22516 24642 22568
rect 24670 22516 24676 22568
rect 24728 22556 24734 22568
rect 25087 22559 25145 22565
rect 24728 22528 24773 22556
rect 24728 22516 24734 22528
rect 25087 22525 25099 22559
rect 25133 22556 25145 22559
rect 25774 22556 25780 22568
rect 25133 22528 25780 22556
rect 25133 22525 25145 22528
rect 25087 22519 25145 22525
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 25866 22516 25872 22568
rect 25924 22556 25930 22568
rect 25961 22559 26019 22565
rect 25961 22556 25973 22559
rect 25924 22528 25973 22556
rect 25924 22516 25930 22528
rect 25961 22525 25973 22528
rect 26007 22525 26019 22559
rect 25961 22519 26019 22525
rect 26050 22559 26108 22565
rect 26050 22525 26062 22559
rect 26096 22525 26108 22559
rect 26050 22519 26108 22525
rect 24854 22488 24860 22500
rect 21416 22460 21461 22488
rect 23768 22460 23980 22488
rect 24815 22460 24860 22488
rect 21416 22448 21422 22460
rect 17736 22392 18092 22420
rect 18417 22423 18475 22429
rect 17736 22380 17742 22392
rect 18417 22389 18429 22423
rect 18463 22420 18475 22423
rect 18782 22420 18788 22432
rect 18463 22392 18788 22420
rect 18463 22389 18475 22392
rect 18417 22383 18475 22389
rect 18782 22380 18788 22392
rect 18840 22380 18846 22432
rect 18966 22380 18972 22432
rect 19024 22420 19030 22432
rect 20714 22420 20720 22432
rect 19024 22392 20720 22420
rect 19024 22380 19030 22392
rect 20714 22380 20720 22392
rect 20772 22380 20778 22432
rect 22741 22423 22799 22429
rect 22741 22389 22753 22423
rect 22787 22420 22799 22423
rect 23842 22420 23848 22432
rect 22787 22392 23848 22420
rect 22787 22389 22799 22392
rect 22741 22383 22799 22389
rect 23842 22380 23848 22392
rect 23900 22380 23906 22432
rect 23952 22420 23980 22460
rect 24854 22448 24860 22460
rect 24912 22448 24918 22500
rect 24946 22448 24952 22500
rect 25004 22488 25010 22500
rect 25004 22460 25049 22488
rect 25004 22448 25010 22460
rect 25130 22420 25136 22432
rect 23952 22392 25136 22420
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 25682 22420 25688 22432
rect 25643 22392 25688 22420
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 26068 22420 26096 22519
rect 26142 22516 26148 22568
rect 26200 22556 26206 22568
rect 26344 22565 26372 22596
rect 26418 22584 26424 22636
rect 26476 22624 26482 22636
rect 29656 22624 29684 22655
rect 30377 22627 30435 22633
rect 26476 22596 29592 22624
rect 29656 22596 30328 22624
rect 26476 22584 26482 22596
rect 26329 22559 26387 22565
rect 26200 22528 26245 22556
rect 26200 22516 26206 22528
rect 26329 22525 26341 22559
rect 26375 22525 26387 22559
rect 26329 22519 26387 22525
rect 27338 22516 27344 22568
rect 27396 22556 27402 22568
rect 27801 22559 27859 22565
rect 27801 22556 27813 22559
rect 27396 22528 27813 22556
rect 27396 22516 27402 22528
rect 27801 22525 27813 22528
rect 27847 22525 27859 22559
rect 27801 22519 27859 22525
rect 28445 22559 28503 22565
rect 28445 22525 28457 22559
rect 28491 22556 28503 22559
rect 28534 22556 28540 22568
rect 28491 22528 28540 22556
rect 28491 22525 28503 22528
rect 28445 22519 28503 22525
rect 28534 22516 28540 22528
rect 28592 22516 28598 22568
rect 28626 22516 28632 22568
rect 28684 22556 28690 22568
rect 28684 22528 28729 22556
rect 28684 22516 28690 22528
rect 28994 22516 29000 22568
rect 29052 22556 29058 22568
rect 29089 22559 29147 22565
rect 29089 22556 29101 22559
rect 29052 22528 29101 22556
rect 29052 22516 29058 22528
rect 29089 22525 29101 22528
rect 29135 22525 29147 22559
rect 29270 22556 29276 22568
rect 29231 22528 29276 22556
rect 29089 22519 29147 22525
rect 29270 22516 29276 22528
rect 29328 22516 29334 22568
rect 29454 22556 29460 22568
rect 29415 22528 29460 22556
rect 29454 22516 29460 22528
rect 29512 22516 29518 22568
rect 29362 22448 29368 22500
rect 29420 22488 29426 22500
rect 29420 22460 29465 22488
rect 29420 22448 29426 22460
rect 27614 22420 27620 22432
rect 26068 22392 27620 22420
rect 27614 22380 27620 22392
rect 27672 22380 27678 22432
rect 27890 22420 27896 22432
rect 27851 22392 27896 22420
rect 27890 22380 27896 22392
rect 27948 22380 27954 22432
rect 29564 22420 29592 22596
rect 30300 22568 30328 22596
rect 30377 22593 30389 22627
rect 30423 22624 30435 22627
rect 30558 22624 30564 22636
rect 30423 22596 30564 22624
rect 30423 22593 30435 22596
rect 30377 22587 30435 22593
rect 30558 22584 30564 22596
rect 30616 22584 30622 22636
rect 31570 22584 31576 22636
rect 31628 22624 31634 22636
rect 32140 22624 32168 22664
rect 34241 22661 34253 22664
rect 34287 22692 34299 22695
rect 34514 22692 34520 22704
rect 34287 22664 34520 22692
rect 34287 22661 34299 22664
rect 34241 22655 34299 22661
rect 34514 22652 34520 22664
rect 34572 22652 34578 22704
rect 54849 22695 54907 22701
rect 54849 22661 54861 22695
rect 54895 22692 54907 22695
rect 54895 22664 55720 22692
rect 54895 22661 54907 22664
rect 54849 22655 54907 22661
rect 31628 22596 32168 22624
rect 31628 22584 31634 22596
rect 32214 22584 32220 22636
rect 32272 22624 32278 22636
rect 33594 22624 33600 22636
rect 32272 22596 33600 22624
rect 32272 22584 32278 22596
rect 33594 22584 33600 22596
rect 33652 22584 33658 22636
rect 34532 22624 34560 22652
rect 55692 22633 55720 22664
rect 55677 22627 55735 22633
rect 34532 22596 36216 22624
rect 30101 22559 30159 22565
rect 30101 22525 30113 22559
rect 30147 22525 30159 22559
rect 30282 22556 30288 22568
rect 30195 22528 30288 22556
rect 30101 22519 30159 22525
rect 30116 22488 30144 22519
rect 30282 22516 30288 22528
rect 30340 22556 30346 22568
rect 30837 22559 30895 22565
rect 30837 22556 30849 22559
rect 30340 22528 30849 22556
rect 30340 22516 30346 22528
rect 30837 22525 30849 22528
rect 30883 22525 30895 22559
rect 30837 22519 30895 22525
rect 31202 22516 31208 22568
rect 31260 22556 31266 22568
rect 31665 22559 31723 22565
rect 31665 22556 31677 22559
rect 31260 22528 31677 22556
rect 31260 22516 31266 22528
rect 31665 22525 31677 22528
rect 31711 22525 31723 22559
rect 31665 22519 31723 22525
rect 31849 22559 31907 22565
rect 31849 22525 31861 22559
rect 31895 22556 31907 22559
rect 33045 22559 33103 22565
rect 31895 22528 32352 22556
rect 31895 22525 31907 22528
rect 31849 22519 31907 22525
rect 30374 22488 30380 22500
rect 30116 22460 30380 22488
rect 30374 22448 30380 22460
rect 30432 22448 30438 22500
rect 31021 22491 31079 22497
rect 31021 22457 31033 22491
rect 31067 22488 31079 22491
rect 31754 22488 31760 22500
rect 31067 22460 31760 22488
rect 31067 22457 31079 22460
rect 31021 22451 31079 22457
rect 31754 22448 31760 22460
rect 31812 22448 31818 22500
rect 32324 22432 32352 22528
rect 33045 22525 33057 22559
rect 33091 22556 33103 22559
rect 33226 22556 33232 22568
rect 33091 22528 33232 22556
rect 33091 22525 33103 22528
rect 33045 22519 33103 22525
rect 33226 22516 33232 22528
rect 33284 22516 33290 22568
rect 34146 22556 34152 22568
rect 34107 22528 34152 22556
rect 34146 22516 34152 22528
rect 34204 22516 34210 22568
rect 35342 22556 35348 22568
rect 35303 22528 35348 22556
rect 35342 22516 35348 22528
rect 35400 22516 35406 22568
rect 35986 22556 35992 22568
rect 35947 22528 35992 22556
rect 35986 22516 35992 22528
rect 36044 22516 36050 22568
rect 36188 22565 36216 22596
rect 55677 22593 55689 22627
rect 55723 22593 55735 22627
rect 57514 22624 57520 22636
rect 57475 22596 57520 22624
rect 55677 22587 55735 22593
rect 57514 22584 57520 22596
rect 57572 22584 57578 22636
rect 36173 22559 36231 22565
rect 36173 22525 36185 22559
rect 36219 22525 36231 22559
rect 55030 22556 55036 22568
rect 54991 22528 55036 22556
rect 36173 22519 36231 22525
rect 55030 22516 55036 22528
rect 55088 22516 55094 22568
rect 55490 22556 55496 22568
rect 55451 22528 55496 22556
rect 55490 22516 55496 22528
rect 55548 22516 55554 22568
rect 56410 22516 56416 22568
rect 56468 22556 56474 22568
rect 57701 22559 57759 22565
rect 57701 22556 57713 22559
rect 56468 22528 57713 22556
rect 56468 22516 56474 22528
rect 57701 22525 57713 22528
rect 57747 22525 57759 22559
rect 57701 22519 57759 22525
rect 32398 22448 32404 22500
rect 32456 22488 32462 22500
rect 34606 22488 34612 22500
rect 32456 22460 34612 22488
rect 32456 22448 32462 22460
rect 34606 22448 34612 22460
rect 34664 22448 34670 22500
rect 56137 22491 56195 22497
rect 56137 22457 56149 22491
rect 56183 22488 56195 22491
rect 56873 22491 56931 22497
rect 56873 22488 56885 22491
rect 56183 22460 56885 22488
rect 56183 22457 56195 22460
rect 56137 22451 56195 22457
rect 56873 22457 56885 22460
rect 56919 22457 56931 22491
rect 57054 22488 57060 22500
rect 57015 22460 57060 22488
rect 56873 22451 56931 22457
rect 57054 22448 57060 22460
rect 57112 22448 57118 22500
rect 31938 22420 31944 22432
rect 29564 22392 31944 22420
rect 31938 22380 31944 22392
rect 31996 22380 32002 22432
rect 32030 22380 32036 22432
rect 32088 22420 32094 22432
rect 32088 22392 32133 22420
rect 32088 22380 32094 22392
rect 32306 22380 32312 22432
rect 32364 22420 32370 22432
rect 33137 22423 33195 22429
rect 33137 22420 33149 22423
rect 32364 22392 33149 22420
rect 32364 22380 32370 22392
rect 33137 22389 33149 22392
rect 33183 22389 33195 22423
rect 35434 22420 35440 22432
rect 35395 22392 35440 22420
rect 33137 22383 33195 22389
rect 35434 22380 35440 22392
rect 35492 22380 35498 22432
rect 1104 22330 58880 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 50326 22330
rect 50378 22278 50390 22330
rect 50442 22278 50454 22330
rect 50506 22278 50518 22330
rect 50570 22278 58880 22330
rect 1104 22256 58880 22278
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 4356 22188 7849 22216
rect 4356 22157 4384 22188
rect 7837 22185 7849 22188
rect 7883 22185 7895 22219
rect 7837 22179 7895 22185
rect 10318 22176 10324 22228
rect 10376 22216 10382 22228
rect 10962 22216 10968 22228
rect 10376 22188 10968 22216
rect 10376 22176 10382 22188
rect 10962 22176 10968 22188
rect 11020 22176 11026 22228
rect 11348 22188 12020 22216
rect 4341 22151 4399 22157
rect 4341 22117 4353 22151
rect 4387 22117 4399 22151
rect 4341 22111 4399 22117
rect 4433 22151 4491 22157
rect 4433 22117 4445 22151
rect 4479 22148 4491 22151
rect 6730 22148 6736 22160
rect 4479 22120 6736 22148
rect 4479 22117 4491 22120
rect 4433 22111 4491 22117
rect 6730 22108 6736 22120
rect 6788 22108 6794 22160
rect 8202 22148 8208 22160
rect 6840 22120 8208 22148
rect 3237 22083 3295 22089
rect 3237 22049 3249 22083
rect 3283 22080 3295 22083
rect 3418 22080 3424 22092
rect 3283 22052 3424 22080
rect 3283 22049 3295 22052
rect 3237 22043 3295 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 5534 22080 5540 22092
rect 5495 22052 5540 22080
rect 5534 22040 5540 22052
rect 5592 22040 5598 22092
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 6638 22080 6644 22092
rect 6599 22052 6644 22080
rect 6638 22040 6644 22052
rect 6696 22040 6702 22092
rect 6840 22089 6868 22120
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 10410 22148 10416 22160
rect 10152 22120 10416 22148
rect 6825 22083 6883 22089
rect 6825 22049 6837 22083
rect 6871 22049 6883 22083
rect 7558 22080 7564 22092
rect 7519 22052 7564 22080
rect 6825 22043 6883 22049
rect 7558 22040 7564 22052
rect 7616 22040 7622 22092
rect 7653 22083 7711 22089
rect 7653 22049 7665 22083
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 9674 22080 9680 22092
rect 8343 22052 9680 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 1949 22015 2007 22021
rect 1949 21981 1961 22015
rect 1995 21981 2007 22015
rect 1949 21975 2007 21981
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 4062 22012 4068 22024
rect 2179 21984 4068 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 1964 21944 1992 21975
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 7668 22012 7696 22043
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10042 22080 10048 22092
rect 9999 22052 10048 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10042 22040 10048 22052
rect 10100 22040 10106 22092
rect 10152 22089 10180 22120
rect 10410 22108 10416 22120
rect 10468 22148 10474 22160
rect 11146 22148 11152 22160
rect 10468 22120 11152 22148
rect 10468 22108 10474 22120
rect 11146 22108 11152 22120
rect 11204 22108 11210 22160
rect 11348 22148 11376 22188
rect 11992 22160 12020 22188
rect 13906 22176 13912 22228
rect 13964 22216 13970 22228
rect 32214 22216 32220 22228
rect 13964 22188 32220 22216
rect 13964 22176 13970 22188
rect 32214 22176 32220 22188
rect 32272 22176 32278 22228
rect 33226 22216 33232 22228
rect 32416 22188 33232 22216
rect 11256 22120 11376 22148
rect 11256 22092 11284 22120
rect 11422 22108 11428 22160
rect 11480 22148 11486 22160
rect 11974 22148 11980 22160
rect 11480 22120 11525 22148
rect 11935 22120 11980 22148
rect 11480 22108 11486 22120
rect 11974 22108 11980 22120
rect 12032 22108 12038 22160
rect 12713 22151 12771 22157
rect 12713 22117 12725 22151
rect 12759 22148 12771 22151
rect 13357 22151 13415 22157
rect 13357 22148 13369 22151
rect 12759 22120 13369 22148
rect 12759 22117 12771 22120
rect 12713 22111 12771 22117
rect 13357 22117 13369 22120
rect 13403 22148 13415 22151
rect 14829 22151 14887 22157
rect 14829 22148 14841 22151
rect 13403 22120 14841 22148
rect 13403 22117 13415 22120
rect 13357 22111 13415 22117
rect 14829 22117 14841 22120
rect 14875 22117 14887 22151
rect 20993 22151 21051 22157
rect 14829 22111 14887 22117
rect 15304 22120 15700 22148
rect 10137 22083 10195 22089
rect 10137 22049 10149 22083
rect 10183 22049 10195 22083
rect 10318 22080 10324 22092
rect 10279 22052 10324 22080
rect 10137 22043 10195 22049
rect 10318 22040 10324 22052
rect 10376 22040 10382 22092
rect 10502 22080 10508 22092
rect 10463 22052 10508 22080
rect 10502 22040 10508 22052
rect 10560 22040 10566 22092
rect 11238 22080 11244 22092
rect 11151 22052 11244 22080
rect 11238 22040 11244 22052
rect 11296 22040 11302 22092
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12342 22080 12348 22092
rect 12124 22052 12348 22080
rect 12124 22040 12130 22052
rect 12342 22040 12348 22052
rect 12400 22080 12406 22092
rect 12621 22083 12679 22089
rect 12621 22080 12633 22083
rect 12400 22052 12633 22080
rect 12400 22040 12406 22052
rect 12621 22049 12633 22052
rect 12667 22049 12679 22083
rect 12621 22043 12679 22049
rect 15010 22040 15016 22092
rect 15068 22080 15074 22092
rect 15304 22080 15332 22120
rect 15068 22052 15332 22080
rect 15068 22040 15074 22052
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 15672 22089 15700 22120
rect 18156 22120 18644 22148
rect 15473 22083 15531 22089
rect 15473 22080 15485 22083
rect 15436 22052 15485 22080
rect 15436 22040 15442 22052
rect 15473 22049 15485 22052
rect 15519 22049 15531 22083
rect 15473 22043 15531 22049
rect 15657 22083 15715 22089
rect 15657 22049 15669 22083
rect 15703 22080 15715 22083
rect 15703 22052 15737 22080
rect 15703 22049 15715 22052
rect 15657 22043 15715 22049
rect 15838 22040 15844 22092
rect 15896 22080 15902 22092
rect 18156 22089 18184 22120
rect 16373 22083 16431 22089
rect 16373 22080 16385 22083
rect 15896 22052 16385 22080
rect 15896 22040 15902 22052
rect 16373 22049 16385 22052
rect 16419 22049 16431 22083
rect 16373 22043 16431 22049
rect 18124 22083 18184 22089
rect 18124 22049 18136 22083
rect 18170 22052 18184 22083
rect 18170 22049 18182 22052
rect 18124 22043 18182 22049
rect 18230 22040 18236 22092
rect 18288 22080 18294 22092
rect 18506 22080 18512 22092
rect 18288 22052 18333 22080
rect 18467 22052 18512 22080
rect 18288 22040 18294 22052
rect 18506 22040 18512 22052
rect 18564 22040 18570 22092
rect 10229 22015 10287 22021
rect 7668 21984 10088 22012
rect 3050 21944 3056 21956
rect 1964 21916 2774 21944
rect 3011 21916 3056 21944
rect 2314 21876 2320 21888
rect 2275 21848 2320 21876
rect 2314 21836 2320 21848
rect 2372 21836 2378 21888
rect 2746 21876 2774 21916
rect 3050 21904 3056 21916
rect 3108 21904 3114 21956
rect 4890 21944 4896 21956
rect 4851 21916 4896 21944
rect 4890 21904 4896 21916
rect 4948 21904 4954 21956
rect 10060 21944 10088 21984
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 14182 22012 14188 22024
rect 10275 21984 14188 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 14182 21972 14188 21984
rect 14240 21972 14246 22024
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15988 21984 16129 22012
rect 15988 21972 15994 21984
rect 16117 21981 16129 21984
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 18380 21984 18429 22012
rect 18380 21972 18386 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 11514 21944 11520 21956
rect 10060 21916 11520 21944
rect 11514 21904 11520 21916
rect 11572 21904 11578 21956
rect 12161 21947 12219 21953
rect 12161 21913 12173 21947
rect 12207 21944 12219 21947
rect 12434 21944 12440 21956
rect 12207 21916 12440 21944
rect 12207 21913 12219 21916
rect 12161 21907 12219 21913
rect 12434 21904 12440 21916
rect 12492 21904 12498 21956
rect 12986 21904 12992 21956
rect 13044 21944 13050 21956
rect 14274 21944 14280 21956
rect 13044 21916 14280 21944
rect 13044 21904 13050 21916
rect 14274 21904 14280 21916
rect 14332 21904 14338 21956
rect 15286 21904 15292 21956
rect 15344 21944 15350 21956
rect 15473 21947 15531 21953
rect 15473 21944 15485 21947
rect 15344 21916 15485 21944
rect 15344 21904 15350 21916
rect 15473 21913 15485 21916
rect 15519 21913 15531 21947
rect 18616 21944 18644 22120
rect 20993 22117 21005 22151
rect 21039 22148 21051 22151
rect 22186 22148 22192 22160
rect 21039 22120 22192 22148
rect 21039 22117 21051 22120
rect 20993 22111 21051 22117
rect 22186 22108 22192 22120
rect 22244 22108 22250 22160
rect 23934 22148 23940 22160
rect 23895 22120 23940 22148
rect 23934 22108 23940 22120
rect 23992 22108 23998 22160
rect 24121 22151 24179 22157
rect 24121 22117 24133 22151
rect 24167 22148 24179 22151
rect 25130 22148 25136 22160
rect 24167 22120 25136 22148
rect 24167 22117 24179 22120
rect 24121 22111 24179 22117
rect 25130 22108 25136 22120
rect 25188 22108 25194 22160
rect 25314 22148 25320 22160
rect 25275 22120 25320 22148
rect 25314 22108 25320 22120
rect 25372 22108 25378 22160
rect 25682 22108 25688 22160
rect 25740 22108 25746 22160
rect 26482 22151 26540 22157
rect 26482 22148 26494 22151
rect 26160 22120 26494 22148
rect 20070 22080 20076 22092
rect 20031 22052 20076 22080
rect 20070 22040 20076 22052
rect 20128 22040 20134 22092
rect 21637 22083 21695 22089
rect 21637 22049 21649 22083
rect 21683 22080 21695 22083
rect 21818 22080 21824 22092
rect 21683 22052 21824 22080
rect 21683 22049 21695 22052
rect 21637 22043 21695 22049
rect 21818 22040 21824 22052
rect 21876 22040 21882 22092
rect 22554 22080 22560 22092
rect 22467 22052 22560 22080
rect 22554 22040 22560 22052
rect 22612 22080 22618 22092
rect 25222 22080 25228 22092
rect 22612 22052 25228 22080
rect 22612 22040 22618 22052
rect 25222 22040 25228 22052
rect 25280 22040 25286 22092
rect 25498 22080 25504 22092
rect 25459 22052 25504 22080
rect 25498 22040 25504 22052
rect 25556 22040 25562 22092
rect 25700 22080 25728 22108
rect 26160 22080 26188 22120
rect 26482 22117 26494 22120
rect 26528 22117 26540 22151
rect 26482 22111 26540 22117
rect 27890 22108 27896 22160
rect 27948 22148 27954 22160
rect 30834 22148 30840 22160
rect 27948 22120 30840 22148
rect 27948 22108 27954 22120
rect 30834 22108 30840 22120
rect 30892 22108 30898 22160
rect 31386 22148 31392 22160
rect 31036 22120 31392 22148
rect 25700 22052 26188 22080
rect 26237 22083 26295 22089
rect 26237 22049 26249 22083
rect 26283 22049 26295 22083
rect 26237 22043 26295 22049
rect 28436 22083 28494 22089
rect 28436 22049 28448 22083
rect 28482 22080 28494 22083
rect 29178 22080 29184 22092
rect 28482 22052 29184 22080
rect 28482 22049 28494 22052
rect 28436 22043 28494 22049
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 20165 22015 20223 22021
rect 20165 22012 20177 22015
rect 19760 21984 20177 22012
rect 19760 21972 19766 21984
rect 20165 21981 20177 21984
rect 20211 22012 20223 22015
rect 20438 22012 20444 22024
rect 20211 21984 20444 22012
rect 20211 21981 20223 21984
rect 20165 21975 20223 21981
rect 20438 21972 20444 21984
rect 20496 21972 20502 22024
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 20772 21984 21741 22012
rect 20772 21972 20778 21984
rect 21729 21981 21741 21984
rect 21775 21981 21787 22015
rect 22830 22012 22836 22024
rect 22791 21984 22836 22012
rect 21729 21975 21787 21981
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 25590 21972 25596 22024
rect 25648 22012 25654 22024
rect 26243 22012 26271 22043
rect 29178 22040 29184 22052
rect 29236 22040 29242 22092
rect 30742 22080 30748 22092
rect 30703 22052 30748 22080
rect 30742 22040 30748 22052
rect 30800 22040 30806 22092
rect 31036 22089 31064 22120
rect 31386 22108 31392 22120
rect 31444 22108 31450 22160
rect 32306 22148 32312 22160
rect 32267 22120 32312 22148
rect 32306 22108 32312 22120
rect 32364 22108 32370 22160
rect 32416 22157 32444 22188
rect 33226 22176 33232 22188
rect 33284 22176 33290 22228
rect 33594 22176 33600 22228
rect 33652 22216 33658 22228
rect 35434 22216 35440 22228
rect 33652 22188 35440 22216
rect 33652 22176 33658 22188
rect 35434 22176 35440 22188
rect 35492 22176 35498 22228
rect 36357 22219 36415 22225
rect 36357 22185 36369 22219
rect 36403 22216 36415 22219
rect 38746 22216 38752 22228
rect 36403 22188 38752 22216
rect 36403 22185 36415 22188
rect 36357 22179 36415 22185
rect 38746 22176 38752 22188
rect 38804 22176 38810 22228
rect 55214 22216 55220 22228
rect 39040 22188 55220 22216
rect 32401 22151 32459 22157
rect 32401 22117 32413 22151
rect 32447 22117 32459 22151
rect 32401 22111 32459 22117
rect 33318 22108 33324 22160
rect 33376 22108 33382 22160
rect 37277 22151 37335 22157
rect 36096 22120 36952 22148
rect 30929 22083 30987 22089
rect 30929 22049 30941 22083
rect 30975 22049 30987 22083
rect 30929 22043 30987 22049
rect 31021 22083 31079 22089
rect 31021 22049 31033 22083
rect 31067 22080 31079 22083
rect 31205 22083 31263 22089
rect 31067 22052 31101 22080
rect 31067 22049 31079 22052
rect 31021 22043 31079 22049
rect 31205 22049 31217 22083
rect 31251 22080 31263 22083
rect 31294 22080 31300 22092
rect 31251 22052 31300 22080
rect 31251 22049 31263 22052
rect 31205 22043 31263 22049
rect 25648 21984 26271 22012
rect 25648 21972 25654 21984
rect 27798 21972 27804 22024
rect 27856 22012 27862 22024
rect 28169 22015 28227 22021
rect 28169 22012 28181 22015
rect 27856 21984 28181 22012
rect 27856 21972 27862 21984
rect 28169 21981 28181 21984
rect 28215 21981 28227 22015
rect 30944 22012 30972 22043
rect 31294 22040 31300 22052
rect 31352 22040 31358 22092
rect 32030 22080 32036 22092
rect 31991 22052 32036 22080
rect 32030 22040 32036 22052
rect 32088 22040 32094 22092
rect 32214 22089 32220 22092
rect 32181 22083 32220 22089
rect 32181 22049 32193 22083
rect 32181 22043 32220 22049
rect 32214 22040 32220 22043
rect 32272 22040 32278 22092
rect 32324 22012 32352 22108
rect 32490 22040 32496 22092
rect 32548 22089 32554 22092
rect 32548 22080 32556 22089
rect 33336 22080 33364 22108
rect 36096 22092 36124 22120
rect 33413 22083 33471 22089
rect 33413 22080 33425 22083
rect 32548 22052 32593 22080
rect 33336 22052 33425 22080
rect 32548 22043 32556 22052
rect 33413 22049 33425 22052
rect 33459 22049 33471 22083
rect 33413 22043 33471 22049
rect 33505 22083 33563 22089
rect 33505 22049 33517 22083
rect 33551 22049 33563 22083
rect 33505 22043 33563 22049
rect 33597 22083 33655 22089
rect 33597 22049 33609 22083
rect 33643 22080 33655 22083
rect 33686 22080 33692 22092
rect 33643 22052 33692 22080
rect 33643 22049 33655 22052
rect 33597 22043 33655 22049
rect 32548 22040 32554 22043
rect 30944 21984 32352 22012
rect 28169 21975 28227 21981
rect 33318 21972 33324 22024
rect 33376 22012 33382 22024
rect 33520 22012 33548 22043
rect 33686 22040 33692 22052
rect 33744 22040 33750 22092
rect 33778 22040 33784 22092
rect 33836 22080 33842 22092
rect 34241 22083 34299 22089
rect 33836 22052 33881 22080
rect 33836 22040 33842 22052
rect 34241 22049 34253 22083
rect 34287 22049 34299 22083
rect 36078 22080 36084 22092
rect 35991 22052 36084 22080
rect 34241 22043 34299 22049
rect 34256 22012 34284 22043
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 36262 22080 36268 22092
rect 36223 22052 36268 22080
rect 36262 22040 36268 22052
rect 36320 22040 36326 22092
rect 36924 22089 36952 22120
rect 37277 22117 37289 22151
rect 37323 22148 37335 22151
rect 39040 22148 39068 22188
rect 55214 22176 55220 22188
rect 55272 22176 55278 22228
rect 37323 22120 39068 22148
rect 37323 22117 37335 22120
rect 37277 22111 37335 22117
rect 39114 22108 39120 22160
rect 39172 22148 39178 22160
rect 55490 22148 55496 22160
rect 39172 22120 55496 22148
rect 39172 22108 39178 22120
rect 55490 22108 55496 22120
rect 55548 22108 55554 22160
rect 36909 22083 36967 22089
rect 36909 22049 36921 22083
rect 36955 22049 36967 22083
rect 36909 22043 36967 22049
rect 37093 22083 37151 22089
rect 37093 22049 37105 22083
rect 37139 22049 37151 22083
rect 37093 22043 37151 22049
rect 33376 21984 34284 22012
rect 33376 21972 33382 21984
rect 23566 21944 23572 21956
rect 18616 21916 23572 21944
rect 15473 21907 15531 21913
rect 23566 21904 23572 21916
rect 23624 21904 23630 21956
rect 27614 21944 27620 21956
rect 27575 21916 27620 21944
rect 27614 21904 27620 21916
rect 27672 21904 27678 21956
rect 31110 21944 31116 21956
rect 31071 21916 31116 21944
rect 31110 21904 31116 21916
rect 31168 21904 31174 21956
rect 32677 21947 32735 21953
rect 32677 21913 32689 21947
rect 32723 21944 32735 21947
rect 32723 21916 33364 21944
rect 32723 21913 32735 21916
rect 32677 21907 32735 21913
rect 7009 21879 7067 21885
rect 7009 21876 7021 21879
rect 2746 21848 7021 21876
rect 7009 21845 7021 21848
rect 7055 21845 7067 21879
rect 7009 21839 7067 21845
rect 8202 21836 8208 21888
rect 8260 21876 8266 21888
rect 8481 21879 8539 21885
rect 8481 21876 8493 21879
rect 8260 21848 8493 21876
rect 8260 21836 8266 21848
rect 8481 21845 8493 21848
rect 8527 21845 8539 21879
rect 8481 21839 8539 21845
rect 8846 21836 8852 21888
rect 8904 21876 8910 21888
rect 10689 21879 10747 21885
rect 10689 21876 10701 21879
rect 8904 21848 10701 21876
rect 8904 21836 8910 21848
rect 10689 21845 10701 21848
rect 10735 21845 10747 21879
rect 10689 21839 10747 21845
rect 11974 21836 11980 21888
rect 12032 21876 12038 21888
rect 13449 21879 13507 21885
rect 13449 21876 13461 21879
rect 12032 21848 13461 21876
rect 12032 21836 12038 21848
rect 13449 21845 13461 21848
rect 13495 21845 13507 21879
rect 13449 21839 13507 21845
rect 14921 21879 14979 21885
rect 14921 21845 14933 21879
rect 14967 21876 14979 21879
rect 15194 21876 15200 21888
rect 14967 21848 15200 21876
rect 14967 21845 14979 21848
rect 14921 21839 14979 21845
rect 15194 21836 15200 21848
rect 15252 21876 15258 21888
rect 15378 21876 15384 21888
rect 15252 21848 15384 21876
rect 15252 21836 15258 21848
rect 15378 21836 15384 21848
rect 15436 21876 15442 21888
rect 16114 21876 16120 21888
rect 15436 21848 16120 21876
rect 15436 21836 15442 21848
rect 16114 21836 16120 21848
rect 16172 21836 16178 21888
rect 17494 21876 17500 21888
rect 17455 21848 17500 21876
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17644 21848 17969 21876
rect 17644 21836 17650 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 18196 21848 20085 21876
rect 18196 21836 18202 21848
rect 20073 21845 20085 21848
rect 20119 21876 20131 21879
rect 20162 21876 20168 21888
rect 20119 21848 20168 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20346 21836 20352 21888
rect 20404 21876 20410 21888
rect 20441 21879 20499 21885
rect 20441 21876 20453 21879
rect 20404 21848 20453 21876
rect 20404 21836 20410 21848
rect 20441 21845 20453 21848
rect 20487 21845 20499 21879
rect 20441 21839 20499 21845
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 21085 21879 21143 21885
rect 21085 21876 21097 21879
rect 20956 21848 21097 21876
rect 20956 21836 20962 21848
rect 21085 21845 21097 21848
rect 21131 21876 21143 21879
rect 23014 21876 23020 21888
rect 21131 21848 23020 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 23014 21836 23020 21848
rect 23072 21836 23078 21888
rect 24305 21879 24363 21885
rect 24305 21845 24317 21879
rect 24351 21876 24363 21879
rect 24394 21876 24400 21888
rect 24351 21848 24400 21876
rect 24351 21845 24363 21848
rect 24305 21839 24363 21845
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 29086 21836 29092 21888
rect 29144 21876 29150 21888
rect 29454 21876 29460 21888
rect 29144 21848 29460 21876
rect 29144 21836 29150 21848
rect 29454 21836 29460 21848
rect 29512 21876 29518 21888
rect 29549 21879 29607 21885
rect 29549 21876 29561 21879
rect 29512 21848 29561 21876
rect 29512 21836 29518 21848
rect 29549 21845 29561 21848
rect 29595 21845 29607 21879
rect 29549 21839 29607 21845
rect 31294 21836 31300 21888
rect 31352 21876 31358 21888
rect 32950 21876 32956 21888
rect 31352 21848 32956 21876
rect 31352 21836 31358 21848
rect 32950 21836 32956 21848
rect 33008 21836 33014 21888
rect 33134 21876 33140 21888
rect 33095 21848 33140 21876
rect 33134 21836 33140 21848
rect 33192 21836 33198 21888
rect 33336 21876 33364 21916
rect 35434 21904 35440 21956
rect 35492 21944 35498 21956
rect 37108 21944 37136 22043
rect 55030 22040 55036 22092
rect 55088 22080 55094 22092
rect 55125 22083 55183 22089
rect 55125 22080 55137 22083
rect 55088 22052 55137 22080
rect 55088 22040 55094 22052
rect 55125 22049 55137 22052
rect 55171 22080 55183 22083
rect 55766 22080 55772 22092
rect 55171 22052 55772 22080
rect 55171 22049 55183 22052
rect 55125 22043 55183 22049
rect 55766 22040 55772 22052
rect 55824 22040 55830 22092
rect 57974 22080 57980 22092
rect 57935 22052 57980 22080
rect 57974 22040 57980 22052
rect 58032 22040 58038 22092
rect 48038 21972 48044 22024
rect 48096 22012 48102 22024
rect 56689 22015 56747 22021
rect 56689 22012 56701 22015
rect 48096 21984 56701 22012
rect 48096 21972 48102 21984
rect 56689 21981 56701 21984
rect 56735 21981 56747 22015
rect 56689 21975 56747 21981
rect 56873 22015 56931 22021
rect 56873 21981 56885 22015
rect 56919 21981 56931 22015
rect 56873 21975 56931 21981
rect 57333 22015 57391 22021
rect 57333 21981 57345 22015
rect 57379 22012 57391 22015
rect 58066 22012 58072 22024
rect 57379 21984 58072 22012
rect 57379 21981 57391 21984
rect 57333 21975 57391 21981
rect 35492 21916 37136 21944
rect 54941 21947 54999 21953
rect 35492 21904 35498 21916
rect 54941 21913 54953 21947
rect 54987 21944 54999 21947
rect 56888 21944 56916 21975
rect 58066 21972 58072 21984
rect 58124 21972 58130 22024
rect 58158 21944 58164 21956
rect 54987 21916 56916 21944
rect 58119 21916 58164 21944
rect 54987 21913 54999 21916
rect 54941 21907 54999 21913
rect 58158 21904 58164 21916
rect 58216 21904 58222 21956
rect 33778 21876 33784 21888
rect 33336 21848 33784 21876
rect 33778 21836 33784 21848
rect 33836 21836 33842 21888
rect 34333 21879 34391 21885
rect 34333 21845 34345 21879
rect 34379 21876 34391 21879
rect 34514 21876 34520 21888
rect 34379 21848 34520 21876
rect 34379 21845 34391 21848
rect 34333 21839 34391 21845
rect 34514 21836 34520 21848
rect 34572 21836 34578 21888
rect 55585 21879 55643 21885
rect 55585 21845 55597 21879
rect 55631 21876 55643 21879
rect 55858 21876 55864 21888
rect 55631 21848 55864 21876
rect 55631 21845 55643 21848
rect 55585 21839 55643 21845
rect 55858 21836 55864 21848
rect 55916 21836 55922 21888
rect 1104 21786 58880 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 58880 21786
rect 1104 21712 58880 21734
rect 1946 21672 1952 21684
rect 1907 21644 1952 21672
rect 1946 21632 1952 21644
rect 2004 21632 2010 21684
rect 2501 21675 2559 21681
rect 2501 21641 2513 21675
rect 2547 21672 2559 21675
rect 2682 21672 2688 21684
rect 2547 21644 2688 21672
rect 2547 21641 2559 21644
rect 2501 21635 2559 21641
rect 2682 21632 2688 21644
rect 2740 21632 2746 21684
rect 4798 21632 4804 21684
rect 4856 21672 4862 21684
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4856 21644 4997 21672
rect 4856 21632 4862 21644
rect 4985 21641 4997 21644
rect 5031 21672 5043 21675
rect 5442 21672 5448 21684
rect 5031 21644 5448 21672
rect 5031 21641 5043 21644
rect 4985 21635 5043 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 6730 21632 6736 21684
rect 6788 21672 6794 21684
rect 6825 21675 6883 21681
rect 6825 21672 6837 21675
rect 6788 21644 6837 21672
rect 6788 21632 6794 21644
rect 6825 21641 6837 21644
rect 6871 21641 6883 21675
rect 6825 21635 6883 21641
rect 14645 21675 14703 21681
rect 14645 21641 14657 21675
rect 14691 21672 14703 21675
rect 15838 21672 15844 21684
rect 14691 21644 15844 21672
rect 14691 21641 14703 21644
rect 14645 21635 14703 21641
rect 15838 21632 15844 21644
rect 15896 21632 15902 21684
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 16172 21644 17816 21672
rect 16172 21632 16178 21644
rect 4709 21607 4767 21613
rect 4709 21573 4721 21607
rect 4755 21604 4767 21607
rect 5994 21604 6000 21616
rect 4755 21576 6000 21604
rect 4755 21573 4767 21576
rect 4709 21567 4767 21573
rect 5994 21564 6000 21576
rect 6052 21564 6058 21616
rect 10594 21564 10600 21616
rect 10652 21604 10658 21616
rect 12434 21604 12440 21616
rect 10652 21576 12440 21604
rect 10652 21564 10658 21576
rect 3418 21536 3424 21548
rect 2700 21508 3424 21536
rect 2700 21477 2728 21508
rect 3418 21496 3424 21508
rect 3476 21496 3482 21548
rect 4062 21496 4068 21548
rect 4120 21536 4126 21548
rect 4120 21508 5488 21536
rect 4120 21496 4126 21508
rect 2685 21471 2743 21477
rect 2685 21437 2697 21471
rect 2731 21437 2743 21471
rect 2685 21431 2743 21437
rect 4709 21471 4767 21477
rect 4709 21437 4721 21471
rect 4755 21468 4767 21471
rect 4801 21471 4859 21477
rect 4801 21468 4813 21471
rect 4755 21440 4813 21468
rect 4755 21437 4767 21440
rect 4709 21431 4767 21437
rect 4801 21437 4813 21440
rect 4847 21437 4859 21471
rect 4801 21431 4859 21437
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21400 1915 21403
rect 2866 21400 2872 21412
rect 1903 21372 2872 21400
rect 1903 21369 1915 21372
rect 1857 21363 1915 21369
rect 2866 21360 2872 21372
rect 2924 21360 2930 21412
rect 3418 21400 3424 21412
rect 3379 21372 3424 21400
rect 3418 21360 3424 21372
rect 3476 21360 3482 21412
rect 3513 21403 3571 21409
rect 3513 21369 3525 21403
rect 3559 21369 3571 21403
rect 4062 21400 4068 21412
rect 4023 21372 4068 21400
rect 3513 21363 3571 21369
rect 3528 21332 3556 21363
rect 4062 21360 4068 21372
rect 4120 21360 4126 21412
rect 4798 21332 4804 21344
rect 3528 21304 4804 21332
rect 4798 21292 4804 21304
rect 4856 21292 4862 21344
rect 5460 21341 5488 21508
rect 6638 21496 6644 21548
rect 6696 21536 6702 21548
rect 7558 21536 7564 21548
rect 6696 21508 7564 21536
rect 6696 21496 6702 21508
rect 7558 21496 7564 21508
rect 7616 21536 7622 21548
rect 8202 21536 8208 21548
rect 7616 21508 8208 21536
rect 7616 21496 7622 21508
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 10796 21545 10824 21576
rect 12434 21564 12440 21576
rect 12492 21564 12498 21616
rect 13449 21607 13507 21613
rect 13449 21573 13461 21607
rect 13495 21573 13507 21607
rect 15749 21607 15807 21613
rect 15749 21604 15761 21607
rect 13449 21567 13507 21573
rect 15672 21576 15761 21604
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21536 12403 21539
rect 13464 21536 13492 21567
rect 12391 21508 13492 21536
rect 13633 21539 13691 21545
rect 12391 21505 12403 21508
rect 12345 21499 12403 21505
rect 13633 21505 13645 21539
rect 13679 21536 13691 21539
rect 13722 21536 13728 21548
rect 13679 21508 13728 21536
rect 13679 21505 13691 21508
rect 13633 21499 13691 21505
rect 13722 21496 13728 21508
rect 13780 21496 13786 21548
rect 15194 21536 15200 21548
rect 14660 21508 15200 21536
rect 5626 21468 5632 21480
rect 5587 21440 5632 21468
rect 5626 21428 5632 21440
rect 5684 21428 5690 21480
rect 6362 21428 6368 21480
rect 6420 21468 6426 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6420 21440 7021 21468
rect 6420 21428 6426 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 7760 21400 7788 21431
rect 7926 21428 7932 21480
rect 7984 21468 7990 21480
rect 8570 21468 8576 21480
rect 7984 21440 8576 21468
rect 7984 21428 7990 21440
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 8846 21477 8852 21480
rect 8840 21468 8852 21477
rect 8807 21440 8852 21468
rect 8840 21431 8852 21440
rect 8846 21428 8852 21431
rect 8904 21428 8910 21480
rect 10134 21428 10140 21480
rect 10192 21468 10198 21480
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 10192 21440 10425 21468
rect 10192 21428 10198 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21437 10655 21471
rect 10597 21431 10655 21437
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21437 10747 21471
rect 10689 21431 10747 21437
rect 7760 21372 8524 21400
rect 5445 21335 5503 21341
rect 5445 21301 5457 21335
rect 5491 21301 5503 21335
rect 7926 21332 7932 21344
rect 7887 21304 7932 21332
rect 5445 21295 5503 21301
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 8496 21332 8524 21372
rect 10318 21360 10324 21412
rect 10376 21400 10382 21412
rect 10612 21400 10640 21431
rect 10376 21372 10640 21400
rect 10704 21400 10732 21431
rect 10870 21428 10876 21480
rect 10928 21468 10934 21480
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 10928 21440 10977 21468
rect 10928 21428 10934 21440
rect 10965 21437 10977 21440
rect 11011 21437 11023 21471
rect 10965 21431 11023 21437
rect 11330 21428 11336 21480
rect 11388 21468 11394 21480
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 11388 21440 12081 21468
rect 11388 21428 11394 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 12250 21468 12256 21480
rect 12211 21440 12256 21468
rect 12069 21431 12127 21437
rect 12250 21428 12256 21440
rect 12308 21428 12314 21480
rect 12434 21468 12440 21480
rect 12395 21440 12440 21468
rect 12434 21428 12440 21440
rect 12492 21428 12498 21480
rect 12618 21468 12624 21480
rect 12579 21440 12624 21468
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 13262 21468 13268 21480
rect 13223 21440 13268 21468
rect 13262 21428 13268 21440
rect 13320 21428 13326 21480
rect 13354 21428 13360 21480
rect 13412 21468 13418 21480
rect 13412 21440 13457 21468
rect 13412 21428 13418 21440
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 13814 21468 13820 21480
rect 13596 21440 13820 21468
rect 13596 21428 13602 21440
rect 13814 21428 13820 21440
rect 13872 21428 13878 21480
rect 14660 21477 14688 21508
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 15672 21536 15700 21576
rect 15749 21573 15761 21576
rect 15795 21573 15807 21607
rect 15749 21567 15807 21573
rect 15436 21508 15700 21536
rect 17788 21536 17816 21644
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18782 21672 18788 21684
rect 18012 21644 18788 21672
rect 18012 21632 18018 21644
rect 18782 21632 18788 21644
rect 18840 21632 18846 21684
rect 19153 21675 19211 21681
rect 19153 21641 19165 21675
rect 19199 21672 19211 21675
rect 19334 21672 19340 21684
rect 19199 21644 19340 21672
rect 19199 21641 19211 21644
rect 19153 21635 19211 21641
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 21545 21675 21603 21681
rect 21545 21672 21557 21675
rect 20496 21644 21557 21672
rect 20496 21632 20502 21644
rect 21545 21641 21557 21644
rect 21591 21641 21603 21675
rect 21545 21635 21603 21641
rect 24026 21632 24032 21684
rect 24084 21672 24090 21684
rect 24213 21675 24271 21681
rect 24213 21672 24225 21675
rect 24084 21644 24225 21672
rect 24084 21632 24090 21644
rect 24213 21641 24225 21644
rect 24259 21641 24271 21675
rect 24213 21635 24271 21641
rect 24394 21632 24400 21684
rect 24452 21672 24458 21684
rect 27246 21672 27252 21684
rect 24452 21644 27252 21672
rect 24452 21632 24458 21644
rect 27246 21632 27252 21644
rect 27304 21632 27310 21684
rect 27338 21632 27344 21684
rect 27396 21672 27402 21684
rect 28994 21672 29000 21684
rect 27396 21644 29000 21672
rect 27396 21632 27402 21644
rect 28994 21632 29000 21644
rect 29052 21672 29058 21684
rect 29181 21675 29239 21681
rect 29181 21672 29193 21675
rect 29052 21644 29193 21672
rect 29052 21632 29058 21644
rect 29181 21641 29193 21644
rect 29227 21641 29239 21675
rect 29181 21635 29239 21641
rect 29825 21675 29883 21681
rect 29825 21641 29837 21675
rect 29871 21672 29883 21675
rect 30837 21675 30895 21681
rect 30837 21672 30849 21675
rect 29871 21644 30849 21672
rect 29871 21641 29883 21644
rect 29825 21635 29883 21641
rect 30837 21641 30849 21644
rect 30883 21672 30895 21675
rect 31386 21672 31392 21684
rect 30883 21644 31392 21672
rect 30883 21641 30895 21644
rect 30837 21635 30895 21641
rect 31386 21632 31392 21644
rect 31444 21632 31450 21684
rect 33137 21675 33195 21681
rect 33137 21641 33149 21675
rect 33183 21672 33195 21675
rect 33226 21672 33232 21684
rect 33183 21644 33232 21672
rect 33183 21641 33195 21644
rect 33137 21635 33195 21641
rect 33226 21632 33232 21644
rect 33284 21632 33290 21684
rect 33594 21672 33600 21684
rect 33555 21644 33600 21672
rect 33594 21632 33600 21644
rect 33652 21632 33658 21684
rect 33686 21632 33692 21684
rect 33744 21672 33750 21684
rect 35342 21672 35348 21684
rect 33744 21644 35348 21672
rect 33744 21632 33750 21644
rect 35342 21632 35348 21644
rect 35400 21672 35406 21684
rect 35529 21675 35587 21681
rect 35529 21672 35541 21675
rect 35400 21644 35541 21672
rect 35400 21632 35406 21644
rect 35529 21641 35541 21644
rect 35575 21641 35587 21675
rect 35529 21635 35587 21641
rect 55033 21675 55091 21681
rect 55033 21641 55045 21675
rect 55079 21672 55091 21675
rect 56410 21672 56416 21684
rect 55079 21644 56416 21672
rect 55079 21641 55091 21644
rect 55033 21635 55091 21641
rect 56410 21632 56416 21644
rect 56468 21632 56474 21684
rect 57974 21672 57980 21684
rect 57935 21644 57980 21672
rect 57974 21632 57980 21644
rect 58032 21632 58038 21684
rect 22554 21604 22560 21616
rect 18800 21576 22560 21604
rect 17788 21508 17908 21536
rect 15436 21496 15442 21508
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21437 14703 21471
rect 14645 21431 14703 21437
rect 14829 21471 14887 21477
rect 14829 21437 14841 21471
rect 14875 21468 14887 21471
rect 15010 21468 15016 21480
rect 14875 21440 15016 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 15010 21428 15016 21440
rect 15068 21428 15074 21480
rect 15286 21468 15292 21480
rect 15247 21440 15292 21468
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 15470 21468 15476 21480
rect 15431 21440 15476 21468
rect 15470 21428 15476 21440
rect 15528 21428 15534 21480
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 15620 21440 15665 21468
rect 15620 21428 15626 21440
rect 15838 21428 15844 21480
rect 15896 21468 15902 21480
rect 17770 21468 17776 21480
rect 15896 21440 15941 21468
rect 17731 21440 17776 21468
rect 15896 21428 15902 21440
rect 17770 21428 17776 21440
rect 17828 21428 17834 21480
rect 17880 21468 17908 21508
rect 18322 21468 18328 21480
rect 17880 21440 18328 21468
rect 18322 21428 18328 21440
rect 18380 21428 18386 21480
rect 12986 21400 12992 21412
rect 10704 21372 12992 21400
rect 10376 21360 10382 21372
rect 12986 21360 12992 21372
rect 13044 21360 13050 21412
rect 13722 21360 13728 21412
rect 13780 21400 13786 21412
rect 18018 21403 18076 21409
rect 18018 21400 18030 21403
rect 13780 21372 18030 21400
rect 13780 21360 13786 21372
rect 18018 21369 18030 21372
rect 18064 21369 18076 21403
rect 18018 21363 18076 21369
rect 9953 21335 10011 21341
rect 9953 21332 9965 21335
rect 8496 21304 9965 21332
rect 9953 21301 9965 21304
rect 9999 21332 10011 21335
rect 10502 21332 10508 21344
rect 9999 21304 10508 21332
rect 9999 21301 10011 21304
rect 9953 21295 10011 21301
rect 10502 21292 10508 21304
rect 10560 21292 10566 21344
rect 11146 21332 11152 21344
rect 11107 21304 11152 21332
rect 11146 21292 11152 21304
rect 11204 21292 11210 21344
rect 12802 21332 12808 21344
rect 12763 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 17034 21292 17040 21344
rect 17092 21332 17098 21344
rect 18800 21332 18828 21576
rect 22554 21564 22560 21576
rect 22612 21564 22618 21616
rect 25222 21564 25228 21616
rect 25280 21604 25286 21616
rect 25280 21576 30880 21604
rect 25280 21564 25286 21576
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 19702 21536 19708 21548
rect 19392 21508 19708 21536
rect 19392 21496 19398 21508
rect 19702 21496 19708 21508
rect 19760 21496 19766 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20119 21508 20668 21536
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20640 21480 20668 21508
rect 23014 21496 23020 21548
rect 23072 21536 23078 21548
rect 23293 21539 23351 21545
rect 23072 21508 23244 21536
rect 23072 21496 23078 21508
rect 19978 21477 19984 21480
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21437 19855 21471
rect 19797 21431 19855 21437
rect 19935 21471 19984 21477
rect 19935 21437 19947 21471
rect 19981 21437 19984 21471
rect 19935 21431 19984 21437
rect 19812 21400 19840 21431
rect 19978 21428 19984 21431
rect 20036 21428 20042 21480
rect 20162 21468 20168 21480
rect 20123 21440 20168 21468
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 20622 21428 20628 21480
rect 20680 21428 20686 21480
rect 20806 21468 20812 21480
rect 20767 21440 20812 21468
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21358 21428 21364 21480
rect 21416 21468 21422 21480
rect 21453 21471 21511 21477
rect 21453 21468 21465 21471
rect 21416 21440 21465 21468
rect 21416 21428 21422 21440
rect 21453 21437 21465 21440
rect 21499 21437 21511 21471
rect 22922 21468 22928 21480
rect 22883 21440 22928 21468
rect 21453 21431 21511 21437
rect 22922 21428 22928 21440
rect 22980 21428 22986 21480
rect 23106 21468 23112 21480
rect 23067 21440 23112 21468
rect 23106 21428 23112 21440
rect 23164 21428 23170 21480
rect 23216 21477 23244 21508
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23842 21536 23848 21548
rect 23339 21508 23848 21536
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 24394 21536 24400 21548
rect 24355 21508 24400 21536
rect 24394 21496 24400 21508
rect 24452 21496 24458 21548
rect 26694 21536 26700 21548
rect 26528 21508 26700 21536
rect 23204 21471 23262 21477
rect 23204 21437 23216 21471
rect 23250 21437 23262 21471
rect 23474 21468 23480 21480
rect 23435 21440 23480 21468
rect 23204 21431 23262 21437
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 24121 21471 24179 21477
rect 24121 21437 24133 21471
rect 24167 21468 24179 21471
rect 24210 21468 24216 21480
rect 24167 21440 24216 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24210 21428 24216 21440
rect 24268 21428 24274 21480
rect 25130 21468 25136 21480
rect 25091 21440 25136 21468
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 26528 21477 26556 21508
rect 26694 21496 26700 21508
rect 26752 21536 26758 21548
rect 28261 21539 28319 21545
rect 28261 21536 28273 21539
rect 26752 21508 28273 21536
rect 26752 21496 26758 21508
rect 28261 21505 28273 21508
rect 28307 21536 28319 21539
rect 30742 21536 30748 21548
rect 28307 21508 30748 21536
rect 28307 21505 28319 21508
rect 28261 21499 28319 21505
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 26513 21471 26571 21477
rect 26513 21437 26525 21471
rect 26559 21437 26571 21471
rect 26513 21431 26571 21437
rect 26605 21471 26663 21477
rect 26605 21437 26617 21471
rect 26651 21468 26663 21471
rect 26651 21440 26740 21468
rect 26651 21437 26663 21440
rect 26605 21431 26663 21437
rect 20254 21400 20260 21412
rect 19812 21372 20260 21400
rect 20254 21360 20260 21372
rect 20312 21360 20318 21412
rect 24854 21360 24860 21412
rect 24912 21400 24918 21412
rect 25317 21403 25375 21409
rect 25317 21400 25329 21403
rect 24912 21372 25329 21400
rect 24912 21360 24918 21372
rect 25317 21369 25329 21372
rect 25363 21400 25375 21403
rect 25406 21400 25412 21412
rect 25363 21372 25412 21400
rect 25363 21369 25375 21372
rect 25317 21363 25375 21369
rect 25406 21360 25412 21372
rect 25464 21360 25470 21412
rect 26712 21400 26740 21440
rect 26786 21428 26792 21480
rect 26844 21477 26850 21480
rect 26844 21471 26859 21477
rect 26847 21437 26859 21471
rect 26844 21431 26859 21437
rect 26891 21471 26949 21477
rect 26891 21437 26903 21471
rect 26937 21468 26949 21471
rect 27062 21468 27068 21480
rect 26937 21440 27068 21468
rect 26937 21437 26949 21440
rect 26891 21431 26949 21437
rect 26844 21428 26850 21431
rect 27062 21428 27068 21440
rect 27120 21428 27126 21480
rect 27614 21428 27620 21480
rect 27672 21468 27678 21480
rect 27985 21471 28043 21477
rect 27985 21468 27997 21471
rect 27672 21440 27997 21468
rect 27672 21428 27678 21440
rect 27985 21437 27997 21440
rect 28031 21437 28043 21471
rect 27985 21431 28043 21437
rect 28077 21471 28135 21477
rect 28077 21437 28089 21471
rect 28123 21437 28135 21471
rect 28077 21431 28135 21437
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21468 28411 21471
rect 28534 21468 28540 21480
rect 28399 21440 28540 21468
rect 28399 21437 28411 21440
rect 28353 21431 28411 21437
rect 26712 21372 26924 21400
rect 26896 21344 26924 21372
rect 26970 21360 26976 21412
rect 27028 21400 27034 21412
rect 27801 21403 27859 21409
rect 27801 21400 27813 21403
rect 27028 21372 27813 21400
rect 27028 21360 27034 21372
rect 27801 21369 27813 21372
rect 27847 21369 27859 21403
rect 28092 21400 28120 21431
rect 28534 21428 28540 21440
rect 28592 21428 28598 21480
rect 29086 21468 29092 21480
rect 29047 21440 29092 21468
rect 29086 21428 29092 21440
rect 29144 21428 29150 21480
rect 29733 21471 29791 21477
rect 29733 21437 29745 21471
rect 29779 21437 29791 21471
rect 30558 21468 30564 21480
rect 30519 21440 30564 21468
rect 29733 21431 29791 21437
rect 28994 21400 29000 21412
rect 28092 21372 29000 21400
rect 27801 21363 27859 21369
rect 28994 21360 29000 21372
rect 29052 21360 29058 21412
rect 29748 21400 29776 21431
rect 30558 21428 30564 21440
rect 30616 21428 30622 21480
rect 30650 21428 30656 21480
rect 30708 21468 30714 21480
rect 30708 21440 30753 21468
rect 30708 21428 30714 21440
rect 30668 21400 30696 21428
rect 29748 21372 30696 21400
rect 17092 21304 18828 21332
rect 19613 21335 19671 21341
rect 17092 21292 17098 21304
rect 19613 21301 19625 21335
rect 19659 21332 19671 21335
rect 19978 21332 19984 21344
rect 19659 21304 19984 21332
rect 19659 21301 19671 21304
rect 19613 21295 19671 21301
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 20070 21292 20076 21344
rect 20128 21332 20134 21344
rect 20901 21335 20959 21341
rect 20901 21332 20913 21335
rect 20128 21304 20913 21332
rect 20128 21292 20134 21304
rect 20901 21301 20913 21304
rect 20947 21301 20959 21335
rect 23658 21332 23664 21344
rect 23619 21304 23664 21332
rect 20901 21295 20959 21301
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 24394 21332 24400 21344
rect 24355 21304 24400 21332
rect 24394 21292 24400 21304
rect 24452 21292 24458 21344
rect 25498 21332 25504 21344
rect 25459 21304 25504 21332
rect 25498 21292 25504 21304
rect 25556 21292 25562 21344
rect 26329 21335 26387 21341
rect 26329 21301 26341 21335
rect 26375 21332 26387 21335
rect 26602 21332 26608 21344
rect 26375 21304 26608 21332
rect 26375 21301 26387 21304
rect 26329 21295 26387 21301
rect 26602 21292 26608 21304
rect 26660 21292 26666 21344
rect 26878 21292 26884 21344
rect 26936 21292 26942 21344
rect 27246 21292 27252 21344
rect 27304 21332 27310 21344
rect 29086 21332 29092 21344
rect 27304 21304 29092 21332
rect 27304 21292 27310 21304
rect 29086 21292 29092 21304
rect 29144 21292 29150 21344
rect 30374 21332 30380 21344
rect 30335 21304 30380 21332
rect 30374 21292 30380 21304
rect 30432 21292 30438 21344
rect 30852 21332 30880 21576
rect 30926 21564 30932 21616
rect 30984 21604 30990 21616
rect 30984 21576 31754 21604
rect 30984 21564 30990 21576
rect 31478 21496 31484 21548
rect 31536 21496 31542 21548
rect 31726 21536 31754 21576
rect 32214 21564 32220 21616
rect 32272 21604 32278 21616
rect 34146 21604 34152 21616
rect 32272 21576 34152 21604
rect 32272 21564 32278 21576
rect 34146 21564 34152 21576
rect 34204 21564 34210 21616
rect 56321 21607 56379 21613
rect 56321 21573 56333 21607
rect 56367 21604 56379 21607
rect 58250 21604 58256 21616
rect 56367 21576 58256 21604
rect 56367 21573 56379 21576
rect 56321 21567 56379 21573
rect 58250 21564 58256 21576
rect 58308 21564 58314 21616
rect 55858 21536 55864 21548
rect 31726 21508 34284 21536
rect 55819 21508 55864 21536
rect 30929 21471 30987 21477
rect 30929 21437 30941 21471
rect 30975 21468 30987 21471
rect 31202 21468 31208 21480
rect 30975 21440 31208 21468
rect 30975 21437 30987 21440
rect 30929 21431 30987 21437
rect 31202 21428 31208 21440
rect 31260 21468 31266 21480
rect 31496 21468 31524 21496
rect 31665 21471 31723 21477
rect 31665 21468 31677 21471
rect 31260 21440 31677 21468
rect 31260 21428 31266 21440
rect 31665 21437 31677 21440
rect 31711 21437 31723 21471
rect 33318 21468 33324 21480
rect 33279 21440 33324 21468
rect 31665 21431 31723 21437
rect 33318 21428 33324 21440
rect 33376 21428 33382 21480
rect 33413 21471 33471 21477
rect 33413 21437 33425 21471
rect 33459 21468 33471 21471
rect 33594 21468 33600 21480
rect 33459 21440 33600 21468
rect 33459 21437 33471 21440
rect 33413 21431 33471 21437
rect 33594 21428 33600 21440
rect 33652 21428 33658 21480
rect 33689 21471 33747 21477
rect 33689 21437 33701 21471
rect 33735 21468 33747 21471
rect 33870 21468 33876 21480
rect 33735 21440 33876 21468
rect 33735 21437 33747 21440
rect 33689 21431 33747 21437
rect 33870 21428 33876 21440
rect 33928 21428 33934 21480
rect 34149 21471 34207 21477
rect 34149 21437 34161 21471
rect 34195 21437 34207 21471
rect 34256 21468 34284 21508
rect 55858 21496 55864 21508
rect 55916 21496 55922 21548
rect 36078 21468 36084 21480
rect 34256 21440 34744 21468
rect 36039 21440 36084 21468
rect 34149 21431 34207 21437
rect 31478 21400 31484 21412
rect 31439 21372 31484 21400
rect 31478 21360 31484 21372
rect 31536 21360 31542 21412
rect 33042 21360 33048 21412
rect 33100 21400 33106 21412
rect 34164 21400 34192 21431
rect 34238 21400 34244 21412
rect 33100 21372 34244 21400
rect 33100 21360 33106 21372
rect 34238 21360 34244 21372
rect 34296 21360 34302 21412
rect 34416 21403 34474 21409
rect 34416 21369 34428 21403
rect 34462 21400 34474 21403
rect 34606 21400 34612 21412
rect 34462 21372 34612 21400
rect 34462 21369 34474 21372
rect 34416 21363 34474 21369
rect 34606 21360 34612 21372
rect 34664 21360 34670 21412
rect 34716 21400 34744 21440
rect 36078 21428 36084 21440
rect 36136 21428 36142 21480
rect 36265 21471 36323 21477
rect 36265 21437 36277 21471
rect 36311 21437 36323 21471
rect 36265 21431 36323 21437
rect 36280 21400 36308 21431
rect 55214 21428 55220 21480
rect 55272 21468 55278 21480
rect 55674 21468 55680 21480
rect 55272 21440 55317 21468
rect 55635 21440 55680 21468
rect 55272 21428 55278 21440
rect 55674 21428 55680 21440
rect 55732 21428 55738 21480
rect 56870 21468 56876 21480
rect 56831 21440 56876 21468
rect 56870 21428 56876 21440
rect 56928 21428 56934 21480
rect 57514 21468 57520 21480
rect 57475 21440 57520 21468
rect 57514 21428 57520 21440
rect 57572 21428 57578 21480
rect 57698 21468 57704 21480
rect 57659 21440 57704 21468
rect 57698 21428 57704 21440
rect 57756 21428 57762 21480
rect 34716 21372 36308 21400
rect 36449 21403 36507 21409
rect 36449 21369 36461 21403
rect 36495 21400 36507 21403
rect 48038 21400 48044 21412
rect 36495 21372 48044 21400
rect 36495 21369 36507 21372
rect 36449 21363 36507 21369
rect 48038 21360 48044 21372
rect 48096 21360 48102 21412
rect 33962 21332 33968 21344
rect 30852 21304 33968 21332
rect 33962 21292 33968 21304
rect 34020 21292 34026 21344
rect 34054 21292 34060 21344
rect 34112 21332 34118 21344
rect 34514 21332 34520 21344
rect 34112 21304 34520 21332
rect 34112 21292 34118 21304
rect 34514 21292 34520 21304
rect 34572 21292 34578 21344
rect 55214 21292 55220 21344
rect 55272 21332 55278 21344
rect 57057 21335 57115 21341
rect 57057 21332 57069 21335
rect 55272 21304 57069 21332
rect 55272 21292 55278 21304
rect 57057 21301 57069 21304
rect 57103 21332 57115 21335
rect 57422 21332 57428 21344
rect 57103 21304 57428 21332
rect 57103 21301 57115 21304
rect 57057 21295 57115 21301
rect 57422 21292 57428 21304
rect 57480 21292 57486 21344
rect 1104 21242 58880 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 50326 21242
rect 50378 21190 50390 21242
rect 50442 21190 50454 21242
rect 50506 21190 50518 21242
rect 50570 21190 58880 21242
rect 1104 21168 58880 21190
rect 3145 21131 3203 21137
rect 3145 21097 3157 21131
rect 3191 21128 3203 21131
rect 3510 21128 3516 21140
rect 3191 21100 3516 21128
rect 3191 21097 3203 21100
rect 3145 21091 3203 21097
rect 3510 21088 3516 21100
rect 3568 21088 3574 21140
rect 4249 21131 4307 21137
rect 4249 21097 4261 21131
rect 4295 21128 4307 21131
rect 4706 21128 4712 21140
rect 4295 21100 4712 21128
rect 4295 21097 4307 21100
rect 4249 21091 4307 21097
rect 4706 21088 4712 21100
rect 4764 21088 4770 21140
rect 4798 21088 4804 21140
rect 4856 21128 4862 21140
rect 6181 21131 6239 21137
rect 6181 21128 6193 21131
rect 4856 21100 6193 21128
rect 4856 21088 4862 21100
rect 6181 21097 6193 21100
rect 6227 21097 6239 21131
rect 8573 21131 8631 21137
rect 8573 21128 8585 21131
rect 6181 21091 6239 21097
rect 7116 21100 8585 21128
rect 1857 21063 1915 21069
rect 1857 21029 1869 21063
rect 1903 21060 1915 21063
rect 2774 21060 2780 21072
rect 1903 21032 2780 21060
rect 1903 21029 1915 21032
rect 1857 21023 1915 21029
rect 2774 21020 2780 21032
rect 2832 21020 2838 21072
rect 5626 21060 5632 21072
rect 5092 21032 5632 21060
rect 2501 20995 2559 21001
rect 2501 20961 2513 20995
rect 2547 20992 2559 20995
rect 2590 20992 2596 21004
rect 2547 20964 2596 20992
rect 2547 20961 2559 20964
rect 2501 20955 2559 20961
rect 2590 20952 2596 20964
rect 2648 20952 2654 21004
rect 2682 20952 2688 21004
rect 2740 20992 2746 21004
rect 5092 21001 5120 21032
rect 5626 21020 5632 21032
rect 5684 21020 5690 21072
rect 7116 21069 7144 21100
rect 8573 21097 8585 21100
rect 8619 21097 8631 21131
rect 15102 21128 15108 21140
rect 8573 21091 8631 21097
rect 13648 21100 15108 21128
rect 7101 21063 7159 21069
rect 7101 21029 7113 21063
rect 7147 21029 7159 21063
rect 7101 21023 7159 21029
rect 7190 21020 7196 21072
rect 7248 21060 7254 21072
rect 9760 21063 9818 21069
rect 7248 21032 7293 21060
rect 7248 21020 7254 21032
rect 9760 21029 9772 21063
rect 9806 21060 9818 21063
rect 11146 21060 11152 21072
rect 9806 21032 11152 21060
rect 9806 21029 9818 21032
rect 9760 21023 9818 21029
rect 11146 21020 11152 21032
rect 11204 21020 11210 21072
rect 11876 21063 11934 21069
rect 11876 21029 11888 21063
rect 11922 21060 11934 21063
rect 12802 21060 12808 21072
rect 11922 21032 12808 21060
rect 11922 21029 11934 21032
rect 11876 21023 11934 21029
rect 12802 21020 12808 21032
rect 12860 21020 12866 21072
rect 3329 20995 3387 21001
rect 3329 20992 3341 20995
rect 2740 20964 3341 20992
rect 2740 20952 2746 20964
rect 3329 20961 3341 20964
rect 3375 20992 3387 20995
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 3375 20964 4445 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 4433 20961 4445 20964
rect 4479 20992 4491 20995
rect 5077 20995 5135 21001
rect 5077 20992 5089 20995
rect 4479 20964 5089 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 5077 20961 5089 20964
rect 5123 20961 5135 20995
rect 5077 20955 5135 20961
rect 5442 20952 5448 21004
rect 5500 20992 5506 21004
rect 5537 20995 5595 21001
rect 5537 20992 5549 20995
rect 5500 20964 5549 20992
rect 5500 20952 5506 20964
rect 5537 20961 5549 20964
rect 5583 20961 5595 20995
rect 6362 20992 6368 21004
rect 6323 20964 6368 20992
rect 5537 20955 5595 20961
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 8202 20992 8208 21004
rect 8163 20964 8208 20992
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 8386 20992 8392 21004
rect 8347 20964 8392 20992
rect 8386 20952 8392 20964
rect 8444 20952 8450 21004
rect 8478 20952 8484 21004
rect 8536 20992 8542 21004
rect 9493 20995 9551 21001
rect 9493 20992 9505 20995
rect 8536 20964 9505 20992
rect 8536 20952 8542 20964
rect 9493 20961 9505 20964
rect 9539 20961 9551 20995
rect 11606 20992 11612 21004
rect 11567 20964 11612 20992
rect 9493 20955 9551 20961
rect 11606 20952 11612 20964
rect 11664 20952 11670 21004
rect 13648 21001 13676 21100
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 15194 21088 15200 21140
rect 15252 21128 15258 21140
rect 17586 21128 17592 21140
rect 15252 21100 17592 21128
rect 15252 21088 15258 21100
rect 17586 21088 17592 21100
rect 17644 21088 17650 21140
rect 17862 21128 17868 21140
rect 17823 21100 17868 21128
rect 17862 21088 17868 21100
rect 17920 21088 17926 21140
rect 18969 21131 19027 21137
rect 18969 21097 18981 21131
rect 19015 21128 19027 21131
rect 20070 21128 20076 21140
rect 19015 21100 20076 21128
rect 19015 21097 19027 21100
rect 18969 21091 19027 21097
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 20254 21128 20260 21140
rect 20215 21100 20260 21128
rect 20254 21088 20260 21100
rect 20312 21088 20318 21140
rect 20806 21088 20812 21140
rect 20864 21128 20870 21140
rect 22097 21131 22155 21137
rect 22097 21128 22109 21131
rect 20864 21100 22109 21128
rect 20864 21088 20870 21100
rect 22097 21097 22109 21100
rect 22143 21097 22155 21131
rect 22097 21091 22155 21097
rect 23106 21088 23112 21140
rect 23164 21128 23170 21140
rect 23164 21100 23796 21128
rect 23164 21088 23170 21100
rect 17678 21060 17684 21072
rect 13832 21032 17684 21060
rect 13832 21001 13860 21032
rect 17678 21020 17684 21032
rect 17736 21020 17742 21072
rect 20272 21060 20300 21088
rect 21542 21060 21548 21072
rect 18892 21032 20300 21060
rect 20732 21032 21548 21060
rect 13633 20995 13691 21001
rect 13633 20961 13645 20995
rect 13679 20961 13691 20995
rect 13633 20955 13691 20961
rect 13817 20995 13875 21001
rect 13817 20961 13829 20995
rect 13863 20961 13875 20995
rect 13817 20955 13875 20961
rect 14826 20952 14832 21004
rect 14884 20992 14890 21004
rect 14993 20995 15051 21001
rect 14993 20992 15005 20995
rect 14884 20964 15005 20992
rect 14884 20952 14890 20964
rect 14993 20961 15005 20964
rect 15039 20961 15051 20995
rect 14993 20955 15051 20961
rect 15470 20952 15476 21004
rect 15528 20992 15534 21004
rect 15528 20964 16988 20992
rect 15528 20952 15534 20964
rect 3786 20884 3792 20936
rect 3844 20924 3850 20936
rect 6380 20924 6408 20952
rect 7374 20924 7380 20936
rect 3844 20896 6408 20924
rect 7335 20896 7380 20924
rect 3844 20884 3850 20896
rect 7374 20884 7380 20896
rect 7432 20884 7438 20936
rect 13722 20924 13728 20936
rect 13683 20896 13728 20924
rect 13722 20884 13728 20896
rect 13780 20884 13786 20936
rect 14550 20884 14556 20936
rect 14608 20924 14614 20936
rect 14737 20927 14795 20933
rect 14737 20924 14749 20927
rect 14608 20896 14749 20924
rect 14608 20884 14614 20896
rect 14737 20893 14749 20896
rect 14783 20893 14795 20927
rect 14737 20887 14795 20893
rect 4614 20816 4620 20868
rect 4672 20856 4678 20868
rect 4893 20859 4951 20865
rect 4893 20856 4905 20859
rect 4672 20828 4905 20856
rect 4672 20816 4678 20828
rect 4893 20825 4905 20828
rect 4939 20825 4951 20859
rect 4893 20819 4951 20825
rect 1946 20788 1952 20800
rect 1907 20760 1952 20788
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 2682 20788 2688 20800
rect 2643 20760 2688 20788
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 5626 20748 5632 20800
rect 5684 20788 5690 20800
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 5684 20760 5733 20788
rect 5684 20748 5690 20760
rect 5721 20757 5733 20760
rect 5767 20757 5779 20791
rect 5721 20751 5779 20757
rect 10778 20748 10784 20800
rect 10836 20788 10842 20800
rect 10873 20791 10931 20797
rect 10873 20788 10885 20791
rect 10836 20760 10885 20788
rect 10836 20748 10842 20760
rect 10873 20757 10885 20760
rect 10919 20757 10931 20791
rect 10873 20751 10931 20757
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 12618 20788 12624 20800
rect 11020 20760 12624 20788
rect 11020 20748 11026 20760
rect 12618 20748 12624 20760
rect 12676 20788 12682 20800
rect 12989 20791 13047 20797
rect 12989 20788 13001 20791
rect 12676 20760 13001 20788
rect 12676 20748 12682 20760
rect 12989 20757 13001 20760
rect 13035 20757 13047 20791
rect 14752 20788 14780 20887
rect 16960 20856 16988 20964
rect 17034 20952 17040 21004
rect 17092 20992 17098 21004
rect 17773 20995 17831 21001
rect 17092 20964 17137 20992
rect 17092 20952 17098 20964
rect 17773 20961 17785 20995
rect 17819 20961 17831 20995
rect 17954 20992 17960 21004
rect 17915 20964 17960 20992
rect 17773 20955 17831 20961
rect 17788 20924 17816 20955
rect 17954 20952 17960 20964
rect 18012 20952 18018 21004
rect 18892 21001 18920 21032
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20961 18935 20995
rect 18877 20955 18935 20961
rect 19242 20952 19248 21004
rect 19300 20992 19306 21004
rect 20732 21001 20760 21032
rect 21542 21020 21548 21032
rect 21600 21060 21606 21072
rect 22824 21063 22882 21069
rect 21600 21032 22600 21060
rect 21600 21020 21606 21032
rect 22572 21001 22600 21032
rect 22824 21029 22836 21063
rect 22870 21060 22882 21063
rect 23658 21060 23664 21072
rect 22870 21032 23664 21060
rect 22870 21029 22882 21032
rect 22824 21023 22882 21029
rect 23658 21020 23664 21032
rect 23716 21020 23722 21072
rect 23768 21060 23796 21100
rect 23842 21088 23848 21140
rect 23900 21128 23906 21140
rect 23937 21131 23995 21137
rect 23937 21128 23949 21131
rect 23900 21100 23949 21128
rect 23900 21088 23906 21100
rect 23937 21097 23949 21100
rect 23983 21097 23995 21131
rect 25406 21128 25412 21140
rect 25367 21100 25412 21128
rect 23937 21091 23995 21097
rect 25406 21088 25412 21100
rect 25464 21088 25470 21140
rect 26145 21131 26203 21137
rect 26145 21097 26157 21131
rect 26191 21128 26203 21131
rect 31018 21128 31024 21140
rect 26191 21100 31024 21128
rect 26191 21097 26203 21100
rect 26145 21091 26203 21097
rect 31018 21088 31024 21100
rect 31076 21128 31082 21140
rect 31478 21128 31484 21140
rect 31076 21100 31484 21128
rect 31076 21088 31082 21100
rect 31478 21088 31484 21100
rect 31536 21088 31542 21140
rect 32950 21088 32956 21140
rect 33008 21128 33014 21140
rect 33873 21131 33931 21137
rect 33873 21128 33885 21131
rect 33008 21100 33885 21128
rect 33008 21088 33014 21100
rect 33873 21097 33885 21100
rect 33919 21097 33931 21131
rect 33873 21091 33931 21097
rect 34146 21088 34152 21140
rect 34204 21128 34210 21140
rect 34425 21131 34483 21137
rect 34425 21128 34437 21131
rect 34204 21100 34437 21128
rect 34204 21088 34210 21100
rect 34425 21097 34437 21100
rect 34471 21097 34483 21131
rect 55585 21131 55643 21137
rect 34425 21091 34483 21097
rect 35728 21100 36952 21128
rect 35728 21072 35756 21100
rect 28902 21060 28908 21072
rect 23768 21032 28908 21060
rect 28902 21020 28908 21032
rect 28960 21060 28966 21072
rect 30374 21060 30380 21072
rect 28960 21032 29040 21060
rect 28960 21020 28966 21032
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19300 20964 19993 20992
rect 19300 20952 19306 20964
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 20717 20995 20775 21001
rect 20717 20961 20729 20995
rect 20763 20961 20775 20995
rect 20973 20995 21031 21001
rect 20973 20992 20985 20995
rect 20717 20955 20775 20961
rect 20824 20964 20985 20992
rect 19150 20924 19156 20936
rect 17788 20896 19156 20924
rect 19150 20884 19156 20896
rect 19208 20884 19214 20936
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 20257 20927 20315 20933
rect 20257 20924 20269 20927
rect 19760 20896 20269 20924
rect 19760 20884 19766 20896
rect 20257 20893 20269 20896
rect 20303 20924 20315 20927
rect 20346 20924 20352 20936
rect 20303 20896 20352 20924
rect 20303 20893 20315 20896
rect 20257 20887 20315 20893
rect 20346 20884 20352 20896
rect 20404 20884 20410 20936
rect 20438 20884 20444 20936
rect 20496 20924 20502 20936
rect 20824 20924 20852 20964
rect 20973 20961 20985 20964
rect 21019 20961 21031 20995
rect 20973 20955 21031 20961
rect 22557 20995 22615 21001
rect 22557 20961 22569 20995
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25314 20992 25320 21004
rect 25004 20964 25320 20992
rect 25004 20952 25010 20964
rect 25314 20952 25320 20964
rect 25372 20952 25378 21004
rect 25866 20952 25872 21004
rect 25924 20992 25930 21004
rect 26375 20995 26433 21001
rect 26375 20992 26387 20995
rect 25924 20964 26387 20992
rect 25924 20952 25930 20964
rect 26375 20961 26387 20964
rect 26421 20961 26433 20995
rect 26510 20992 26516 21004
rect 26471 20964 26516 20992
rect 26375 20955 26433 20961
rect 26510 20952 26516 20964
rect 26568 20952 26574 21004
rect 26602 20952 26608 21004
rect 26660 20992 26666 21004
rect 27341 20995 27399 21001
rect 26660 20964 26705 20992
rect 26660 20952 26666 20964
rect 27341 20961 27353 20995
rect 27387 20992 27399 20995
rect 27614 20992 27620 21004
rect 27387 20964 27620 20992
rect 27387 20961 27399 20964
rect 27341 20955 27399 20961
rect 27614 20952 27620 20964
rect 27672 20952 27678 21004
rect 28169 20995 28227 21001
rect 28169 20961 28181 20995
rect 28215 20961 28227 20995
rect 28169 20955 28227 20961
rect 26878 20924 26884 20936
rect 20496 20896 20852 20924
rect 26791 20896 26884 20924
rect 20496 20884 20502 20896
rect 26878 20884 26884 20896
rect 26936 20924 26942 20936
rect 28184 20924 28212 20955
rect 28718 20952 28724 21004
rect 28776 20992 28782 21004
rect 29012 21001 29040 21032
rect 29104 21032 30380 21060
rect 29104 21001 29132 21032
rect 30374 21020 30380 21032
rect 30432 21020 30438 21072
rect 32861 21063 32919 21069
rect 32861 21029 32873 21063
rect 32907 21060 32919 21063
rect 33318 21060 33324 21072
rect 32907 21032 33324 21060
rect 32907 21029 32919 21032
rect 32861 21023 32919 21029
rect 33318 21020 33324 21032
rect 33376 21060 33382 21072
rect 33376 21032 33640 21060
rect 33376 21020 33382 21032
rect 28813 20995 28871 21001
rect 28813 20992 28825 20995
rect 28776 20964 28825 20992
rect 28776 20952 28782 20964
rect 28813 20961 28825 20964
rect 28859 20961 28871 20995
rect 28813 20955 28871 20961
rect 28997 20995 29055 21001
rect 28997 20961 29009 20995
rect 29043 20961 29055 20995
rect 28997 20955 29055 20961
rect 29089 20995 29147 21001
rect 29089 20961 29101 20995
rect 29135 20961 29147 20995
rect 29089 20955 29147 20961
rect 29270 20952 29276 21004
rect 29328 20992 29334 21004
rect 29365 20995 29423 21001
rect 29365 20992 29377 20995
rect 29328 20964 29377 20992
rect 29328 20952 29334 20964
rect 29365 20961 29377 20964
rect 29411 20961 29423 20995
rect 31202 20992 31208 21004
rect 31163 20964 31208 20992
rect 29365 20955 29423 20961
rect 31202 20952 31208 20964
rect 31260 20952 31266 21004
rect 31297 20995 31355 21001
rect 31297 20961 31309 20995
rect 31343 20992 31355 20995
rect 31386 20992 31392 21004
rect 31343 20964 31392 20992
rect 31343 20961 31355 20964
rect 31297 20955 31355 20961
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 31570 20992 31576 21004
rect 31531 20964 31576 20992
rect 31570 20952 31576 20964
rect 31628 20952 31634 21004
rect 32582 20992 32588 21004
rect 32543 20964 32588 20992
rect 32582 20952 32588 20964
rect 32640 20952 32646 21004
rect 33612 21001 33640 21032
rect 33962 21020 33968 21072
rect 34020 21060 34026 21072
rect 35710 21060 35716 21072
rect 34020 21032 35716 21060
rect 34020 21020 34026 21032
rect 35710 21020 35716 21032
rect 35768 21020 35774 21072
rect 32769 20995 32827 21001
rect 32769 20961 32781 20995
rect 32815 20961 32827 20995
rect 32769 20955 32827 20961
rect 32977 20995 33035 21001
rect 32977 20961 32989 20995
rect 33023 20992 33035 20995
rect 33597 20995 33655 21001
rect 33023 20964 33272 20992
rect 33023 20961 33035 20964
rect 32977 20955 33035 20961
rect 29181 20927 29239 20933
rect 26936 20896 27476 20924
rect 28184 20896 29040 20924
rect 26936 20884 26942 20896
rect 19794 20856 19800 20868
rect 16960 20828 19800 20856
rect 19794 20816 19800 20828
rect 19852 20816 19858 20868
rect 20070 20856 20076 20868
rect 19983 20828 20076 20856
rect 20070 20816 20076 20828
rect 20128 20856 20134 20868
rect 20714 20856 20720 20868
rect 20128 20828 20720 20856
rect 20128 20816 20134 20828
rect 20714 20816 20720 20828
rect 20772 20816 20778 20868
rect 27448 20865 27476 20896
rect 29012 20868 29040 20896
rect 29181 20893 29193 20927
rect 29227 20924 29239 20927
rect 30926 20924 30932 20936
rect 29227 20896 30932 20924
rect 29227 20893 29239 20896
rect 29181 20887 29239 20893
rect 30926 20884 30932 20896
rect 30984 20924 30990 20936
rect 32784 20924 32812 20955
rect 30984 20896 32812 20924
rect 33244 20924 33272 20964
rect 33597 20961 33609 20995
rect 33643 20961 33655 20995
rect 34330 20992 34336 21004
rect 34291 20964 34336 20992
rect 33597 20955 33655 20961
rect 34330 20952 34336 20964
rect 34388 20952 34394 21004
rect 36078 20992 36084 21004
rect 36039 20964 36084 20992
rect 36078 20952 36084 20964
rect 36136 20952 36142 21004
rect 36924 21001 36952 21100
rect 55585 21097 55597 21131
rect 55631 21128 55643 21131
rect 57698 21128 57704 21140
rect 55631 21100 57704 21128
rect 55631 21097 55643 21100
rect 55585 21091 55643 21097
rect 57698 21088 57704 21100
rect 57756 21088 57762 21140
rect 57514 21060 57520 21072
rect 55140 21032 57520 21060
rect 55140 21001 55168 21032
rect 57514 21020 57520 21032
rect 57572 21020 57578 21072
rect 36265 20995 36323 21001
rect 36265 20961 36277 20995
rect 36311 20961 36323 20995
rect 36265 20955 36323 20961
rect 36909 20995 36967 21001
rect 36909 20961 36921 20995
rect 36955 20961 36967 20995
rect 36909 20955 36967 20961
rect 55125 20995 55183 21001
rect 55125 20961 55137 20995
rect 55171 20961 55183 20995
rect 55125 20955 55183 20961
rect 33686 20924 33692 20936
rect 33244 20896 33692 20924
rect 30984 20884 30990 20896
rect 33686 20884 33692 20896
rect 33744 20884 33750 20936
rect 33873 20927 33931 20933
rect 33873 20893 33885 20927
rect 33919 20893 33931 20927
rect 33873 20887 33931 20893
rect 27433 20859 27491 20865
rect 27433 20825 27445 20859
rect 27479 20856 27491 20859
rect 28534 20856 28540 20868
rect 27479 20828 28540 20856
rect 27479 20825 27491 20828
rect 27433 20819 27491 20825
rect 28534 20816 28540 20828
rect 28592 20816 28598 20868
rect 28994 20816 29000 20868
rect 29052 20816 29058 20868
rect 31021 20859 31079 20865
rect 31021 20825 31033 20859
rect 31067 20856 31079 20859
rect 32490 20856 32496 20868
rect 31067 20828 32496 20856
rect 31067 20825 31079 20828
rect 31021 20819 31079 20825
rect 32490 20816 32496 20828
rect 32548 20816 32554 20868
rect 33137 20859 33195 20865
rect 33137 20825 33149 20859
rect 33183 20856 33195 20859
rect 33888 20856 33916 20887
rect 33962 20884 33968 20936
rect 34020 20924 34026 20936
rect 36280 20924 36308 20955
rect 55214 20952 55220 21004
rect 55272 20992 55278 21004
rect 55769 20995 55827 21001
rect 55769 20992 55781 20995
rect 55272 20964 55781 20992
rect 55272 20952 55278 20964
rect 55769 20961 55781 20964
rect 55815 20961 55827 20995
rect 55769 20955 55827 20961
rect 56042 20952 56048 21004
rect 56100 20992 56106 21004
rect 56873 20995 56931 21001
rect 56873 20992 56885 20995
rect 56100 20964 56885 20992
rect 56100 20952 56106 20964
rect 56873 20961 56885 20964
rect 56919 20961 56931 20995
rect 56873 20955 56931 20961
rect 57333 20995 57391 21001
rect 57333 20961 57345 20995
rect 57379 20992 57391 20995
rect 57977 20995 58035 21001
rect 57977 20992 57989 20995
rect 57379 20964 57989 20992
rect 57379 20961 57391 20964
rect 57333 20955 57391 20961
rect 57977 20961 57989 20964
rect 58023 20961 58035 20995
rect 58158 20992 58164 21004
rect 58119 20964 58164 20992
rect 57977 20955 58035 20961
rect 58158 20952 58164 20964
rect 58216 20952 58222 21004
rect 34020 20896 36308 20924
rect 34020 20884 34026 20896
rect 36446 20884 36452 20936
rect 36504 20924 36510 20936
rect 56597 20927 56655 20933
rect 56597 20924 56609 20927
rect 36504 20896 56609 20924
rect 36504 20884 36510 20896
rect 56597 20893 56609 20896
rect 56643 20924 56655 20927
rect 56689 20927 56747 20933
rect 56689 20924 56701 20927
rect 56643 20896 56701 20924
rect 56643 20893 56655 20896
rect 56597 20887 56655 20893
rect 56689 20893 56701 20896
rect 56735 20893 56747 20927
rect 56689 20887 56747 20893
rect 33183 20828 33916 20856
rect 36357 20859 36415 20865
rect 33183 20825 33195 20828
rect 33137 20819 33195 20825
rect 36357 20825 36369 20859
rect 36403 20856 36415 20859
rect 55674 20856 55680 20868
rect 36403 20828 41414 20856
rect 36403 20825 36415 20828
rect 36357 20819 36415 20825
rect 15470 20788 15476 20800
rect 14752 20760 15476 20788
rect 12989 20751 13047 20757
rect 15470 20748 15476 20760
rect 15528 20788 15534 20800
rect 15930 20788 15936 20800
rect 15528 20760 15936 20788
rect 15528 20748 15534 20760
rect 15930 20748 15936 20760
rect 15988 20748 15994 20800
rect 16114 20788 16120 20800
rect 16075 20760 16120 20788
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16264 20760 17141 20788
rect 16264 20748 16270 20760
rect 17129 20757 17141 20760
rect 17175 20757 17187 20791
rect 17129 20751 17187 20757
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 19702 20788 19708 20800
rect 17460 20760 19708 20788
rect 17460 20748 17466 20760
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 26694 20748 26700 20800
rect 26752 20788 26758 20800
rect 26789 20791 26847 20797
rect 26789 20788 26801 20791
rect 26752 20760 26801 20788
rect 26752 20748 26758 20760
rect 26789 20757 26801 20760
rect 26835 20788 26847 20791
rect 28261 20791 28319 20797
rect 28261 20788 28273 20791
rect 26835 20760 28273 20788
rect 26835 20757 26847 20760
rect 26789 20751 26847 20757
rect 28261 20757 28273 20760
rect 28307 20757 28319 20791
rect 28261 20751 28319 20757
rect 29549 20791 29607 20797
rect 29549 20757 29561 20791
rect 29595 20788 29607 20791
rect 29730 20788 29736 20800
rect 29595 20760 29736 20788
rect 29595 20757 29607 20760
rect 29549 20751 29607 20757
rect 29730 20748 29736 20760
rect 29788 20748 29794 20800
rect 31481 20791 31539 20797
rect 31481 20757 31493 20791
rect 31527 20788 31539 20791
rect 31938 20788 31944 20800
rect 31527 20760 31944 20788
rect 31527 20757 31539 20760
rect 31481 20751 31539 20757
rect 31938 20748 31944 20760
rect 31996 20748 32002 20800
rect 36078 20748 36084 20800
rect 36136 20788 36142 20800
rect 37093 20791 37151 20797
rect 37093 20788 37105 20791
rect 36136 20760 37105 20788
rect 36136 20748 36142 20760
rect 37093 20757 37105 20760
rect 37139 20757 37151 20791
rect 41386 20788 41414 20828
rect 45526 20828 55680 20856
rect 45526 20788 45554 20828
rect 55674 20816 55680 20828
rect 55732 20816 55738 20868
rect 41386 20760 45554 20788
rect 37093 20751 37151 20757
rect 1104 20698 58880 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 58880 20698
rect 1104 20624 58880 20646
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2038 20584 2044 20596
rect 1995 20556 2044 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 7190 20544 7196 20596
rect 7248 20584 7254 20596
rect 8021 20587 8079 20593
rect 8021 20584 8033 20587
rect 7248 20556 8033 20584
rect 7248 20544 7254 20556
rect 8021 20553 8033 20556
rect 8067 20553 8079 20587
rect 8021 20547 8079 20553
rect 10318 20544 10324 20596
rect 10376 20584 10382 20596
rect 11790 20584 11796 20596
rect 10376 20556 11796 20584
rect 10376 20544 10382 20556
rect 11790 20544 11796 20556
rect 11848 20584 11854 20596
rect 12250 20584 12256 20596
rect 11848 20556 12256 20584
rect 11848 20544 11854 20556
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 13262 20584 13268 20596
rect 13223 20556 13268 20584
rect 13262 20544 13268 20556
rect 13320 20584 13326 20596
rect 14001 20587 14059 20593
rect 14001 20584 14013 20587
rect 13320 20556 14013 20584
rect 13320 20544 13326 20556
rect 14001 20553 14013 20556
rect 14047 20584 14059 20587
rect 14090 20584 14096 20596
rect 14047 20556 14096 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 14826 20584 14832 20596
rect 14787 20556 14832 20584
rect 14826 20544 14832 20556
rect 14884 20544 14890 20596
rect 22922 20584 22928 20596
rect 14936 20556 22928 20584
rect 4433 20519 4491 20525
rect 4433 20485 4445 20519
rect 4479 20485 4491 20519
rect 4433 20479 4491 20485
rect 4448 20448 4476 20479
rect 5994 20476 6000 20528
rect 6052 20516 6058 20528
rect 13357 20519 13415 20525
rect 13357 20516 13369 20519
rect 6052 20488 8984 20516
rect 6052 20476 6058 20488
rect 5261 20451 5319 20457
rect 5261 20448 5273 20451
rect 4448 20420 5273 20448
rect 5261 20417 5273 20420
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20448 6975 20451
rect 8757 20451 8815 20457
rect 8757 20448 8769 20451
rect 6963 20420 8769 20448
rect 6963 20417 6975 20420
rect 6917 20411 6975 20417
rect 8757 20417 8769 20420
rect 8803 20417 8815 20451
rect 8757 20411 8815 20417
rect 2133 20383 2191 20389
rect 2133 20349 2145 20383
rect 2179 20380 2191 20383
rect 2682 20380 2688 20392
rect 2179 20352 2688 20380
rect 2179 20349 2191 20352
rect 2133 20343 2191 20349
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20349 4675 20383
rect 5074 20380 5080 20392
rect 5035 20352 5080 20380
rect 4617 20343 4675 20349
rect 2961 20315 3019 20321
rect 2961 20281 2973 20315
rect 3007 20281 3019 20315
rect 2961 20275 3019 20281
rect 2976 20244 3004 20275
rect 3050 20272 3056 20324
rect 3108 20312 3114 20324
rect 3602 20312 3608 20324
rect 3108 20284 3153 20312
rect 3563 20284 3608 20312
rect 3108 20272 3114 20284
rect 3602 20272 3608 20284
rect 3660 20272 3666 20324
rect 4632 20312 4660 20343
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 7668 20352 8217 20380
rect 5350 20312 5356 20324
rect 4632 20284 5356 20312
rect 5350 20272 5356 20284
rect 5408 20312 5414 20324
rect 5626 20312 5632 20324
rect 5408 20284 5632 20312
rect 5408 20272 5414 20284
rect 5626 20272 5632 20284
rect 5684 20312 5690 20324
rect 5684 20284 6960 20312
rect 5684 20272 5690 20284
rect 5442 20244 5448 20256
rect 2976 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 5534 20204 5540 20256
rect 5592 20244 5598 20256
rect 5721 20247 5779 20253
rect 5721 20244 5733 20247
rect 5592 20216 5733 20244
rect 5592 20204 5598 20216
rect 5721 20213 5733 20216
rect 5767 20213 5779 20247
rect 6932 20244 6960 20284
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 7558 20312 7564 20324
rect 7064 20284 7109 20312
rect 7519 20284 7564 20312
rect 7064 20272 7070 20284
rect 7558 20272 7564 20284
rect 7616 20272 7622 20324
rect 7668 20244 7696 20352
rect 8205 20349 8217 20352
rect 8251 20380 8263 20383
rect 8478 20380 8484 20392
rect 8251 20352 8484 20380
rect 8251 20349 8263 20352
rect 8205 20343 8263 20349
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 8665 20383 8723 20389
rect 8665 20349 8677 20383
rect 8711 20349 8723 20383
rect 8846 20380 8852 20392
rect 8807 20352 8852 20380
rect 8665 20343 8723 20349
rect 8018 20272 8024 20324
rect 8076 20312 8082 20324
rect 8680 20312 8708 20343
rect 8846 20340 8852 20352
rect 8904 20340 8910 20392
rect 8076 20284 8708 20312
rect 8956 20312 8984 20488
rect 10428 20488 13369 20516
rect 10428 20457 10456 20488
rect 13357 20485 13369 20488
rect 13403 20485 13415 20519
rect 13357 20479 13415 20485
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 14936 20516 14964 20556
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 23014 20544 23020 20596
rect 23072 20584 23078 20596
rect 23474 20584 23480 20596
rect 23072 20556 23117 20584
rect 23308 20556 23480 20584
rect 23072 20544 23078 20556
rect 13964 20488 14964 20516
rect 19061 20519 19119 20525
rect 13964 20476 13970 20488
rect 19061 20485 19073 20519
rect 19107 20485 19119 20519
rect 19061 20479 19119 20485
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 10594 20448 10600 20460
rect 10551 20420 10600 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13538 20448 13544 20460
rect 13495 20420 13544 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 13538 20408 13544 20420
rect 13596 20448 13602 20460
rect 14185 20451 14243 20457
rect 14185 20448 14197 20451
rect 13596 20420 14197 20448
rect 13596 20408 13602 20420
rect 14185 20417 14197 20420
rect 14231 20448 14243 20451
rect 14274 20448 14280 20460
rect 14231 20420 14280 20448
rect 14231 20417 14243 20420
rect 14185 20411 14243 20417
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 15286 20448 15292 20460
rect 14844 20420 15292 20448
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9493 20383 9551 20389
rect 9493 20380 9505 20383
rect 9180 20352 9505 20380
rect 9180 20340 9186 20352
rect 9493 20349 9505 20352
rect 9539 20349 9551 20383
rect 10134 20380 10140 20392
rect 10095 20352 10140 20380
rect 9493 20343 9551 20349
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 10318 20380 10324 20392
rect 10279 20352 10324 20380
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 10686 20380 10692 20392
rect 10647 20352 10692 20380
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 12066 20380 12072 20392
rect 12027 20352 12072 20380
rect 12066 20340 12072 20352
rect 12124 20340 12130 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13814 20380 13820 20392
rect 13219 20352 13820 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13814 20340 13820 20352
rect 13872 20340 13878 20392
rect 14844 20389 14872 20420
rect 15286 20408 15292 20420
rect 15344 20408 15350 20460
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16301 20451 16359 20457
rect 16301 20448 16313 20451
rect 16080 20420 16313 20448
rect 16080 20408 16086 20420
rect 16301 20417 16313 20420
rect 16347 20448 16359 20451
rect 16347 20420 17816 20448
rect 16347 20417 16359 20420
rect 16301 20411 16359 20417
rect 13909 20383 13967 20389
rect 13909 20349 13921 20383
rect 13955 20349 13967 20383
rect 13909 20343 13967 20349
rect 14829 20383 14887 20389
rect 14829 20349 14841 20383
rect 14875 20349 14887 20383
rect 15010 20380 15016 20392
rect 14971 20352 15016 20380
rect 14829 20343 14887 20349
rect 12342 20312 12348 20324
rect 8956 20284 12348 20312
rect 8076 20272 8082 20284
rect 12342 20272 12348 20284
rect 12400 20272 12406 20324
rect 13924 20312 13952 20343
rect 15010 20340 15016 20352
rect 15068 20340 15074 20392
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20380 15623 20383
rect 16114 20380 16120 20392
rect 15611 20352 16120 20380
rect 15611 20349 15623 20352
rect 15565 20343 15623 20349
rect 16114 20340 16120 20352
rect 16172 20340 16178 20392
rect 16209 20383 16267 20389
rect 16209 20349 16221 20383
rect 16255 20380 16267 20383
rect 17494 20380 17500 20392
rect 16255 20352 17500 20380
rect 16255 20349 16267 20352
rect 16209 20343 16267 20349
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 17678 20380 17684 20392
rect 17639 20352 17684 20380
rect 17678 20340 17684 20352
rect 17736 20340 17742 20392
rect 17788 20380 17816 20420
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19076 20448 19104 20479
rect 19518 20476 19524 20528
rect 19576 20516 19582 20528
rect 20990 20516 20996 20528
rect 19576 20488 20996 20516
rect 19576 20476 19582 20488
rect 20990 20476 20996 20488
rect 21048 20476 21054 20528
rect 21266 20476 21272 20528
rect 21324 20516 21330 20528
rect 23308 20516 23336 20556
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23934 20544 23940 20596
rect 23992 20584 23998 20596
rect 25406 20593 25412 20596
rect 24213 20587 24271 20593
rect 24213 20584 24225 20587
rect 23992 20556 24225 20584
rect 23992 20544 23998 20556
rect 24213 20553 24225 20556
rect 24259 20553 24271 20587
rect 24213 20547 24271 20553
rect 25390 20587 25412 20593
rect 25390 20553 25402 20587
rect 25390 20547 25412 20553
rect 25406 20544 25412 20547
rect 25464 20544 25470 20596
rect 25866 20584 25872 20596
rect 25827 20556 25872 20584
rect 25866 20544 25872 20556
rect 25924 20544 25930 20596
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 26789 20587 26847 20593
rect 26789 20584 26801 20587
rect 26568 20556 26801 20584
rect 26568 20544 26574 20556
rect 26789 20553 26801 20556
rect 26835 20553 26847 20587
rect 26789 20547 26847 20553
rect 28994 20544 29000 20596
rect 29052 20584 29058 20596
rect 29181 20587 29239 20593
rect 29181 20584 29193 20587
rect 29052 20556 29193 20584
rect 29052 20544 29058 20556
rect 29181 20553 29193 20556
rect 29227 20553 29239 20587
rect 29181 20547 29239 20553
rect 30650 20544 30656 20596
rect 30708 20584 30714 20596
rect 31481 20587 31539 20593
rect 31481 20584 31493 20587
rect 30708 20556 31493 20584
rect 30708 20544 30714 20556
rect 31481 20553 31493 20556
rect 31527 20553 31539 20587
rect 31481 20547 31539 20553
rect 33318 20544 33324 20596
rect 33376 20584 33382 20596
rect 34425 20587 34483 20593
rect 34425 20584 34437 20587
rect 33376 20556 34437 20584
rect 33376 20544 33382 20556
rect 34425 20553 34437 20556
rect 34471 20553 34483 20587
rect 34425 20547 34483 20553
rect 34606 20544 34612 20596
rect 34664 20584 34670 20596
rect 34885 20587 34943 20593
rect 34885 20584 34897 20587
rect 34664 20556 34897 20584
rect 34664 20544 34670 20556
rect 34885 20553 34897 20556
rect 34931 20553 34943 20587
rect 34885 20547 34943 20553
rect 55033 20587 55091 20593
rect 55033 20553 55045 20587
rect 55079 20584 55091 20587
rect 56042 20584 56048 20596
rect 55079 20556 56048 20584
rect 55079 20553 55091 20556
rect 55033 20547 55091 20553
rect 56042 20544 56048 20556
rect 56100 20544 56106 20596
rect 56870 20584 56876 20596
rect 56831 20556 56876 20584
rect 56870 20544 56876 20556
rect 56928 20544 56934 20596
rect 24026 20516 24032 20528
rect 21324 20488 23336 20516
rect 23492 20488 24032 20516
rect 21324 20476 21330 20488
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 18932 20420 19901 20448
rect 18932 20408 18938 20420
rect 19889 20417 19901 20420
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 19978 20408 19984 20460
rect 20036 20408 20042 20460
rect 20530 20448 20536 20460
rect 20088 20420 20536 20448
rect 18506 20380 18512 20392
rect 17788 20352 18512 20380
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 19518 20380 19524 20392
rect 19479 20352 19524 20380
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 19610 20340 19616 20392
rect 19668 20380 19674 20392
rect 19705 20383 19763 20389
rect 19705 20380 19717 20383
rect 19668 20352 19717 20380
rect 19668 20340 19674 20352
rect 19705 20349 19717 20352
rect 19751 20349 19763 20383
rect 19705 20343 19763 20349
rect 19806 20383 19864 20389
rect 19806 20349 19818 20383
rect 19852 20380 19864 20383
rect 19996 20380 20024 20408
rect 20088 20389 20116 20420
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20622 20408 20628 20460
rect 20680 20448 20686 20460
rect 21177 20451 21235 20457
rect 20680 20420 21036 20448
rect 20680 20408 20686 20420
rect 19852 20352 20024 20380
rect 20073 20383 20131 20389
rect 19852 20349 19864 20352
rect 19806 20343 19864 20349
rect 20073 20349 20085 20383
rect 20119 20349 20131 20383
rect 20073 20343 20131 20349
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20898 20380 20904 20392
rect 20220 20352 20904 20380
rect 20220 20340 20226 20352
rect 20898 20340 20904 20352
rect 20956 20340 20962 20392
rect 21008 20389 21036 20420
rect 21177 20417 21189 20451
rect 21223 20448 21235 20451
rect 21542 20448 21548 20460
rect 21223 20420 21548 20448
rect 21223 20417 21235 20420
rect 21177 20411 21235 20417
rect 21542 20408 21548 20420
rect 21600 20408 21606 20460
rect 23492 20457 23520 20488
rect 24026 20476 24032 20488
rect 24084 20516 24090 20528
rect 24489 20519 24547 20525
rect 24489 20516 24501 20519
rect 24084 20488 24501 20516
rect 24084 20476 24090 20488
rect 24489 20485 24501 20488
rect 24535 20516 24547 20519
rect 25501 20519 25559 20525
rect 25501 20516 25513 20519
rect 24535 20488 25513 20516
rect 24535 20485 24547 20488
rect 24489 20479 24547 20485
rect 25501 20485 25513 20488
rect 25547 20516 25559 20519
rect 27706 20516 27712 20528
rect 25547 20488 27712 20516
rect 25547 20485 25559 20488
rect 25501 20479 25559 20485
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 30926 20476 30932 20528
rect 30984 20516 30990 20528
rect 31021 20519 31079 20525
rect 31021 20516 31033 20519
rect 30984 20488 31033 20516
rect 30984 20476 30990 20488
rect 31021 20485 31033 20488
rect 31067 20485 31079 20519
rect 31021 20479 31079 20485
rect 23477 20451 23535 20457
rect 23477 20417 23489 20451
rect 23523 20417 23535 20451
rect 25590 20448 25596 20460
rect 23477 20411 23535 20417
rect 24412 20420 25596 20448
rect 20993 20383 21051 20389
rect 20993 20349 21005 20383
rect 21039 20349 21051 20383
rect 21269 20383 21327 20389
rect 21269 20380 21281 20383
rect 20993 20343 21051 20349
rect 21192 20352 21281 20380
rect 21192 20324 21220 20352
rect 21269 20349 21281 20352
rect 21315 20349 21327 20383
rect 21269 20343 21327 20349
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20349 23259 20383
rect 23201 20343 23259 20349
rect 17948 20315 18006 20321
rect 13924 20284 17908 20312
rect 9674 20244 9680 20256
rect 6932 20216 7696 20244
rect 9635 20216 9680 20244
rect 5721 20207 5779 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 10870 20244 10876 20256
rect 10831 20216 10876 20244
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 14182 20244 14188 20256
rect 14143 20216 14188 20244
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 15562 20204 15568 20256
rect 15620 20244 15626 20256
rect 15657 20247 15715 20253
rect 15657 20244 15669 20247
rect 15620 20216 15669 20244
rect 15620 20204 15626 20216
rect 15657 20213 15669 20216
rect 15703 20244 15715 20247
rect 15838 20244 15844 20256
rect 15703 20216 15844 20244
rect 15703 20213 15715 20216
rect 15657 20207 15715 20213
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 17880 20244 17908 20284
rect 17948 20281 17960 20315
rect 17994 20312 18006 20315
rect 20257 20315 20315 20321
rect 20257 20312 20269 20315
rect 17994 20284 20269 20312
rect 17994 20281 18006 20284
rect 17948 20275 18006 20281
rect 20257 20281 20269 20284
rect 20303 20281 20315 20315
rect 20257 20275 20315 20281
rect 21174 20272 21180 20324
rect 21232 20272 21238 20324
rect 23216 20312 23244 20343
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23566 20380 23572 20392
rect 23348 20352 23393 20380
rect 23527 20352 23572 20380
rect 23348 20340 23354 20352
rect 23566 20340 23572 20352
rect 23624 20380 23630 20392
rect 24412 20389 24440 20420
rect 25590 20408 25596 20420
rect 25648 20408 25654 20460
rect 27798 20448 27804 20460
rect 27759 20420 27804 20448
rect 27798 20408 27804 20420
rect 27856 20408 27862 20460
rect 24397 20383 24455 20389
rect 23624 20352 24348 20380
rect 23624 20340 23630 20352
rect 23658 20312 23664 20324
rect 23216 20284 23664 20312
rect 23658 20272 23664 20284
rect 23716 20272 23722 20324
rect 24320 20312 24348 20352
rect 24397 20349 24409 20383
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 24581 20383 24639 20389
rect 24581 20349 24593 20383
rect 24627 20349 24639 20383
rect 24581 20343 24639 20349
rect 24673 20383 24731 20389
rect 24673 20349 24685 20383
rect 24719 20380 24731 20383
rect 24719 20352 25452 20380
rect 24719 20349 24731 20352
rect 24673 20343 24731 20349
rect 24596 20312 24624 20343
rect 25225 20315 25283 20321
rect 25225 20312 25237 20315
rect 24320 20284 25237 20312
rect 25225 20281 25237 20284
rect 25271 20281 25283 20315
rect 25424 20312 25452 20352
rect 25498 20340 25504 20392
rect 25556 20380 25562 20392
rect 26605 20383 26663 20389
rect 26605 20380 26617 20383
rect 25556 20352 26617 20380
rect 25556 20340 25562 20352
rect 26605 20349 26617 20352
rect 26651 20349 26663 20383
rect 27816 20380 27844 20408
rect 29641 20383 29699 20389
rect 29641 20380 29653 20383
rect 27816 20352 29653 20380
rect 26605 20343 26663 20349
rect 29641 20349 29653 20352
rect 29687 20349 29699 20383
rect 29641 20343 29699 20349
rect 26418 20312 26424 20324
rect 25424 20284 26424 20312
rect 25225 20275 25283 20281
rect 20070 20244 20076 20256
rect 17880 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20622 20204 20628 20256
rect 20680 20244 20686 20256
rect 20717 20247 20775 20253
rect 20717 20244 20729 20247
rect 20680 20216 20729 20244
rect 20680 20204 20686 20216
rect 20717 20213 20729 20216
rect 20763 20213 20775 20247
rect 20717 20207 20775 20213
rect 20898 20204 20904 20256
rect 20956 20244 20962 20256
rect 21266 20244 21272 20256
rect 20956 20216 21272 20244
rect 20956 20204 20962 20216
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 22186 20204 22192 20256
rect 22244 20244 22250 20256
rect 24578 20244 24584 20256
rect 22244 20216 24584 20244
rect 22244 20204 22250 20216
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 25240 20244 25268 20275
rect 26418 20272 26424 20284
rect 26476 20272 26482 20324
rect 28068 20315 28126 20321
rect 28068 20281 28080 20315
rect 28114 20312 28126 20315
rect 29270 20312 29276 20324
rect 28114 20284 29276 20312
rect 28114 20281 28126 20284
rect 28068 20275 28126 20281
rect 29270 20272 29276 20284
rect 29328 20272 29334 20324
rect 29656 20312 29684 20343
rect 29730 20340 29736 20392
rect 29788 20380 29794 20392
rect 29897 20383 29955 20389
rect 29897 20380 29909 20383
rect 29788 20352 29909 20380
rect 29788 20340 29794 20352
rect 29897 20349 29909 20352
rect 29943 20349 29955 20383
rect 31036 20380 31064 20479
rect 31570 20408 31576 20460
rect 31628 20448 31634 20460
rect 31628 20420 31892 20448
rect 31628 20408 31634 20420
rect 31478 20380 31484 20392
rect 31036 20352 31484 20380
rect 29897 20343 29955 20349
rect 31478 20340 31484 20352
rect 31536 20380 31542 20392
rect 31665 20383 31723 20389
rect 31665 20380 31677 20383
rect 31536 20352 31677 20380
rect 31536 20340 31542 20352
rect 31665 20349 31677 20352
rect 31711 20349 31723 20383
rect 31665 20343 31723 20349
rect 31757 20383 31815 20389
rect 31757 20349 31769 20383
rect 31803 20349 31815 20383
rect 31864 20380 31892 20420
rect 31938 20408 31944 20460
rect 31996 20448 32002 20460
rect 32858 20448 32864 20460
rect 31996 20420 32864 20448
rect 31996 20408 32002 20420
rect 32858 20408 32864 20420
rect 32916 20408 32922 20460
rect 34514 20408 34520 20460
rect 34572 20448 34578 20460
rect 36446 20448 36452 20460
rect 34572 20420 35112 20448
rect 36407 20420 36452 20448
rect 34572 20408 34578 20420
rect 32033 20383 32091 20389
rect 32033 20380 32045 20383
rect 31864 20352 32045 20380
rect 31757 20343 31815 20349
rect 32033 20349 32045 20352
rect 32079 20349 32091 20383
rect 33042 20380 33048 20392
rect 33003 20352 33048 20380
rect 32033 20343 32091 20349
rect 30926 20312 30932 20324
rect 29656 20284 30932 20312
rect 30926 20272 30932 20284
rect 30984 20272 30990 20324
rect 31772 20312 31800 20343
rect 33042 20340 33048 20352
rect 33100 20340 33106 20392
rect 33134 20340 33140 20392
rect 33192 20380 33198 20392
rect 35084 20389 35112 20420
rect 36446 20408 36452 20420
rect 36504 20408 36510 20460
rect 33301 20383 33359 20389
rect 33301 20380 33313 20383
rect 33192 20352 33313 20380
rect 33192 20340 33198 20352
rect 33301 20349 33313 20352
rect 33347 20349 33359 20383
rect 33301 20343 33359 20349
rect 34885 20383 34943 20389
rect 34885 20349 34897 20383
rect 34931 20349 34943 20383
rect 34885 20343 34943 20349
rect 35069 20383 35127 20389
rect 35069 20349 35081 20383
rect 35115 20349 35127 20383
rect 36078 20380 36084 20392
rect 36039 20352 36084 20380
rect 35069 20343 35127 20349
rect 32582 20312 32588 20324
rect 31772 20284 32588 20312
rect 32582 20272 32588 20284
rect 32640 20272 32646 20324
rect 34900 20312 34928 20343
rect 36078 20340 36084 20352
rect 36136 20340 36142 20392
rect 36262 20380 36268 20392
rect 36223 20352 36268 20380
rect 36262 20340 36268 20352
rect 36320 20340 36326 20392
rect 54389 20383 54447 20389
rect 54389 20349 54401 20383
rect 54435 20349 54447 20383
rect 54389 20343 54447 20349
rect 35986 20312 35992 20324
rect 34900 20284 35992 20312
rect 26878 20244 26884 20256
rect 25240 20216 26884 20244
rect 26878 20204 26884 20216
rect 26936 20204 26942 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 29638 20244 29644 20256
rect 29420 20216 29644 20244
rect 29420 20204 29426 20216
rect 29638 20204 29644 20216
rect 29696 20244 29702 20256
rect 34900 20244 34928 20284
rect 35986 20272 35992 20284
rect 36044 20272 36050 20324
rect 54404 20312 54432 20343
rect 55214 20340 55220 20392
rect 55272 20380 55278 20392
rect 55272 20352 55317 20380
rect 55272 20340 55278 20352
rect 55398 20340 55404 20392
rect 55456 20380 55462 20392
rect 55677 20383 55735 20389
rect 55677 20380 55689 20383
rect 55456 20352 55689 20380
rect 55456 20340 55462 20352
rect 55677 20349 55689 20352
rect 55723 20380 55735 20383
rect 56042 20380 56048 20392
rect 55723 20352 56048 20380
rect 55723 20349 55735 20352
rect 55677 20343 55735 20349
rect 56042 20340 56048 20352
rect 56100 20340 56106 20392
rect 56962 20340 56968 20392
rect 57020 20380 57026 20392
rect 57517 20383 57575 20389
rect 57517 20380 57529 20383
rect 57020 20352 57529 20380
rect 57020 20340 57026 20352
rect 57517 20349 57529 20352
rect 57563 20349 57575 20383
rect 57698 20380 57704 20392
rect 57659 20352 57704 20380
rect 57517 20343 57575 20349
rect 57698 20340 57704 20352
rect 57756 20340 57762 20392
rect 56502 20312 56508 20324
rect 54404 20284 56508 20312
rect 56502 20272 56508 20284
rect 56560 20272 56566 20324
rect 56778 20312 56784 20324
rect 56739 20284 56784 20312
rect 56778 20272 56784 20284
rect 56836 20272 56842 20324
rect 29696 20216 34928 20244
rect 29696 20204 29702 20216
rect 55214 20204 55220 20256
rect 55272 20244 55278 20256
rect 55766 20244 55772 20256
rect 55272 20216 55772 20244
rect 55272 20204 55278 20216
rect 55766 20204 55772 20216
rect 55824 20244 55830 20256
rect 55861 20247 55919 20253
rect 55861 20244 55873 20247
rect 55824 20216 55873 20244
rect 55824 20204 55830 20216
rect 55861 20213 55873 20216
rect 55907 20244 55919 20247
rect 56134 20244 56140 20256
rect 55907 20216 56140 20244
rect 55907 20213 55919 20216
rect 55861 20207 55919 20213
rect 56134 20204 56140 20216
rect 56192 20204 56198 20256
rect 57974 20204 57980 20256
rect 58032 20244 58038 20256
rect 58161 20247 58219 20253
rect 58161 20244 58173 20247
rect 58032 20216 58173 20244
rect 58032 20204 58038 20216
rect 58161 20213 58173 20216
rect 58207 20213 58219 20247
rect 58161 20207 58219 20213
rect 1104 20154 58880 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 50326 20154
rect 50378 20102 50390 20154
rect 50442 20102 50454 20154
rect 50506 20102 50518 20154
rect 50570 20102 58880 20154
rect 1104 20080 58880 20102
rect 2958 20040 2964 20052
rect 1688 20012 2964 20040
rect 1688 19981 1716 20012
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 7926 20040 7932 20052
rect 4172 20012 7932 20040
rect 1673 19975 1731 19981
rect 1673 19941 1685 19975
rect 1719 19941 1731 19975
rect 2498 19972 2504 19984
rect 2459 19944 2504 19972
rect 1673 19935 1731 19941
rect 2498 19932 2504 19944
rect 2556 19932 2562 19984
rect 2409 19839 2467 19845
rect 2409 19805 2421 19839
rect 2455 19836 2467 19839
rect 4172 19836 4200 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 8297 20043 8355 20049
rect 8297 20009 8309 20043
rect 8343 20009 8355 20043
rect 12250 20040 12256 20052
rect 8297 20003 8355 20009
rect 11624 20012 12256 20040
rect 4433 19975 4491 19981
rect 4433 19941 4445 19975
rect 4479 19972 4491 19975
rect 4614 19972 4620 19984
rect 4479 19944 4620 19972
rect 4479 19941 4491 19944
rect 4433 19935 4491 19941
rect 4614 19932 4620 19944
rect 4672 19932 4678 19984
rect 7285 19975 7343 19981
rect 7285 19941 7297 19975
rect 7331 19972 7343 19975
rect 8312 19972 8340 20003
rect 7331 19944 8340 19972
rect 9760 19975 9818 19981
rect 7331 19941 7343 19944
rect 7285 19935 7343 19941
rect 9760 19941 9772 19975
rect 9806 19972 9818 19975
rect 10870 19972 10876 19984
rect 9806 19944 10876 19972
rect 9806 19941 9818 19944
rect 9760 19935 9818 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19904 5503 19907
rect 5718 19904 5724 19916
rect 5491 19876 5724 19904
rect 5491 19873 5503 19876
rect 5445 19867 5503 19873
rect 5718 19864 5724 19876
rect 5776 19864 5782 19916
rect 8478 19904 8484 19916
rect 8439 19876 8484 19904
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 8570 19864 8576 19916
rect 8628 19904 8634 19916
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 8628 19876 9505 19904
rect 8628 19864 8634 19876
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 11330 19864 11336 19916
rect 11388 19904 11394 19916
rect 11624 19913 11652 20012
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 50982 20040 50988 20052
rect 12400 20012 50988 20040
rect 12400 20000 12406 20012
rect 50982 20000 50988 20012
rect 51040 20000 51046 20052
rect 14182 19972 14188 19984
rect 11900 19944 14188 19972
rect 11609 19907 11667 19913
rect 11609 19904 11621 19907
rect 11388 19876 11621 19904
rect 11388 19864 11394 19876
rect 11609 19873 11621 19876
rect 11655 19873 11667 19907
rect 11790 19904 11796 19916
rect 11751 19876 11796 19904
rect 11609 19867 11667 19873
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 11900 19913 11928 19944
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 15841 19975 15899 19981
rect 15841 19941 15853 19975
rect 15887 19972 15899 19975
rect 16638 19975 16696 19981
rect 16638 19972 16650 19975
rect 15887 19944 16650 19972
rect 15887 19941 15899 19944
rect 15841 19935 15899 19941
rect 16638 19941 16650 19944
rect 16684 19941 16696 19975
rect 16638 19935 16696 19941
rect 18325 19975 18383 19981
rect 18325 19941 18337 19975
rect 18371 19972 18383 19975
rect 21450 19972 21456 19984
rect 18371 19944 21456 19972
rect 18371 19941 18383 19944
rect 18325 19935 18383 19941
rect 21450 19932 21456 19944
rect 21508 19932 21514 19984
rect 22186 19972 22192 19984
rect 21567 19944 22192 19972
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 11885 19867 11943 19873
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 12161 19907 12219 19913
rect 12161 19904 12173 19907
rect 12124 19876 12173 19904
rect 12124 19864 12130 19876
rect 12161 19873 12173 19876
rect 12207 19873 12219 19907
rect 12161 19867 12219 19873
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 12805 19907 12863 19913
rect 12805 19904 12817 19907
rect 12308 19876 12817 19904
rect 12308 19864 12314 19876
rect 12805 19873 12817 19876
rect 12851 19873 12863 19907
rect 12805 19867 12863 19873
rect 12989 19907 13047 19913
rect 12989 19873 13001 19907
rect 13035 19873 13047 19907
rect 13354 19904 13360 19916
rect 13315 19876 13360 19904
rect 12989 19867 13047 19873
rect 2455 19808 4200 19836
rect 4341 19839 4399 19845
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 4341 19805 4353 19839
rect 4387 19805 4399 19839
rect 4798 19836 4804 19848
rect 4759 19808 4804 19836
rect 4341 19799 4399 19805
rect 1854 19768 1860 19780
rect 1815 19740 1860 19768
rect 1854 19728 1860 19740
rect 1912 19728 1918 19780
rect 2958 19768 2964 19780
rect 2919 19740 2964 19768
rect 2958 19728 2964 19740
rect 3016 19728 3022 19780
rect 4356 19768 4384 19799
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 5626 19836 5632 19848
rect 5587 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 7193 19839 7251 19845
rect 7193 19805 7205 19839
rect 7239 19836 7251 19839
rect 7282 19836 7288 19848
rect 7239 19808 7288 19836
rect 7239 19805 7251 19808
rect 7193 19799 7251 19805
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7466 19836 7472 19848
rect 7427 19808 7472 19836
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 6362 19768 6368 19780
rect 4356 19740 6368 19768
rect 6362 19728 6368 19740
rect 6420 19728 6426 19780
rect 11808 19768 11836 19864
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19836 12035 19839
rect 12434 19836 12440 19848
rect 12023 19808 12440 19836
rect 12023 19805 12035 19808
rect 11977 19799 12035 19805
rect 12434 19796 12440 19808
rect 12492 19836 12498 19848
rect 12894 19836 12900 19848
rect 12492 19808 12900 19836
rect 12492 19796 12498 19808
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 13004 19768 13032 19867
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19904 14887 19907
rect 14918 19904 14924 19916
rect 14875 19876 14924 19904
rect 14875 19873 14887 19876
rect 14829 19867 14887 19873
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 15010 19864 15016 19916
rect 15068 19904 15074 19916
rect 15746 19904 15752 19916
rect 15068 19876 15161 19904
rect 15707 19876 15752 19904
rect 15068 19864 15074 19876
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 15933 19907 15991 19913
rect 15933 19873 15945 19907
rect 15979 19904 15991 19907
rect 16206 19904 16212 19916
rect 15979 19876 16212 19904
rect 15979 19873 15991 19876
rect 15933 19867 15991 19873
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 11808 19740 13032 19768
rect 13096 19768 13124 19799
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 15028 19836 15056 19864
rect 15948 19836 15976 19867
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19873 18291 19907
rect 18874 19904 18880 19916
rect 18835 19876 18880 19904
rect 18233 19867 18291 19873
rect 13228 19808 13273 19836
rect 15028 19808 15976 19836
rect 16393 19839 16451 19845
rect 13228 19796 13234 19808
rect 16393 19805 16405 19839
rect 16439 19805 16451 19839
rect 18248 19836 18276 19867
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 20717 19907 20775 19913
rect 20717 19873 20729 19907
rect 20763 19904 20775 19907
rect 20806 19904 20812 19916
rect 20763 19876 20812 19904
rect 20763 19873 20775 19876
rect 20717 19867 20775 19873
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 20990 19904 20996 19916
rect 20951 19876 20996 19904
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 21567 19913 21595 19944
rect 22186 19932 22192 19944
rect 22244 19932 22250 19984
rect 24118 19972 24124 19984
rect 22894 19944 24124 19972
rect 21545 19907 21603 19913
rect 21545 19873 21557 19907
rect 21591 19873 21603 19907
rect 21545 19867 21603 19873
rect 21638 19907 21696 19913
rect 21638 19873 21650 19907
rect 21684 19873 21696 19907
rect 21638 19867 21696 19873
rect 20622 19836 20628 19848
rect 18248 19808 20628 19836
rect 16393 19799 16451 19805
rect 14182 19768 14188 19780
rect 13096 19740 14188 19768
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 15470 19728 15476 19780
rect 15528 19768 15534 19780
rect 16408 19768 16436 19799
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 19978 19768 19984 19780
rect 15528 19740 16436 19768
rect 17328 19740 19984 19768
rect 15528 19728 15534 19740
rect 5810 19700 5816 19712
rect 5771 19672 5816 19700
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 10686 19660 10692 19712
rect 10744 19700 10750 19712
rect 10873 19703 10931 19709
rect 10873 19700 10885 19703
rect 10744 19672 10885 19700
rect 10744 19660 10750 19672
rect 10873 19669 10885 19672
rect 10919 19669 10931 19703
rect 10873 19663 10931 19669
rect 12345 19703 12403 19709
rect 12345 19669 12357 19703
rect 12391 19700 12403 19703
rect 12434 19700 12440 19712
rect 12391 19672 12440 19700
rect 12391 19669 12403 19672
rect 12345 19663 12403 19669
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 13538 19700 13544 19712
rect 13499 19672 13544 19700
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 14826 19700 14832 19712
rect 14787 19672 14832 19700
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 15010 19660 15016 19712
rect 15068 19700 15074 19712
rect 17328 19700 17356 19740
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 15068 19672 17356 19700
rect 17773 19703 17831 19709
rect 15068 19660 15074 19672
rect 17773 19669 17785 19703
rect 17819 19700 17831 19703
rect 18230 19700 18236 19712
rect 17819 19672 18236 19700
rect 17819 19669 17831 19672
rect 17773 19663 17831 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 18966 19700 18972 19712
rect 18927 19672 18972 19700
rect 18966 19660 18972 19672
rect 19024 19660 19030 19712
rect 19058 19660 19064 19712
rect 19116 19700 19122 19712
rect 19886 19700 19892 19712
rect 19116 19672 19892 19700
rect 19116 19660 19122 19672
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 20640 19700 20668 19796
rect 20714 19728 20720 19780
rect 20772 19768 20778 19780
rect 20813 19771 20871 19777
rect 20813 19768 20825 19771
rect 20772 19740 20825 19768
rect 20772 19728 20778 19740
rect 20813 19737 20825 19740
rect 20859 19737 20871 19771
rect 20813 19731 20871 19737
rect 20901 19771 20959 19777
rect 20901 19737 20913 19771
rect 20947 19768 20959 19771
rect 21266 19768 21272 19780
rect 20947 19740 21272 19768
rect 20947 19737 20959 19740
rect 20901 19731 20959 19737
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 21450 19728 21456 19780
rect 21508 19768 21514 19780
rect 21653 19768 21681 19867
rect 21726 19864 21732 19916
rect 21784 19913 21790 19916
rect 21784 19907 21833 19913
rect 21784 19873 21787 19907
rect 21821 19873 21833 19907
rect 21910 19904 21916 19916
rect 21871 19876 21916 19904
rect 21784 19867 21833 19873
rect 21784 19864 21790 19867
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 22894 19913 22922 19944
rect 24118 19932 24124 19944
rect 24176 19972 24182 19984
rect 24486 19972 24492 19984
rect 24176 19944 24492 19972
rect 24176 19932 24182 19944
rect 24486 19932 24492 19944
rect 24544 19932 24550 19984
rect 25593 19975 25651 19981
rect 25593 19941 25605 19975
rect 25639 19972 25651 19975
rect 26602 19972 26608 19984
rect 25639 19944 26608 19972
rect 25639 19941 25651 19944
rect 25593 19935 25651 19941
rect 26602 19932 26608 19944
rect 26660 19932 26666 19984
rect 27706 19972 27712 19984
rect 27667 19944 27712 19972
rect 27706 19932 27712 19944
rect 27764 19932 27770 19984
rect 28350 19972 28356 19984
rect 28311 19944 28356 19972
rect 28350 19932 28356 19944
rect 28408 19932 28414 19984
rect 28718 19932 28724 19984
rect 28776 19972 28782 19984
rect 36262 19972 36268 19984
rect 28776 19944 36268 19972
rect 28776 19932 28782 19944
rect 36262 19932 36268 19944
rect 36320 19932 36326 19984
rect 51000 19972 51028 20000
rect 54941 19975 54999 19981
rect 54941 19972 54953 19975
rect 51000 19944 54953 19972
rect 54941 19941 54953 19944
rect 54987 19941 54999 19975
rect 54941 19935 54999 19941
rect 55309 19975 55367 19981
rect 55309 19941 55321 19975
rect 55355 19972 55367 19975
rect 56778 19972 56784 19984
rect 55355 19944 56784 19972
rect 55355 19941 55367 19944
rect 55309 19935 55367 19941
rect 22051 19907 22109 19913
rect 22051 19873 22063 19907
rect 22097 19873 22109 19907
rect 22051 19867 22109 19873
rect 22879 19907 22937 19913
rect 22879 19873 22891 19907
rect 22925 19873 22937 19907
rect 23014 19904 23020 19916
rect 22975 19876 23020 19904
rect 22879 19867 22937 19873
rect 22066 19836 22094 19867
rect 23014 19864 23020 19876
rect 23072 19864 23078 19916
rect 23109 19907 23167 19913
rect 23109 19873 23121 19907
rect 23155 19904 23167 19907
rect 23198 19904 23204 19916
rect 23155 19876 23204 19904
rect 23155 19873 23167 19876
rect 23109 19867 23167 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 23293 19907 23351 19913
rect 23293 19873 23305 19907
rect 23339 19873 23351 19907
rect 23293 19867 23351 19873
rect 23308 19836 23336 19867
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 23937 19907 23995 19913
rect 23937 19904 23949 19907
rect 23624 19876 23949 19904
rect 23624 19864 23630 19876
rect 23937 19873 23949 19876
rect 23983 19873 23995 19907
rect 23937 19867 23995 19873
rect 24026 19864 24032 19916
rect 24084 19904 24090 19916
rect 24084 19876 24129 19904
rect 24084 19864 24090 19876
rect 24210 19864 24216 19916
rect 24268 19904 24274 19916
rect 24305 19907 24363 19913
rect 24305 19904 24317 19907
rect 24268 19876 24317 19904
rect 24268 19864 24274 19876
rect 24305 19873 24317 19876
rect 24351 19873 24363 19907
rect 24305 19867 24363 19873
rect 24578 19864 24584 19916
rect 24636 19904 24642 19916
rect 25225 19907 25283 19913
rect 25225 19904 25237 19907
rect 24636 19876 25237 19904
rect 24636 19864 24642 19876
rect 25225 19873 25237 19876
rect 25271 19873 25283 19907
rect 25225 19867 25283 19873
rect 25314 19864 25320 19916
rect 25372 19904 25378 19916
rect 25498 19904 25504 19916
rect 25372 19876 25417 19904
rect 25459 19876 25504 19904
rect 25372 19864 25378 19876
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 25690 19907 25748 19913
rect 25690 19904 25702 19907
rect 25608 19876 25702 19904
rect 21508 19740 21681 19768
rect 21836 19808 22094 19836
rect 22204 19808 23336 19836
rect 23753 19839 23811 19845
rect 21508 19728 21514 19740
rect 21836 19700 21864 19808
rect 22204 19777 22232 19808
rect 23753 19805 23765 19839
rect 23799 19836 23811 19839
rect 25130 19836 25136 19848
rect 23799 19808 25136 19836
rect 23799 19805 23811 19808
rect 23753 19799 23811 19805
rect 25130 19796 25136 19808
rect 25188 19836 25194 19848
rect 25608 19836 25636 19876
rect 25690 19873 25702 19876
rect 25736 19873 25748 19907
rect 25690 19867 25748 19873
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 26789 19907 26847 19913
rect 26789 19904 26801 19907
rect 26752 19876 26801 19904
rect 26752 19864 26758 19876
rect 26789 19873 26801 19876
rect 26835 19873 26847 19907
rect 26789 19867 26847 19873
rect 26881 19907 26939 19913
rect 26881 19873 26893 19907
rect 26927 19904 26939 19907
rect 26970 19904 26976 19916
rect 26927 19876 26976 19904
rect 26927 19873 26939 19876
rect 26881 19867 26939 19873
rect 26970 19864 26976 19876
rect 27028 19864 27034 19916
rect 27157 19907 27215 19913
rect 27157 19873 27169 19907
rect 27203 19873 27215 19907
rect 27614 19904 27620 19916
rect 27575 19876 27620 19904
rect 27157 19867 27215 19873
rect 25188 19808 25636 19836
rect 25188 19796 25194 19808
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 27062 19836 27068 19848
rect 25832 19808 27068 19836
rect 25832 19796 25838 19808
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 27172 19836 27200 19867
rect 27614 19864 27620 19876
rect 27672 19864 27678 19916
rect 28258 19904 28264 19916
rect 28219 19876 28264 19904
rect 28258 19864 28264 19876
rect 28316 19864 28322 19916
rect 28445 19907 28503 19913
rect 28445 19873 28457 19907
rect 28491 19904 28503 19907
rect 28626 19904 28632 19916
rect 28491 19876 28632 19904
rect 28491 19873 28503 19876
rect 28445 19867 28503 19873
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 28810 19864 28816 19916
rect 28868 19904 28874 19916
rect 28905 19907 28963 19913
rect 28905 19904 28917 19907
rect 28868 19876 28917 19904
rect 28868 19864 28874 19876
rect 28905 19873 28917 19876
rect 28951 19873 28963 19907
rect 28905 19867 28963 19873
rect 31018 19864 31024 19916
rect 31076 19904 31082 19916
rect 31185 19907 31243 19913
rect 31185 19904 31197 19907
rect 31076 19876 31197 19904
rect 31076 19864 31082 19876
rect 31185 19873 31197 19876
rect 31231 19873 31243 19907
rect 31185 19867 31243 19873
rect 32582 19864 32588 19916
rect 32640 19904 32646 19916
rect 32769 19907 32827 19913
rect 32769 19904 32781 19907
rect 32640 19876 32781 19904
rect 32640 19864 32646 19876
rect 32769 19873 32781 19876
rect 32815 19873 32827 19907
rect 32769 19867 32827 19873
rect 32858 19864 32864 19916
rect 32916 19904 32922 19916
rect 33962 19904 33968 19916
rect 32916 19876 33968 19904
rect 32916 19864 32922 19876
rect 33962 19864 33968 19876
rect 34020 19864 34026 19916
rect 53742 19904 53748 19916
rect 53655 19876 53748 19904
rect 53742 19864 53748 19876
rect 53800 19904 53806 19916
rect 55324 19904 55352 19935
rect 56778 19932 56784 19944
rect 56836 19932 56842 19984
rect 57974 19972 57980 19984
rect 57935 19944 57980 19972
rect 57974 19932 57980 19944
rect 58032 19932 58038 19984
rect 58158 19904 58164 19916
rect 53800 19876 55352 19904
rect 58119 19876 58164 19904
rect 53800 19864 53806 19876
rect 58158 19864 58164 19876
rect 58216 19864 58222 19916
rect 27890 19836 27896 19848
rect 27172 19808 27896 19836
rect 27890 19796 27896 19808
rect 27948 19796 27954 19848
rect 30926 19836 30932 19848
rect 30887 19808 30932 19836
rect 30926 19796 30932 19808
rect 30984 19796 30990 19848
rect 22189 19771 22247 19777
rect 22189 19737 22201 19771
rect 22235 19737 22247 19771
rect 22189 19731 22247 19737
rect 25682 19728 25688 19780
rect 25740 19768 25746 19780
rect 28997 19771 29055 19777
rect 28997 19768 29009 19771
rect 25740 19740 29009 19768
rect 25740 19728 25746 19740
rect 28997 19737 29009 19740
rect 29043 19737 29055 19771
rect 28997 19731 29055 19737
rect 32309 19771 32367 19777
rect 32309 19737 32321 19771
rect 32355 19768 32367 19771
rect 32600 19768 32628 19864
rect 54294 19836 54300 19848
rect 54255 19808 54300 19836
rect 54294 19796 54300 19808
rect 54352 19796 54358 19848
rect 56686 19836 56692 19848
rect 56647 19808 56692 19836
rect 56686 19796 56692 19808
rect 56744 19796 56750 19848
rect 56870 19836 56876 19848
rect 56831 19808 56876 19836
rect 56870 19796 56876 19808
rect 56928 19796 56934 19848
rect 32355 19740 32628 19768
rect 32355 19737 32367 19740
rect 32309 19731 32367 19737
rect 22646 19700 22652 19712
rect 20640 19672 21864 19700
rect 22607 19672 22652 19700
rect 22646 19660 22652 19672
rect 22704 19660 22710 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 24213 19703 24271 19709
rect 24213 19700 24225 19703
rect 23532 19672 24225 19700
rect 23532 19660 23538 19672
rect 24213 19669 24225 19672
rect 24259 19700 24271 19703
rect 24670 19700 24676 19712
rect 24259 19672 24676 19700
rect 24259 19669 24271 19672
rect 24213 19663 24271 19669
rect 24670 19660 24676 19672
rect 24728 19660 24734 19712
rect 25869 19703 25927 19709
rect 25869 19669 25881 19703
rect 25915 19700 25927 19703
rect 26142 19700 26148 19712
rect 25915 19672 26148 19700
rect 25915 19669 25927 19672
rect 25869 19663 25927 19669
rect 26142 19660 26148 19672
rect 26200 19660 26206 19712
rect 57333 19703 57391 19709
rect 57333 19669 57345 19703
rect 57379 19700 57391 19703
rect 57974 19700 57980 19712
rect 57379 19672 57980 19700
rect 57379 19669 57391 19672
rect 57333 19663 57391 19669
rect 57974 19660 57980 19672
rect 58032 19660 58038 19712
rect 1104 19610 58880 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 58880 19610
rect 1104 19536 58880 19558
rect 1949 19499 2007 19505
rect 1949 19465 1961 19499
rect 1995 19496 2007 19499
rect 2498 19496 2504 19508
rect 1995 19468 2504 19496
rect 1995 19465 2007 19468
rect 1949 19459 2007 19465
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 4525 19499 4583 19505
rect 4525 19465 4537 19499
rect 4571 19496 4583 19499
rect 5074 19496 5080 19508
rect 4571 19468 5080 19496
rect 4571 19465 4583 19468
rect 4525 19459 4583 19465
rect 5074 19456 5080 19468
rect 5132 19456 5138 19508
rect 6825 19499 6883 19505
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 7006 19496 7012 19508
rect 6871 19468 7012 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 13998 19496 14004 19508
rect 7668 19468 14004 19496
rect 5442 19388 5448 19440
rect 5500 19428 5506 19440
rect 7668 19428 7696 19468
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 14182 19496 14188 19508
rect 14143 19468 14188 19496
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14918 19456 14924 19508
rect 14976 19496 14982 19508
rect 15105 19499 15163 19505
rect 15105 19496 15117 19499
rect 14976 19468 15117 19496
rect 14976 19456 14982 19468
rect 15105 19465 15117 19468
rect 15151 19465 15163 19499
rect 15105 19459 15163 19465
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 17313 19499 17371 19505
rect 17313 19496 17325 19499
rect 15804 19468 17325 19496
rect 15804 19456 15810 19468
rect 17313 19465 17325 19468
rect 17359 19465 17371 19499
rect 19058 19496 19064 19508
rect 19019 19468 19064 19496
rect 17313 19459 17371 19465
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19521 19499 19579 19505
rect 19521 19465 19533 19499
rect 19567 19496 19579 19499
rect 20070 19496 20076 19508
rect 19567 19468 20076 19496
rect 19567 19465 19579 19468
rect 19521 19459 19579 19465
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19496 20223 19499
rect 20714 19496 20720 19508
rect 20211 19468 20720 19496
rect 20211 19465 20223 19468
rect 20165 19459 20223 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 20864 19468 21281 19496
rect 20864 19456 20870 19468
rect 21269 19465 21281 19468
rect 21315 19496 21327 19499
rect 21726 19496 21732 19508
rect 21315 19468 21732 19496
rect 21315 19465 21327 19468
rect 21269 19459 21327 19465
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 23290 19456 23296 19508
rect 23348 19496 23354 19508
rect 24213 19499 24271 19505
rect 24213 19496 24225 19499
rect 23348 19468 24225 19496
rect 23348 19456 23354 19468
rect 24213 19465 24225 19468
rect 24259 19465 24271 19499
rect 24670 19496 24676 19508
rect 24631 19468 24676 19496
rect 24213 19459 24271 19465
rect 14090 19428 14096 19440
rect 5500 19400 7696 19428
rect 14051 19400 14096 19428
rect 5500 19388 5506 19400
rect 14090 19388 14096 19400
rect 14148 19388 14154 19440
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 16117 19431 16175 19437
rect 15436 19400 15608 19428
rect 15436 19388 15442 19400
rect 9674 19320 9680 19372
rect 9732 19360 9738 19372
rect 9769 19363 9827 19369
rect 9769 19360 9781 19363
rect 9732 19332 9781 19360
rect 9732 19320 9738 19332
rect 9769 19329 9781 19332
rect 9815 19360 9827 19363
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 9815 19332 10609 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 10597 19329 10609 19332
rect 10643 19329 10655 19363
rect 14274 19360 14280 19372
rect 14235 19332 14280 19360
rect 10597 19323 10655 19329
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 15580 19369 15608 19400
rect 16117 19397 16129 19431
rect 16163 19428 16175 19431
rect 20438 19428 20444 19440
rect 16163 19400 20444 19428
rect 16163 19397 16175 19400
rect 16117 19391 16175 19397
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 24228 19428 24256 19459
rect 24670 19456 24676 19468
rect 24728 19456 24734 19508
rect 25498 19456 25504 19508
rect 25556 19496 25562 19508
rect 26697 19499 26755 19505
rect 26697 19496 26709 19499
rect 25556 19468 26709 19496
rect 25556 19456 25562 19468
rect 26697 19465 26709 19468
rect 26743 19465 26755 19499
rect 26697 19459 26755 19465
rect 27062 19456 27068 19508
rect 27120 19496 27126 19508
rect 28718 19496 28724 19508
rect 27120 19468 28724 19496
rect 27120 19456 27126 19468
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 29914 19496 29920 19508
rect 29875 19468 29920 19496
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 30926 19456 30932 19508
rect 30984 19496 30990 19508
rect 33042 19496 33048 19508
rect 30984 19468 33048 19496
rect 30984 19456 30990 19468
rect 33042 19456 33048 19468
rect 33100 19456 33106 19508
rect 56781 19499 56839 19505
rect 56781 19465 56793 19499
rect 56827 19496 56839 19499
rect 56962 19496 56968 19508
rect 56827 19468 56968 19496
rect 56827 19465 56839 19468
rect 56781 19459 56839 19465
rect 56962 19456 56968 19468
rect 57020 19456 57026 19508
rect 57241 19499 57299 19505
rect 57241 19465 57253 19499
rect 57287 19496 57299 19499
rect 57698 19496 57704 19508
rect 57287 19468 57704 19496
rect 57287 19465 57299 19468
rect 57241 19459 57299 19465
rect 57698 19456 57704 19468
rect 57756 19456 57762 19508
rect 27614 19428 27620 19440
rect 24228 19400 27620 19428
rect 27614 19388 27620 19400
rect 27672 19388 27678 19440
rect 15565 19363 15623 19369
rect 15120 19332 15516 19360
rect 2133 19295 2191 19301
rect 2133 19261 2145 19295
rect 2179 19261 2191 19295
rect 2590 19292 2596 19304
rect 2551 19264 2596 19292
rect 2133 19255 2191 19261
rect 2148 19224 2176 19255
rect 2590 19252 2596 19264
rect 2648 19252 2654 19304
rect 3786 19292 3792 19304
rect 3747 19264 3792 19292
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19261 4583 19295
rect 4706 19292 4712 19304
rect 4667 19264 4712 19292
rect 4525 19255 4583 19261
rect 3142 19224 3148 19236
rect 2148 19196 3148 19224
rect 2792 19165 2820 19196
rect 3142 19184 3148 19196
rect 3200 19224 3206 19236
rect 3804 19224 3832 19252
rect 3200 19196 3832 19224
rect 4540 19224 4568 19255
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 5350 19292 5356 19304
rect 5311 19264 5356 19292
rect 5350 19252 5356 19264
rect 5408 19292 5414 19304
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 5408 19264 7021 19292
rect 5408 19252 5414 19264
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19261 10011 19295
rect 10778 19292 10784 19304
rect 10739 19264 10784 19292
rect 9953 19255 10011 19261
rect 5258 19224 5264 19236
rect 4540 19196 5264 19224
rect 3200 19184 3206 19196
rect 5258 19184 5264 19196
rect 5316 19184 5322 19236
rect 7929 19227 7987 19233
rect 7929 19193 7941 19227
rect 7975 19193 7987 19227
rect 7929 19187 7987 19193
rect 2777 19159 2835 19165
rect 2777 19125 2789 19159
rect 2823 19156 2835 19159
rect 3605 19159 3663 19165
rect 2823 19128 2857 19156
rect 2823 19125 2835 19128
rect 2777 19119 2835 19125
rect 3605 19125 3617 19159
rect 3651 19156 3663 19159
rect 4522 19156 4528 19168
rect 3651 19128 4528 19156
rect 3651 19125 3663 19128
rect 3605 19119 3663 19125
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 5169 19159 5227 19165
rect 5169 19125 5181 19159
rect 5215 19156 5227 19159
rect 5626 19156 5632 19168
rect 5215 19128 5632 19156
rect 5215 19125 5227 19128
rect 5169 19119 5227 19125
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 7944 19156 7972 19187
rect 8018 19184 8024 19236
rect 8076 19224 8082 19236
rect 8938 19224 8944 19236
rect 8076 19196 8121 19224
rect 8899 19196 8944 19224
rect 8076 19184 8082 19196
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 9968 19224 9996 19255
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 11146 19252 11152 19304
rect 11204 19292 11210 19304
rect 11606 19292 11612 19304
rect 11204 19264 11612 19292
rect 11204 19252 11210 19264
rect 11606 19252 11612 19264
rect 11664 19292 11670 19304
rect 12158 19292 12164 19304
rect 11664 19264 12164 19292
rect 11664 19252 11670 19264
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12434 19301 12440 19304
rect 12428 19255 12440 19301
rect 12492 19292 12498 19304
rect 14001 19295 14059 19301
rect 12492 19264 12528 19292
rect 12434 19252 12440 19255
rect 12492 19252 12498 19264
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 15010 19292 15016 19304
rect 14047 19264 15016 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 12066 19224 12072 19236
rect 9968 19196 12072 19224
rect 12066 19184 12072 19196
rect 12124 19224 12130 19236
rect 12124 19196 12434 19224
rect 12124 19184 12130 19196
rect 10042 19156 10048 19168
rect 7944 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10134 19116 10140 19168
rect 10192 19156 10198 19168
rect 10192 19128 10237 19156
rect 10192 19116 10198 19128
rect 10502 19116 10508 19168
rect 10560 19156 10566 19168
rect 10965 19159 11023 19165
rect 10965 19156 10977 19159
rect 10560 19128 10977 19156
rect 10560 19116 10566 19128
rect 10965 19125 10977 19128
rect 11011 19125 11023 19159
rect 12406 19156 12434 19196
rect 12986 19184 12992 19236
rect 13044 19224 13050 19236
rect 15120 19224 15148 19332
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19261 15439 19295
rect 15488 19292 15516 19332
rect 15565 19329 15577 19363
rect 15611 19360 15623 19363
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 15611 19332 16773 19360
rect 15611 19329 15623 19332
rect 15565 19323 15623 19329
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 17420 19332 17632 19360
rect 15657 19295 15715 19301
rect 15657 19292 15669 19295
rect 15488 19264 15669 19292
rect 15381 19255 15439 19261
rect 13044 19196 15148 19224
rect 13044 19184 13050 19196
rect 13541 19159 13599 19165
rect 13541 19156 13553 19159
rect 12406 19128 13553 19156
rect 10965 19119 11023 19125
rect 13541 19125 13553 19128
rect 13587 19125 13599 19159
rect 15396 19156 15424 19255
rect 15580 19224 15608 19264
rect 15657 19261 15669 19264
rect 15703 19261 15715 19295
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 15657 19255 15715 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16301 19295 16359 19301
rect 16301 19261 16313 19295
rect 16347 19292 16359 19295
rect 16390 19292 16396 19304
rect 16347 19264 16396 19292
rect 16347 19261 16359 19264
rect 16301 19255 16359 19261
rect 16390 19252 16396 19264
rect 16448 19252 16454 19304
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 17420 19292 17448 19332
rect 17604 19301 17632 19332
rect 17678 19320 17684 19372
rect 17736 19360 17742 19372
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17736 19332 17785 19360
rect 17736 19320 17742 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 18800 19332 20208 19360
rect 16540 19264 17448 19292
rect 17497 19295 17555 19301
rect 16540 19252 16546 19264
rect 17497 19261 17509 19295
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 17589 19295 17647 19301
rect 17589 19261 17601 19295
rect 17635 19261 17647 19295
rect 17862 19292 17868 19304
rect 17823 19264 17868 19292
rect 17589 19255 17647 19261
rect 16666 19224 16672 19236
rect 15580 19196 16672 19224
rect 16666 19184 16672 19196
rect 16724 19184 16730 19236
rect 17512 19224 17540 19255
rect 17862 19252 17868 19264
rect 17920 19252 17926 19304
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19292 18567 19295
rect 18800 19292 18828 19332
rect 18555 19264 18828 19292
rect 18555 19261 18567 19264
rect 18509 19255 18567 19261
rect 18874 19252 18880 19304
rect 18932 19292 18938 19304
rect 19245 19295 19303 19301
rect 19245 19292 19257 19295
rect 18932 19264 19257 19292
rect 18932 19252 18938 19264
rect 19245 19261 19257 19264
rect 19291 19261 19303 19295
rect 19245 19255 19303 19261
rect 19334 19252 19340 19304
rect 19392 19301 19398 19304
rect 19392 19295 19425 19301
rect 19413 19261 19425 19295
rect 19392 19255 19425 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 19392 19252 19398 19255
rect 19518 19224 19524 19236
rect 17512 19196 19524 19224
rect 19518 19184 19524 19196
rect 19576 19184 19582 19236
rect 16482 19156 16488 19168
rect 15396 19128 16488 19156
rect 13541 19119 13599 19125
rect 16482 19116 16488 19128
rect 16540 19116 16546 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17678 19156 17684 19168
rect 16807 19128 17684 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 19150 19156 19156 19168
rect 19024 19128 19156 19156
rect 19024 19116 19030 19128
rect 19150 19116 19156 19128
rect 19208 19156 19214 19168
rect 19628 19156 19656 19255
rect 19886 19252 19892 19304
rect 19944 19292 19950 19304
rect 20073 19295 20131 19301
rect 20073 19292 20085 19295
rect 19944 19264 20085 19292
rect 19944 19252 19950 19264
rect 20073 19261 20085 19264
rect 20119 19261 20131 19295
rect 20180 19292 20208 19332
rect 24210 19320 24216 19372
rect 24268 19360 24274 19372
rect 26970 19360 26976 19372
rect 24268 19332 24624 19360
rect 24268 19320 24274 19332
rect 20898 19292 20904 19304
rect 20180 19264 20904 19292
rect 20073 19255 20131 19261
rect 20898 19252 20904 19264
rect 20956 19252 20962 19304
rect 21177 19295 21235 19301
rect 21177 19261 21189 19295
rect 21223 19292 21235 19295
rect 21450 19292 21456 19304
rect 21223 19264 21456 19292
rect 21223 19261 21235 19264
rect 21177 19255 21235 19261
rect 21450 19252 21456 19264
rect 21508 19292 21514 19304
rect 21910 19292 21916 19304
rect 21508 19264 21916 19292
rect 21508 19252 21514 19264
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23017 19295 23075 19301
rect 23017 19292 23029 19295
rect 22888 19264 23029 19292
rect 22888 19252 22894 19264
rect 23017 19261 23029 19264
rect 23063 19261 23075 19295
rect 23474 19292 23480 19304
rect 23435 19264 23480 19292
rect 23017 19255 23075 19261
rect 23474 19252 23480 19264
rect 23532 19252 23538 19304
rect 23842 19252 23848 19304
rect 23900 19292 23906 19304
rect 24397 19295 24455 19301
rect 24397 19292 24409 19295
rect 23900 19264 24409 19292
rect 23900 19252 23906 19264
rect 23750 19224 23756 19236
rect 23711 19196 23756 19224
rect 23750 19184 23756 19196
rect 23808 19184 23814 19236
rect 21174 19156 21180 19168
rect 19208 19128 21180 19156
rect 19208 19116 19214 19128
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 24320 19156 24348 19264
rect 24397 19261 24409 19264
rect 24443 19261 24455 19295
rect 24397 19255 24455 19261
rect 24489 19295 24547 19301
rect 24489 19261 24501 19295
rect 24535 19261 24547 19295
rect 24596 19292 24624 19332
rect 26497 19332 26976 19360
rect 24765 19295 24823 19301
rect 24765 19292 24777 19295
rect 24596 19264 24777 19292
rect 24489 19255 24547 19261
rect 24765 19261 24777 19264
rect 24811 19261 24823 19295
rect 24765 19255 24823 19261
rect 25593 19295 25651 19301
rect 25593 19261 25605 19295
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 25961 19295 26019 19301
rect 25961 19261 25973 19295
rect 26007 19292 26019 19295
rect 26497 19292 26525 19332
rect 26970 19320 26976 19332
rect 27028 19320 27034 19372
rect 27154 19320 27160 19372
rect 27212 19360 27218 19372
rect 27212 19332 27936 19360
rect 27212 19320 27218 19332
rect 26602 19292 26608 19304
rect 26007 19264 26525 19292
rect 26563 19264 26608 19292
rect 26007 19261 26019 19264
rect 25961 19255 26019 19261
rect 24504 19224 24532 19255
rect 24670 19224 24676 19236
rect 24504 19196 24676 19224
rect 24670 19184 24676 19196
rect 24728 19224 24734 19236
rect 25608 19224 25636 19255
rect 26602 19252 26608 19264
rect 26660 19252 26666 19304
rect 26694 19252 26700 19304
rect 26752 19292 26758 19304
rect 27801 19295 27859 19301
rect 27801 19292 27813 19295
rect 26752 19264 27813 19292
rect 26752 19252 26758 19264
rect 27801 19261 27813 19264
rect 27847 19261 27859 19295
rect 27908 19292 27936 19332
rect 28552 19332 29040 19360
rect 28552 19292 28580 19332
rect 27908 19264 28580 19292
rect 28629 19295 28687 19301
rect 27801 19255 27859 19261
rect 28629 19261 28641 19295
rect 28675 19292 28687 19295
rect 28902 19292 28908 19304
rect 28675 19264 28908 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 24728 19196 25636 19224
rect 25777 19227 25835 19233
rect 24728 19184 24734 19196
rect 25777 19193 25789 19227
rect 25823 19193 25835 19227
rect 25777 19187 25835 19193
rect 25869 19227 25927 19233
rect 25869 19193 25881 19227
rect 25915 19224 25927 19227
rect 26712 19224 26740 19252
rect 25915 19196 26740 19224
rect 25915 19193 25927 19196
rect 25869 19187 25927 19193
rect 25792 19156 25820 19187
rect 26970 19184 26976 19236
rect 27028 19224 27034 19236
rect 28644 19224 28672 19255
rect 28902 19252 28908 19264
rect 28960 19252 28966 19304
rect 27028 19196 28672 19224
rect 29012 19224 29040 19332
rect 29086 19252 29092 19304
rect 29144 19292 29150 19304
rect 29273 19295 29331 19301
rect 29273 19292 29285 19295
rect 29144 19264 29285 19292
rect 29144 19252 29150 19264
rect 29273 19261 29285 19264
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 29365 19295 29423 19301
rect 29365 19261 29377 19295
rect 29411 19292 29423 19295
rect 29546 19292 29552 19304
rect 29411 19264 29552 19292
rect 29411 19261 29423 19264
rect 29365 19255 29423 19261
rect 29546 19252 29552 19264
rect 29604 19252 29610 19304
rect 29822 19252 29828 19304
rect 29880 19292 29886 19304
rect 29917 19295 29975 19301
rect 29917 19292 29929 19295
rect 29880 19264 29929 19292
rect 29880 19252 29886 19264
rect 29917 19261 29929 19264
rect 29963 19261 29975 19295
rect 29917 19255 29975 19261
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19261 30159 19295
rect 30101 19255 30159 19261
rect 30653 19295 30711 19301
rect 30653 19261 30665 19295
rect 30699 19292 30711 19295
rect 31202 19292 31208 19304
rect 30699 19264 31208 19292
rect 30699 19261 30711 19264
rect 30653 19255 30711 19261
rect 30116 19224 30144 19255
rect 31202 19252 31208 19264
rect 31260 19252 31266 19304
rect 31478 19292 31484 19304
rect 31439 19264 31484 19292
rect 31478 19252 31484 19264
rect 31536 19252 31542 19304
rect 56134 19292 56140 19304
rect 56095 19264 56140 19292
rect 56134 19252 56140 19264
rect 56192 19252 56198 19304
rect 57422 19292 57428 19304
rect 57383 19264 57428 19292
rect 57422 19252 57428 19264
rect 57480 19252 57486 19304
rect 57974 19292 57980 19304
rect 57935 19264 57980 19292
rect 57974 19252 57980 19264
rect 58032 19252 58038 19304
rect 58158 19292 58164 19304
rect 58119 19264 58164 19292
rect 58158 19252 58164 19264
rect 58216 19252 58222 19304
rect 29012 19196 30144 19224
rect 27028 19184 27034 19196
rect 30558 19184 30564 19236
rect 30616 19224 30622 19236
rect 30745 19227 30803 19233
rect 30745 19224 30757 19227
rect 30616 19196 30757 19224
rect 30616 19184 30622 19196
rect 30745 19193 30757 19196
rect 30791 19193 30803 19227
rect 30745 19187 30803 19193
rect 24320 19128 25820 19156
rect 26145 19159 26203 19165
rect 26145 19125 26157 19159
rect 26191 19156 26203 19159
rect 26510 19156 26516 19168
rect 26191 19128 26516 19156
rect 26191 19125 26203 19128
rect 26145 19119 26203 19125
rect 26510 19116 26516 19128
rect 26568 19116 26574 19168
rect 27890 19156 27896 19168
rect 27803 19128 27896 19156
rect 27890 19116 27896 19128
rect 27948 19156 27954 19168
rect 28626 19156 28632 19168
rect 27948 19128 28632 19156
rect 27948 19116 27954 19128
rect 28626 19116 28632 19128
rect 28684 19116 28690 19168
rect 31110 19116 31116 19168
rect 31168 19156 31174 19168
rect 31570 19156 31576 19168
rect 31168 19128 31576 19156
rect 31168 19116 31174 19128
rect 31570 19116 31576 19128
rect 31628 19116 31634 19168
rect 55953 19159 56011 19165
rect 55953 19125 55965 19159
rect 55999 19156 56011 19159
rect 56870 19156 56876 19168
rect 55999 19128 56876 19156
rect 55999 19125 56011 19128
rect 55953 19119 56011 19125
rect 56870 19116 56876 19128
rect 56928 19116 56934 19168
rect 1104 19066 58880 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 50326 19066
rect 50378 19014 50390 19066
rect 50442 19014 50454 19066
rect 50506 19014 50518 19066
rect 50570 19014 58880 19066
rect 1104 18992 58880 19014
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 3050 18952 3056 18964
rect 2915 18924 3056 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 3050 18912 3056 18924
rect 3108 18912 3114 18964
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 5813 18955 5871 18961
rect 5813 18952 5825 18955
rect 4764 18924 5825 18952
rect 4764 18912 4770 18924
rect 5813 18921 5825 18924
rect 5859 18921 5871 18955
rect 6362 18952 6368 18964
rect 6323 18924 6368 18952
rect 5813 18915 5871 18921
rect 2038 18884 2044 18896
rect 1999 18856 2044 18884
rect 2038 18844 2044 18856
rect 2096 18844 2102 18896
rect 5828 18884 5856 18915
rect 6362 18912 6368 18924
rect 6420 18912 6426 18964
rect 6914 18912 6920 18964
rect 6972 18952 6978 18964
rect 7009 18955 7067 18961
rect 7009 18952 7021 18955
rect 6972 18924 7021 18952
rect 6972 18912 6978 18924
rect 7009 18921 7021 18924
rect 7055 18921 7067 18955
rect 7009 18915 7067 18921
rect 7745 18955 7803 18961
rect 7745 18921 7757 18955
rect 7791 18952 7803 18955
rect 8018 18952 8024 18964
rect 7791 18924 8024 18952
rect 7791 18921 7803 18924
rect 7745 18915 7803 18921
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 10042 18912 10048 18964
rect 10100 18952 10106 18964
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 10100 18924 10241 18952
rect 10100 18912 10106 18924
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 12434 18952 12440 18964
rect 10229 18915 10287 18921
rect 10336 18924 12440 18952
rect 5902 18884 5908 18896
rect 5815 18856 5908 18884
rect 5902 18844 5908 18856
rect 5960 18884 5966 18896
rect 8846 18884 8852 18896
rect 5960 18856 8852 18884
rect 5960 18844 5966 18856
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2130 18816 2136 18828
rect 1903 18788 2136 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 3142 18816 3148 18828
rect 3099 18788 3148 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 3142 18776 3148 18788
rect 3200 18776 3206 18828
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18816 5687 18819
rect 6086 18816 6092 18828
rect 5675 18788 6092 18816
rect 5675 18785 5687 18788
rect 5629 18779 5687 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6270 18816 6276 18828
rect 6231 18788 6276 18816
rect 6270 18776 6276 18788
rect 6328 18776 6334 18828
rect 6472 18825 6500 18856
rect 6457 18819 6515 18825
rect 6457 18785 6469 18819
rect 6503 18785 6515 18819
rect 6457 18779 6515 18785
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 7006 18816 7012 18828
rect 6963 18788 7012 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7116 18825 7144 18856
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 10336 18884 10364 18924
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 13354 18952 13360 18964
rect 12584 18924 13360 18952
rect 12584 18912 12590 18924
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 16117 18955 16175 18961
rect 13504 18924 16068 18952
rect 13504 18912 13510 18924
rect 9968 18856 10364 18884
rect 11416 18887 11474 18893
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 7561 18819 7619 18825
rect 7561 18785 7573 18819
rect 7607 18816 7619 18819
rect 8110 18816 8116 18828
rect 7607 18788 8116 18816
rect 7607 18785 7619 18788
rect 7561 18779 7619 18785
rect 8110 18776 8116 18788
rect 8168 18816 8174 18828
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 8168 18788 8217 18816
rect 8168 18776 8174 18788
rect 8205 18785 8217 18788
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9861 18819 9919 18825
rect 9861 18816 9873 18819
rect 9732 18788 9873 18816
rect 9732 18776 9738 18788
rect 9861 18785 9873 18788
rect 9907 18785 9919 18819
rect 9861 18779 9919 18785
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 9968 18748 9996 18856
rect 11416 18853 11428 18887
rect 11462 18884 11474 18887
rect 13538 18884 13544 18896
rect 11462 18856 13544 18884
rect 11462 18853 11474 18856
rect 11416 18847 11474 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 14826 18844 14832 18896
rect 14884 18884 14890 18896
rect 14982 18887 15040 18893
rect 14982 18884 14994 18887
rect 14884 18856 14994 18884
rect 14884 18844 14890 18856
rect 14982 18853 14994 18856
rect 15028 18853 15040 18887
rect 14982 18847 15040 18853
rect 15194 18844 15200 18896
rect 15252 18884 15258 18896
rect 15470 18884 15476 18896
rect 15252 18856 15476 18884
rect 15252 18844 15258 18856
rect 15470 18844 15476 18856
rect 15528 18844 15534 18896
rect 10045 18819 10103 18825
rect 10045 18785 10057 18819
rect 10091 18816 10103 18819
rect 12986 18816 12992 18828
rect 10091 18788 12434 18816
rect 12947 18788 12992 18816
rect 10091 18785 10103 18788
rect 10045 18779 10103 18785
rect 11146 18748 11152 18760
rect 3476 18720 9996 18748
rect 11107 18720 11152 18748
rect 3476 18708 3482 18720
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 12406 18680 12434 18788
rect 12986 18776 12992 18788
rect 13044 18776 13050 18828
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13630 18816 13636 18828
rect 13219 18788 13492 18816
rect 13591 18788 13636 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 12526 18680 12532 18692
rect 12406 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 12894 18640 12900 18692
rect 12952 18680 12958 18692
rect 13354 18680 13360 18692
rect 12952 18652 13360 18680
rect 12952 18640 12958 18652
rect 13354 18640 13360 18652
rect 13412 18640 13418 18692
rect 13464 18680 13492 18788
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18816 14795 18819
rect 15212 18816 15240 18844
rect 14783 18788 15240 18816
rect 14783 18785 14795 18788
rect 14737 18779 14795 18785
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 15344 18788 15976 18816
rect 15344 18776 15350 18788
rect 13464 18652 13860 18680
rect 13832 18624 13860 18652
rect 8389 18615 8447 18621
rect 8389 18581 8401 18615
rect 8435 18612 8447 18615
rect 8478 18612 8484 18624
rect 8435 18584 8484 18612
rect 8435 18581 8447 18584
rect 8389 18575 8447 18581
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 12986 18612 12992 18624
rect 12947 18584 12992 18612
rect 12986 18572 12992 18584
rect 13044 18572 13050 18624
rect 13814 18612 13820 18624
rect 13727 18584 13820 18612
rect 13814 18572 13820 18584
rect 13872 18612 13878 18624
rect 14918 18612 14924 18624
rect 13872 18584 14924 18612
rect 13872 18572 13878 18584
rect 14918 18572 14924 18584
rect 14976 18572 14982 18624
rect 15948 18612 15976 18788
rect 16040 18748 16068 18924
rect 16117 18921 16129 18955
rect 16163 18921 16175 18955
rect 16666 18952 16672 18964
rect 16627 18924 16672 18952
rect 16117 18915 16175 18921
rect 16132 18884 16160 18915
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 19061 18955 19119 18961
rect 19061 18921 19073 18955
rect 19107 18952 19119 18955
rect 19334 18952 19340 18964
rect 19107 18924 19340 18952
rect 19107 18921 19119 18924
rect 19061 18915 19119 18921
rect 19334 18912 19340 18924
rect 19392 18952 19398 18964
rect 20070 18952 20076 18964
rect 19392 18924 19932 18952
rect 20031 18924 20076 18952
rect 19392 18912 19398 18924
rect 16132 18856 16344 18884
rect 16316 18816 16344 18856
rect 16390 18844 16396 18896
rect 16448 18884 16454 18896
rect 19242 18884 19248 18896
rect 16448 18856 19248 18884
rect 16448 18844 16454 18856
rect 19242 18844 19248 18856
rect 19300 18844 19306 18896
rect 16577 18819 16635 18825
rect 16577 18816 16589 18819
rect 16316 18788 16589 18816
rect 16577 18785 16589 18788
rect 16623 18785 16635 18819
rect 16577 18779 16635 18785
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 17770 18816 17776 18828
rect 17727 18788 17776 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 17770 18776 17776 18788
rect 17828 18776 17834 18828
rect 17948 18819 18006 18825
rect 17948 18785 17960 18819
rect 17994 18816 18006 18819
rect 18966 18816 18972 18828
rect 17994 18788 18972 18816
rect 17994 18785 18006 18788
rect 17948 18779 18006 18785
rect 18966 18776 18972 18788
rect 19024 18776 19030 18828
rect 19904 18816 19932 18924
rect 20070 18912 20076 18924
rect 20128 18912 20134 18964
rect 20625 18955 20683 18961
rect 20625 18921 20637 18955
rect 20671 18952 20683 18955
rect 20990 18952 20996 18964
rect 20671 18924 20996 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 28902 18952 28908 18964
rect 28863 18924 28908 18952
rect 28902 18912 28908 18924
rect 28960 18912 28966 18964
rect 29178 18912 29184 18964
rect 29236 18952 29242 18964
rect 29457 18955 29515 18961
rect 29457 18952 29469 18955
rect 29236 18924 29469 18952
rect 29236 18912 29242 18924
rect 29457 18921 29469 18924
rect 29503 18921 29515 18955
rect 31018 18952 31024 18964
rect 30979 18924 31024 18952
rect 29457 18915 29515 18921
rect 31018 18912 31024 18924
rect 31076 18912 31082 18964
rect 22272 18887 22330 18893
rect 20088 18856 22094 18884
rect 19981 18819 20039 18825
rect 19981 18816 19993 18819
rect 19904 18788 19993 18816
rect 19981 18785 19993 18788
rect 20027 18785 20039 18819
rect 19981 18779 20039 18785
rect 16850 18748 16856 18760
rect 16040 18720 16856 18748
rect 16850 18708 16856 18720
rect 16908 18708 16914 18760
rect 20088 18748 20116 18856
rect 20809 18819 20867 18825
rect 20809 18785 20821 18819
rect 20855 18816 20867 18819
rect 21174 18816 21180 18828
rect 20855 18788 21180 18816
rect 20855 18785 20867 18788
rect 20809 18779 20867 18785
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 21269 18819 21327 18825
rect 21269 18785 21281 18819
rect 21315 18816 21327 18819
rect 21910 18816 21916 18828
rect 21315 18788 21916 18816
rect 21315 18785 21327 18788
rect 21269 18779 21327 18785
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 22066 18816 22094 18856
rect 22272 18853 22284 18887
rect 22318 18884 22330 18887
rect 22646 18884 22652 18896
rect 22318 18856 22652 18884
rect 22318 18853 22330 18856
rect 22272 18847 22330 18853
rect 22646 18844 22652 18856
rect 22704 18844 22710 18896
rect 23750 18844 23756 18896
rect 23808 18884 23814 18896
rect 56686 18884 56692 18896
rect 23808 18856 56692 18884
rect 23808 18844 23814 18856
rect 56686 18844 56692 18856
rect 56744 18844 56750 18896
rect 23474 18816 23480 18828
rect 22066 18788 23480 18816
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 23842 18776 23848 18828
rect 23900 18816 23906 18828
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23900 18788 24041 18816
rect 23900 18776 23906 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24029 18779 24087 18785
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 25731 18819 25789 18825
rect 25731 18816 25743 18819
rect 24176 18788 25743 18816
rect 24176 18776 24182 18788
rect 25731 18785 25743 18788
rect 25777 18785 25789 18819
rect 25731 18779 25789 18785
rect 25850 18819 25908 18825
rect 25850 18785 25862 18819
rect 25896 18816 25908 18819
rect 25896 18785 25912 18816
rect 25850 18779 25912 18785
rect 20990 18748 20996 18760
rect 19996 18720 20116 18748
rect 20951 18720 20996 18748
rect 19996 18612 20024 18720
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21634 18748 21640 18760
rect 21131 18720 21640 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 22002 18748 22008 18760
rect 21744 18720 22008 18748
rect 20070 18640 20076 18692
rect 20128 18680 20134 18692
rect 20901 18683 20959 18689
rect 20901 18680 20913 18683
rect 20128 18652 20913 18680
rect 20128 18640 20134 18652
rect 20901 18649 20913 18652
rect 20947 18680 20959 18683
rect 21542 18680 21548 18692
rect 20947 18652 21548 18680
rect 20947 18649 20959 18652
rect 20901 18643 20959 18649
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 15948 18584 20024 18612
rect 20254 18572 20260 18624
rect 20312 18612 20318 18624
rect 21744 18612 21772 18720
rect 22002 18708 22008 18720
rect 22060 18708 22066 18760
rect 25884 18748 25912 18779
rect 25958 18776 25964 18828
rect 26016 18825 26022 18828
rect 26016 18819 26040 18825
rect 26028 18785 26040 18819
rect 26142 18816 26148 18828
rect 26103 18788 26148 18816
rect 26016 18779 26040 18785
rect 26016 18776 26022 18779
rect 26142 18776 26148 18788
rect 26200 18776 26206 18828
rect 26602 18816 26608 18828
rect 26252 18788 26608 18816
rect 26252 18748 26280 18788
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 26697 18819 26755 18825
rect 26697 18785 26709 18819
rect 26743 18816 26755 18819
rect 26970 18816 26976 18828
rect 26743 18788 26976 18816
rect 26743 18785 26755 18788
rect 26697 18779 26755 18785
rect 26970 18776 26976 18788
rect 27028 18776 27034 18828
rect 27792 18819 27850 18825
rect 27792 18785 27804 18819
rect 27838 18816 27850 18819
rect 28350 18816 28356 18828
rect 27838 18788 28356 18816
rect 27838 18785 27850 18788
rect 27792 18779 27850 18785
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 29362 18816 29368 18828
rect 29323 18788 29368 18816
rect 29362 18776 29368 18788
rect 29420 18776 29426 18828
rect 29549 18819 29607 18825
rect 29549 18785 29561 18819
rect 29595 18816 29607 18819
rect 30466 18816 30472 18828
rect 29595 18788 30472 18816
rect 29595 18785 29607 18788
rect 29549 18779 29607 18785
rect 30466 18776 30472 18788
rect 30524 18776 30530 18828
rect 30926 18816 30932 18828
rect 30887 18788 30932 18816
rect 30926 18776 30932 18788
rect 30984 18776 30990 18828
rect 31110 18816 31116 18828
rect 31071 18788 31116 18816
rect 31110 18776 31116 18788
rect 31168 18776 31174 18828
rect 55582 18816 55588 18828
rect 55543 18788 55588 18816
rect 55582 18776 55588 18788
rect 55640 18776 55646 18828
rect 57974 18816 57980 18828
rect 57935 18788 57980 18816
rect 57974 18776 57980 18788
rect 58032 18776 58038 18828
rect 25884 18720 26280 18748
rect 26510 18708 26516 18760
rect 26568 18748 26574 18760
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26568 18720 26893 18748
rect 26568 18708 26574 18720
rect 26881 18717 26893 18720
rect 26927 18717 26939 18751
rect 26881 18711 26939 18717
rect 27525 18751 27583 18757
rect 27525 18717 27537 18751
rect 27571 18717 27583 18751
rect 27525 18711 27583 18717
rect 26142 18640 26148 18692
rect 26200 18680 26206 18692
rect 27540 18680 27568 18711
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 31938 18748 31944 18760
rect 28776 18720 31944 18748
rect 28776 18708 28782 18720
rect 31938 18708 31944 18720
rect 31996 18708 32002 18760
rect 58158 18680 58164 18692
rect 26200 18652 27568 18680
rect 58119 18652 58164 18680
rect 26200 18640 26206 18652
rect 58158 18640 58164 18652
rect 58216 18640 58222 18692
rect 20312 18584 21772 18612
rect 20312 18572 20318 18584
rect 21818 18572 21824 18624
rect 21876 18612 21882 18624
rect 23014 18612 23020 18624
rect 21876 18584 23020 18612
rect 21876 18572 21882 18584
rect 23014 18572 23020 18584
rect 23072 18612 23078 18624
rect 23385 18615 23443 18621
rect 23385 18612 23397 18615
rect 23072 18584 23397 18612
rect 23072 18572 23078 18584
rect 23385 18581 23397 18584
rect 23431 18581 23443 18615
rect 23385 18575 23443 18581
rect 24121 18615 24179 18621
rect 24121 18581 24133 18615
rect 24167 18612 24179 18615
rect 24210 18612 24216 18624
rect 24167 18584 24216 18612
rect 24167 18581 24179 18584
rect 24121 18575 24179 18581
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 25498 18612 25504 18624
rect 25459 18584 25504 18612
rect 25498 18572 25504 18584
rect 25556 18572 25562 18624
rect 26418 18572 26424 18624
rect 26476 18612 26482 18624
rect 26789 18615 26847 18621
rect 26789 18612 26801 18615
rect 26476 18584 26801 18612
rect 26476 18572 26482 18584
rect 26789 18581 26801 18584
rect 26835 18581 26847 18615
rect 26789 18575 26847 18581
rect 57425 18615 57483 18621
rect 57425 18581 57437 18615
rect 57471 18612 57483 18615
rect 57514 18612 57520 18624
rect 57471 18584 57520 18612
rect 57471 18581 57483 18584
rect 57425 18575 57483 18581
rect 57514 18572 57520 18584
rect 57572 18572 57578 18624
rect 1104 18522 58880 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 58880 18522
rect 1104 18448 58880 18470
rect 5718 18408 5724 18420
rect 5679 18380 5724 18408
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 12434 18408 12440 18420
rect 6144 18380 12440 18408
rect 6144 18368 6150 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12526 18368 12532 18420
rect 12584 18408 12590 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 12584 18380 16129 18408
rect 12584 18368 12590 18380
rect 16117 18377 16129 18380
rect 16163 18377 16175 18411
rect 16117 18371 16175 18377
rect 16758 18368 16764 18420
rect 16816 18408 16822 18420
rect 17313 18411 17371 18417
rect 17313 18408 17325 18411
rect 16816 18380 17325 18408
rect 16816 18368 16822 18380
rect 17313 18377 17325 18380
rect 17359 18377 17371 18411
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 17313 18371 17371 18377
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 21358 18408 21364 18420
rect 21284 18380 21364 18408
rect 12250 18300 12256 18352
rect 12308 18300 12314 18352
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 13630 18340 13636 18352
rect 12676 18312 13636 18340
rect 12676 18300 12682 18312
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 15562 18340 15568 18352
rect 14568 18312 15568 18340
rect 6178 18272 6184 18284
rect 5736 18244 6184 18272
rect 5736 18213 5764 18244
rect 6178 18232 6184 18244
rect 6236 18232 6242 18284
rect 7834 18232 7840 18284
rect 7892 18272 7898 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 7892 18244 8677 18272
rect 7892 18232 7898 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9732 18244 9965 18272
rect 9732 18232 9738 18244
rect 9953 18241 9965 18244
rect 9999 18272 10011 18275
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 9999 18244 10793 18272
rect 9999 18241 10011 18244
rect 9953 18235 10011 18241
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 5721 18207 5779 18213
rect 5721 18173 5733 18207
rect 5767 18173 5779 18207
rect 5902 18204 5908 18216
rect 5863 18176 5908 18204
rect 5721 18167 5779 18173
rect 5902 18164 5908 18176
rect 5960 18164 5966 18216
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10686 18204 10692 18216
rect 10183 18176 10692 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10686 18164 10692 18176
rect 10744 18164 10750 18216
rect 10962 18204 10968 18216
rect 10923 18176 10968 18204
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 12268 18204 12296 18300
rect 13814 18272 13820 18284
rect 13188 18244 13820 18272
rect 12333 18207 12391 18213
rect 12333 18204 12345 18207
rect 12268 18176 12345 18204
rect 12333 18173 12345 18176
rect 12379 18173 12391 18207
rect 12333 18167 12391 18173
rect 12529 18207 12587 18213
rect 12529 18173 12541 18207
rect 12575 18204 12587 18207
rect 12894 18204 12900 18216
rect 12575 18176 12900 18204
rect 12575 18173 12587 18176
rect 12529 18167 12587 18173
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13188 18213 13216 18244
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18173 13047 18207
rect 12989 18167 13047 18173
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18105 8447 18139
rect 8389 18099 8447 18105
rect 8404 18068 8432 18099
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 12434 18136 12440 18148
rect 8536 18108 8581 18136
rect 12395 18108 12440 18136
rect 8536 18096 8542 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 10134 18068 10140 18080
rect 8404 18040 10140 18068
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10318 18068 10324 18080
rect 10279 18040 10324 18068
rect 10318 18028 10324 18040
rect 10376 18028 10382 18080
rect 11149 18071 11207 18077
rect 11149 18037 11161 18071
rect 11195 18068 11207 18071
rect 11238 18068 11244 18080
rect 11195 18040 11244 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 13004 18068 13032 18167
rect 13081 18139 13139 18145
rect 13081 18105 13093 18139
rect 13127 18136 13139 18139
rect 13725 18139 13783 18145
rect 13725 18136 13737 18139
rect 13127 18108 13737 18136
rect 13127 18105 13139 18108
rect 13081 18099 13139 18105
rect 13725 18105 13737 18108
rect 13771 18105 13783 18139
rect 13725 18099 13783 18105
rect 13817 18139 13875 18145
rect 13817 18105 13829 18139
rect 13863 18136 13875 18139
rect 13906 18136 13912 18148
rect 13863 18108 13912 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 14568 18136 14596 18312
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 18414 18300 18420 18352
rect 18472 18340 18478 18352
rect 21284 18340 21312 18380
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 26053 18411 26111 18417
rect 23716 18380 25636 18408
rect 23716 18368 23722 18380
rect 21450 18340 21456 18352
rect 18472 18312 21312 18340
rect 21411 18312 21456 18340
rect 18472 18300 18478 18312
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 22002 18300 22008 18352
rect 22060 18340 22066 18352
rect 25608 18340 25636 18380
rect 26053 18377 26065 18411
rect 26099 18408 26111 18411
rect 26326 18408 26332 18420
rect 26099 18380 26332 18408
rect 26099 18377 26111 18380
rect 26053 18371 26111 18377
rect 26326 18368 26332 18380
rect 26384 18368 26390 18420
rect 28350 18368 28356 18420
rect 28408 18408 28414 18420
rect 28445 18411 28503 18417
rect 28445 18408 28457 18411
rect 28408 18380 28457 18408
rect 28408 18368 28414 18380
rect 28445 18377 28457 18380
rect 28491 18377 28503 18411
rect 29270 18408 29276 18420
rect 29231 18380 29276 18408
rect 28445 18371 28503 18377
rect 29270 18368 29276 18380
rect 29328 18368 29334 18420
rect 57974 18408 57980 18420
rect 57935 18380 57980 18408
rect 57974 18368 57980 18380
rect 58032 18368 58038 18420
rect 27893 18343 27951 18349
rect 27893 18340 27905 18343
rect 22060 18312 23980 18340
rect 25608 18312 27905 18340
rect 22060 18300 22066 18312
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 14976 18244 16344 18272
rect 14976 18232 14982 18244
rect 15396 18213 15424 18244
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 14108 18108 14596 18136
rect 14108 18068 14136 18108
rect 14642 18096 14648 18148
rect 14700 18136 14706 18148
rect 14737 18139 14795 18145
rect 14737 18136 14749 18139
rect 14700 18108 14749 18136
rect 14700 18096 14706 18108
rect 14737 18105 14749 18108
rect 14783 18105 14795 18139
rect 15212 18136 15240 18167
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16316 18213 16344 18244
rect 17770 18232 17776 18284
rect 17828 18272 17834 18284
rect 19978 18272 19984 18284
rect 17828 18244 19984 18272
rect 17828 18232 17834 18244
rect 19978 18232 19984 18244
rect 20036 18272 20042 18284
rect 20254 18272 20260 18284
rect 20036 18244 20260 18272
rect 20036 18232 20042 18244
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 20993 18275 21051 18281
rect 20993 18272 21005 18275
rect 20364 18244 21005 18272
rect 16117 18207 16175 18213
rect 16117 18204 16129 18207
rect 16080 18176 16129 18204
rect 16080 18164 16086 18176
rect 16117 18173 16129 18176
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 16301 18207 16359 18213
rect 16301 18173 16313 18207
rect 16347 18173 16359 18207
rect 17310 18204 17316 18216
rect 17271 18176 17316 18204
rect 16301 18167 16359 18173
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18204 17555 18207
rect 17954 18204 17960 18216
rect 17543 18176 17960 18204
rect 17543 18173 17555 18176
rect 17497 18167 17555 18173
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18230 18164 18236 18216
rect 18288 18204 18294 18216
rect 18325 18207 18383 18213
rect 18325 18204 18337 18207
rect 18288 18176 18337 18204
rect 18288 18164 18294 18176
rect 18325 18173 18337 18176
rect 18371 18173 18383 18207
rect 18325 18167 18383 18173
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18173 19027 18207
rect 19150 18204 19156 18216
rect 19111 18176 19156 18204
rect 18969 18167 19027 18173
rect 17862 18136 17868 18148
rect 15212 18108 17868 18136
rect 14737 18099 14795 18105
rect 17862 18096 17868 18108
rect 17920 18136 17926 18148
rect 18417 18139 18475 18145
rect 18417 18136 18429 18139
rect 17920 18108 18429 18136
rect 17920 18096 17926 18108
rect 18417 18105 18429 18108
rect 18463 18105 18475 18139
rect 18417 18099 18475 18105
rect 18984 18136 19012 18167
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 20364 18213 20392 18244
rect 20993 18241 21005 18244
rect 21039 18272 21051 18275
rect 21358 18272 21364 18284
rect 21039 18244 21364 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21358 18232 21364 18244
rect 21416 18232 21422 18284
rect 21818 18272 21824 18284
rect 21468 18244 21824 18272
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 20349 18207 20407 18213
rect 19935 18176 20300 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 19720 18136 19748 18167
rect 18984 18108 19748 18136
rect 13004 18040 14136 18068
rect 14182 18028 14188 18080
rect 14240 18068 14246 18080
rect 15289 18071 15347 18077
rect 15289 18068 15301 18071
rect 14240 18040 15301 18068
rect 14240 18028 14246 18040
rect 15289 18037 15301 18040
rect 15335 18037 15347 18071
rect 15289 18031 15347 18037
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18984 18068 19012 18108
rect 16172 18040 19012 18068
rect 19797 18071 19855 18077
rect 16172 18028 16178 18040
rect 19797 18037 19809 18071
rect 19843 18068 19855 18071
rect 20162 18068 20168 18080
rect 19843 18040 20168 18068
rect 19843 18037 19855 18040
rect 19797 18031 19855 18037
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20272 18068 20300 18176
rect 20349 18173 20361 18207
rect 20395 18173 20407 18207
rect 20349 18167 20407 18173
rect 20533 18207 20591 18213
rect 20533 18173 20545 18207
rect 20579 18204 20591 18207
rect 21177 18207 21235 18213
rect 21177 18204 21189 18207
rect 20579 18176 21189 18204
rect 20579 18173 20591 18176
rect 20533 18167 20591 18173
rect 21177 18173 21189 18176
rect 21223 18204 21235 18207
rect 21468 18204 21496 18244
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 23382 18272 23388 18284
rect 23343 18244 23388 18272
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 21223 18176 21496 18204
rect 21545 18207 21603 18213
rect 21223 18173 21235 18176
rect 21177 18167 21235 18173
rect 21545 18173 21557 18207
rect 21591 18173 21603 18207
rect 22830 18204 22836 18216
rect 22791 18176 22836 18204
rect 21545 18167 21603 18173
rect 20441 18139 20499 18145
rect 20441 18105 20453 18139
rect 20487 18136 20499 18139
rect 20990 18136 20996 18148
rect 20487 18108 20996 18136
rect 20487 18105 20499 18108
rect 20441 18099 20499 18105
rect 20990 18096 20996 18108
rect 21048 18136 21054 18148
rect 21560 18136 21588 18167
rect 22830 18164 22836 18176
rect 22888 18164 22894 18216
rect 23952 18213 23980 18312
rect 27893 18309 27905 18312
rect 27939 18309 27951 18343
rect 27893 18303 27951 18309
rect 56873 18343 56931 18349
rect 56873 18309 56885 18343
rect 56919 18340 56931 18343
rect 56919 18312 57744 18340
rect 56919 18309 56931 18312
rect 56873 18303 56931 18309
rect 26142 18272 26148 18284
rect 24964 18244 26148 18272
rect 23201 18207 23259 18213
rect 23201 18173 23213 18207
rect 23247 18173 23259 18207
rect 23201 18167 23259 18173
rect 23937 18207 23995 18213
rect 23937 18173 23949 18207
rect 23983 18204 23995 18207
rect 24964 18204 24992 18244
rect 26142 18232 26148 18244
rect 26200 18232 26206 18284
rect 28534 18232 28540 18284
rect 28592 18272 28598 18284
rect 57514 18272 57520 18284
rect 28592 18244 29500 18272
rect 57475 18244 57520 18272
rect 28592 18232 28598 18244
rect 26050 18204 26056 18216
rect 23983 18176 24992 18204
rect 26011 18176 26056 18204
rect 23983 18173 23995 18176
rect 23937 18167 23995 18173
rect 21048 18108 21588 18136
rect 21048 18096 21054 18108
rect 21634 18096 21640 18148
rect 21692 18136 21698 18148
rect 23216 18136 23244 18167
rect 26050 18164 26056 18176
rect 26108 18164 26114 18216
rect 26237 18207 26295 18213
rect 26237 18173 26249 18207
rect 26283 18204 26295 18207
rect 26786 18204 26792 18216
rect 26283 18176 26792 18204
rect 26283 18173 26295 18176
rect 26237 18167 26295 18173
rect 26786 18164 26792 18176
rect 26844 18164 26850 18216
rect 26878 18164 26884 18216
rect 26936 18204 26942 18216
rect 27801 18207 27859 18213
rect 27801 18204 27813 18207
rect 26936 18176 27813 18204
rect 26936 18164 26942 18176
rect 27801 18173 27813 18176
rect 27847 18173 27859 18207
rect 27801 18167 27859 18173
rect 28445 18207 28503 18213
rect 28445 18173 28457 18207
rect 28491 18173 28503 18207
rect 28626 18204 28632 18216
rect 28587 18176 28632 18204
rect 28445 18167 28503 18173
rect 21692 18108 23244 18136
rect 24204 18139 24262 18145
rect 21692 18096 21698 18108
rect 24204 18105 24216 18139
rect 24250 18136 24262 18139
rect 24762 18136 24768 18148
rect 24250 18108 24768 18136
rect 24250 18105 24262 18108
rect 24204 18099 24262 18105
rect 24762 18096 24768 18108
rect 24820 18096 24826 18148
rect 25774 18096 25780 18148
rect 25832 18136 25838 18148
rect 26068 18136 26096 18164
rect 28460 18136 28488 18167
rect 28626 18164 28632 18176
rect 28684 18164 28690 18216
rect 29472 18213 29500 18244
rect 57514 18232 57520 18244
rect 57572 18232 57578 18284
rect 57716 18281 57744 18312
rect 57701 18275 57759 18281
rect 57701 18241 57713 18275
rect 57747 18241 57759 18275
rect 57701 18235 57759 18241
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18173 29331 18207
rect 29273 18167 29331 18173
rect 29457 18207 29515 18213
rect 29457 18173 29469 18207
rect 29503 18173 29515 18207
rect 56226 18204 56232 18216
rect 56187 18176 56232 18204
rect 29457 18167 29515 18173
rect 29288 18136 29316 18167
rect 56226 18164 56232 18176
rect 56284 18164 56290 18216
rect 57054 18204 57060 18216
rect 56967 18176 57060 18204
rect 57054 18164 57060 18176
rect 57112 18204 57118 18216
rect 57422 18204 57428 18216
rect 57112 18176 57428 18204
rect 57112 18164 57118 18176
rect 57422 18164 57428 18176
rect 57480 18164 57486 18216
rect 30926 18136 30932 18148
rect 25832 18108 30932 18136
rect 25832 18096 25838 18108
rect 30926 18096 30932 18108
rect 30984 18096 30990 18148
rect 21910 18068 21916 18080
rect 20272 18040 21916 18068
rect 21910 18028 21916 18040
rect 21968 18028 21974 18080
rect 24026 18028 24032 18080
rect 24084 18068 24090 18080
rect 24670 18068 24676 18080
rect 24084 18040 24676 18068
rect 24084 18028 24090 18040
rect 24670 18028 24676 18040
rect 24728 18068 24734 18080
rect 25317 18071 25375 18077
rect 25317 18068 25329 18071
rect 24728 18040 25329 18068
rect 24728 18028 24734 18040
rect 25317 18037 25329 18040
rect 25363 18037 25375 18071
rect 25317 18031 25375 18037
rect 1104 17978 58880 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 50326 17978
rect 50378 17926 50390 17978
rect 50442 17926 50454 17978
rect 50506 17926 50518 17978
rect 50570 17926 58880 17978
rect 1104 17904 58880 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 13998 17824 14004 17876
rect 14056 17864 14062 17876
rect 14829 17867 14887 17873
rect 14829 17864 14841 17867
rect 14056 17836 14841 17864
rect 14056 17824 14062 17836
rect 14829 17833 14841 17836
rect 14875 17833 14887 17867
rect 14829 17827 14887 17833
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 16025 17867 16083 17873
rect 16025 17864 16037 17867
rect 15252 17836 16037 17864
rect 15252 17824 15258 17836
rect 16025 17833 16037 17836
rect 16071 17833 16083 17867
rect 16025 17827 16083 17833
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 21358 17864 21364 17876
rect 20128 17836 20392 17864
rect 21319 17836 21364 17864
rect 20128 17824 20134 17836
rect 1857 17799 1915 17805
rect 1857 17765 1869 17799
rect 1903 17796 1915 17799
rect 2314 17796 2320 17808
rect 1903 17768 2320 17796
rect 1903 17765 1915 17768
rect 1857 17759 1915 17765
rect 2314 17756 2320 17768
rect 2372 17756 2378 17808
rect 10594 17796 10600 17808
rect 10555 17768 10600 17796
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 15654 17796 15660 17808
rect 14752 17768 15660 17796
rect 12066 17728 12072 17740
rect 12027 17700 12072 17728
rect 12066 17688 12072 17700
rect 12124 17728 12130 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 12124 17700 13829 17728
rect 12124 17688 12130 17700
rect 13817 17697 13829 17700
rect 13863 17728 13875 17731
rect 13998 17728 14004 17740
rect 13863 17700 14004 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 14752 17737 14780 17768
rect 15654 17756 15660 17768
rect 15712 17756 15718 17808
rect 20162 17756 20168 17808
rect 20220 17805 20226 17808
rect 20220 17799 20284 17805
rect 20220 17765 20238 17799
rect 20272 17765 20284 17799
rect 20364 17796 20392 17836
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 21910 17864 21916 17876
rect 21871 17836 21916 17864
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 24121 17867 24179 17873
rect 24121 17864 24133 17867
rect 23532 17836 24133 17864
rect 23532 17824 23538 17836
rect 24121 17833 24133 17836
rect 24167 17833 24179 17867
rect 25314 17864 25320 17876
rect 25275 17836 25320 17864
rect 24121 17827 24179 17833
rect 25314 17824 25320 17836
rect 25372 17824 25378 17876
rect 26602 17824 26608 17876
rect 26660 17864 26666 17876
rect 27249 17867 27307 17873
rect 27249 17864 27261 17867
rect 26660 17836 27261 17864
rect 26660 17824 26666 17836
rect 27249 17833 27261 17836
rect 27295 17833 27307 17867
rect 27249 17827 27307 17833
rect 20364 17768 23336 17796
rect 20220 17759 20284 17765
rect 20220 17756 20226 17759
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17697 14795 17731
rect 14918 17728 14924 17740
rect 14879 17700 14924 17728
rect 14737 17691 14795 17697
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 16209 17731 16267 17737
rect 16209 17728 16221 17731
rect 15611 17700 16221 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 16209 17697 16221 17700
rect 16255 17728 16267 17731
rect 16298 17728 16304 17740
rect 16255 17700 16304 17728
rect 16255 17697 16267 17700
rect 16209 17691 16267 17697
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 19978 17728 19984 17740
rect 19939 17700 19984 17728
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 21818 17728 21824 17740
rect 21779 17700 21824 17728
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 22830 17728 22836 17740
rect 22791 17700 22836 17728
rect 22830 17688 22836 17700
rect 22888 17688 22894 17740
rect 23308 17737 23336 17768
rect 23382 17756 23388 17808
rect 23440 17796 23446 17808
rect 23440 17768 25360 17796
rect 23440 17756 23446 17768
rect 23293 17731 23351 17737
rect 23293 17697 23305 17731
rect 23339 17697 23351 17731
rect 24026 17728 24032 17740
rect 23987 17700 24032 17728
rect 23293 17691 23351 17697
rect 24026 17688 24032 17700
rect 24084 17688 24090 17740
rect 25130 17688 25136 17740
rect 25188 17728 25194 17740
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 25188 17700 25237 17728
rect 25188 17688 25194 17700
rect 25225 17697 25237 17700
rect 25271 17697 25283 17731
rect 25332 17728 25360 17768
rect 25498 17756 25504 17808
rect 25556 17796 25562 17808
rect 26114 17799 26172 17805
rect 26114 17796 26126 17799
rect 25556 17768 26126 17796
rect 25556 17756 25562 17768
rect 26114 17765 26126 17768
rect 26160 17765 26172 17799
rect 56597 17799 56655 17805
rect 56597 17796 56609 17799
rect 26114 17759 26172 17765
rect 31726 17768 56609 17796
rect 31726 17728 31754 17768
rect 56597 17765 56609 17768
rect 56643 17796 56655 17799
rect 58158 17796 58164 17808
rect 56643 17768 56732 17796
rect 58119 17768 58164 17796
rect 56643 17765 56655 17768
rect 56597 17759 56655 17765
rect 56704 17737 56732 17768
rect 58158 17756 58164 17768
rect 58216 17756 58222 17808
rect 25332 17700 31754 17728
rect 56689 17731 56747 17737
rect 25225 17691 25283 17697
rect 56689 17697 56701 17731
rect 56735 17697 56747 17731
rect 56689 17691 56747 17697
rect 57333 17731 57391 17737
rect 57333 17697 57345 17731
rect 57379 17728 57391 17731
rect 57977 17731 58035 17737
rect 57977 17728 57989 17731
rect 57379 17700 57989 17728
rect 57379 17697 57391 17700
rect 57333 17691 57391 17697
rect 57977 17697 57989 17700
rect 58023 17697 58035 17731
rect 57977 17691 58035 17697
rect 10502 17660 10508 17672
rect 10463 17632 10508 17660
rect 10502 17620 10508 17632
rect 10560 17620 10566 17672
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17629 10839 17663
rect 10781 17623 10839 17629
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 25774 17660 25780 17672
rect 23615 17632 25780 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 1762 17552 1768 17604
rect 1820 17592 1826 17604
rect 10796 17592 10824 17623
rect 25774 17620 25780 17632
rect 25832 17620 25838 17672
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17629 25927 17663
rect 25869 17623 25927 17629
rect 1820 17564 10824 17592
rect 1820 17552 1826 17564
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 15381 17595 15439 17601
rect 15381 17592 15393 17595
rect 12216 17564 15393 17592
rect 12216 17552 12222 17564
rect 15381 17561 15393 17564
rect 15427 17561 15439 17595
rect 15381 17555 15439 17561
rect 12250 17524 12256 17536
rect 12211 17496 12256 17524
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 13633 17527 13691 17533
rect 13633 17493 13645 17527
rect 13679 17524 13691 17527
rect 13814 17524 13820 17536
rect 13679 17496 13820 17524
rect 13679 17493 13691 17496
rect 13633 17487 13691 17493
rect 13814 17484 13820 17496
rect 13872 17484 13878 17536
rect 25884 17524 25912 17623
rect 55398 17620 55404 17672
rect 55456 17660 55462 17672
rect 56873 17663 56931 17669
rect 56873 17660 56885 17663
rect 55456 17632 56885 17660
rect 55456 17620 55462 17632
rect 56873 17629 56885 17632
rect 56919 17629 56931 17663
rect 56873 17623 56931 17629
rect 26142 17524 26148 17536
rect 25884 17496 26148 17524
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 1104 17434 58880 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 58880 17434
rect 1104 17360 58880 17382
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 15013 17323 15071 17329
rect 15013 17320 15025 17323
rect 14056 17292 15025 17320
rect 14056 17280 14062 17292
rect 15013 17289 15025 17292
rect 15059 17289 15071 17323
rect 15013 17283 15071 17289
rect 21361 17323 21419 17329
rect 21361 17289 21373 17323
rect 21407 17320 21419 17323
rect 21634 17320 21640 17332
rect 21407 17292 21640 17320
rect 21407 17289 21419 17292
rect 21361 17283 21419 17289
rect 21634 17280 21640 17292
rect 21692 17280 21698 17332
rect 24762 17320 24768 17332
rect 24723 17292 24768 17320
rect 24762 17280 24768 17292
rect 24820 17280 24826 17332
rect 25774 17280 25780 17332
rect 25832 17320 25838 17332
rect 55214 17320 55220 17332
rect 25832 17292 55220 17320
rect 25832 17280 25838 17292
rect 55214 17280 55220 17292
rect 55272 17280 55278 17332
rect 55398 17320 55404 17332
rect 55359 17292 55404 17320
rect 55398 17280 55404 17292
rect 55456 17280 55462 17332
rect 56318 17252 56324 17264
rect 56279 17224 56324 17252
rect 56318 17212 56324 17224
rect 56376 17212 56382 17264
rect 56873 17255 56931 17261
rect 56873 17221 56885 17255
rect 56919 17221 56931 17255
rect 56873 17215 56931 17221
rect 10318 17184 10324 17196
rect 10279 17156 10324 17184
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10410 17144 10416 17196
rect 10468 17184 10474 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10468 17156 10609 17184
rect 10468 17144 10474 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17184 12219 17187
rect 12986 17184 12992 17196
rect 12207 17156 12992 17184
rect 12207 17153 12219 17156
rect 12161 17147 12219 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 14182 17184 14188 17196
rect 13771 17156 14188 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 20346 17144 20352 17196
rect 20404 17184 20410 17196
rect 23382 17184 23388 17196
rect 20404 17156 23244 17184
rect 23343 17156 23388 17184
rect 20404 17144 20410 17156
rect 1857 17119 1915 17125
rect 1857 17085 1869 17119
rect 1903 17116 1915 17119
rect 5534 17116 5540 17128
rect 1903 17088 5540 17116
rect 1903 17085 1915 17088
rect 1857 17079 1915 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 9766 17116 9772 17128
rect 9727 17088 9772 17116
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17085 14887 17119
rect 14829 17079 14887 17085
rect 21269 17119 21327 17125
rect 21269 17085 21281 17119
rect 21315 17116 21327 17119
rect 21358 17116 21364 17128
rect 21315 17088 21364 17116
rect 21315 17085 21327 17088
rect 21269 17079 21327 17085
rect 2038 17048 2044 17060
rect 1999 17020 2044 17048
rect 2038 17008 2044 17020
rect 2096 17008 2102 17060
rect 10413 17051 10471 17057
rect 10413 17048 10425 17051
rect 9600 17020 10425 17048
rect 9600 16989 9628 17020
rect 10413 17017 10425 17020
rect 10459 17017 10471 17051
rect 10413 17011 10471 17017
rect 12250 17008 12256 17060
rect 12308 17048 12314 17060
rect 13170 17048 13176 17060
rect 12308 17020 12353 17048
rect 13131 17020 13176 17048
rect 12308 17008 12314 17020
rect 13170 17008 13176 17020
rect 13228 17008 13234 17060
rect 13814 17008 13820 17060
rect 13872 17048 13878 17060
rect 14369 17051 14427 17057
rect 13872 17020 13917 17048
rect 13872 17008 13878 17020
rect 14369 17017 14381 17051
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 9585 16983 9643 16989
rect 9585 16949 9597 16983
rect 9631 16949 9643 16983
rect 9585 16943 9643 16949
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 14384 16980 14412 17011
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 14844 17048 14872 17079
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 22830 17116 22836 17128
rect 22791 17088 22836 17116
rect 22830 17076 22836 17088
rect 22888 17076 22894 17128
rect 23216 17125 23244 17156
rect 23382 17144 23388 17156
rect 23440 17144 23446 17196
rect 56888 17184 56916 17215
rect 57701 17187 57759 17193
rect 57701 17184 57713 17187
rect 56888 17156 57713 17184
rect 57701 17153 57713 17156
rect 57747 17153 57759 17187
rect 57701 17147 57759 17153
rect 23201 17119 23259 17125
rect 23201 17085 23213 17119
rect 23247 17085 23259 17119
rect 24118 17116 24124 17128
rect 24079 17088 24124 17116
rect 23201 17079 23259 17085
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 55585 17119 55643 17125
rect 55585 17085 55597 17119
rect 55631 17116 55643 17119
rect 55766 17116 55772 17128
rect 55631 17088 55772 17116
rect 55631 17085 55643 17088
rect 55585 17079 55643 17085
rect 55766 17076 55772 17088
rect 55824 17076 55830 17128
rect 57054 17116 57060 17128
rect 57015 17088 57060 17116
rect 57054 17076 57060 17088
rect 57112 17076 57118 17128
rect 57514 17116 57520 17128
rect 57475 17088 57520 17116
rect 57514 17076 57520 17088
rect 57572 17076 57578 17128
rect 53742 17048 53748 17060
rect 14792 17020 53748 17048
rect 14792 17008 14798 17020
rect 53742 17008 53748 17020
rect 53800 17048 53806 17060
rect 56137 17051 56195 17057
rect 56137 17048 56149 17051
rect 53800 17020 56149 17048
rect 53800 17008 53806 17020
rect 56137 17017 56149 17020
rect 56183 17017 56195 17051
rect 56137 17011 56195 17017
rect 9732 16952 14412 16980
rect 9732 16940 9738 16952
rect 57974 16940 57980 16992
rect 58032 16980 58038 16992
rect 58161 16983 58219 16989
rect 58161 16980 58173 16983
rect 58032 16952 58173 16980
rect 58032 16940 58038 16952
rect 58161 16949 58173 16952
rect 58207 16949 58219 16983
rect 58161 16943 58219 16949
rect 1104 16890 58880 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 50326 16890
rect 50378 16838 50390 16890
rect 50442 16838 50454 16890
rect 50506 16838 50518 16890
rect 50570 16838 58880 16890
rect 1104 16816 58880 16838
rect 1854 16736 1860 16788
rect 1912 16776 1918 16788
rect 9674 16776 9680 16788
rect 1912 16748 9680 16776
rect 1912 16736 1918 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10594 16776 10600 16788
rect 10555 16748 10600 16776
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 13906 16776 13912 16788
rect 13863 16748 13912 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 24118 16776 24124 16788
rect 24079 16748 24124 16776
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 55585 16779 55643 16785
rect 31726 16748 45554 16776
rect 2130 16668 2136 16720
rect 2188 16708 2194 16720
rect 10410 16708 10416 16720
rect 2188 16680 10416 16708
rect 2188 16668 2194 16680
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 21542 16668 21548 16720
rect 21600 16708 21606 16720
rect 23569 16711 23627 16717
rect 21600 16680 23336 16708
rect 21600 16668 21606 16680
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 9824 16612 10793 16640
rect 9824 16600 9830 16612
rect 10781 16609 10793 16612
rect 10827 16640 10839 16643
rect 12066 16640 12072 16652
rect 10827 16612 12072 16640
rect 10827 16609 10839 16612
rect 10781 16603 10839 16609
rect 12066 16600 12072 16612
rect 12124 16640 12130 16652
rect 13633 16643 13691 16649
rect 13633 16640 13645 16643
rect 12124 16612 13645 16640
rect 12124 16600 12130 16612
rect 13633 16609 13645 16612
rect 13679 16609 13691 16643
rect 22830 16640 22836 16652
rect 22791 16612 22836 16640
rect 13633 16603 13691 16609
rect 22830 16600 22836 16612
rect 22888 16600 22894 16652
rect 23308 16649 23336 16680
rect 23569 16677 23581 16711
rect 23615 16708 23627 16711
rect 31726 16708 31754 16748
rect 23615 16680 31754 16708
rect 23615 16677 23627 16680
rect 23569 16671 23627 16677
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16609 23351 16643
rect 23293 16603 23351 16609
rect 24029 16643 24087 16649
rect 24029 16609 24041 16643
rect 24075 16609 24087 16643
rect 24210 16640 24216 16652
rect 24171 16612 24216 16640
rect 24029 16603 24087 16609
rect 24044 16572 24072 16603
rect 24210 16600 24216 16612
rect 24268 16600 24274 16652
rect 26050 16640 26056 16652
rect 24320 16612 26056 16640
rect 24320 16572 24348 16612
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 45526 16640 45554 16748
rect 55585 16745 55597 16779
rect 55631 16776 55643 16779
rect 55631 16748 57008 16776
rect 55631 16745 55643 16748
rect 55585 16739 55643 16745
rect 55766 16640 55772 16652
rect 45526 16612 55628 16640
rect 55727 16612 55772 16640
rect 24044 16544 24348 16572
rect 55600 16572 55628 16612
rect 55766 16600 55772 16612
rect 55824 16600 55830 16652
rect 56980 16649 57008 16748
rect 57974 16708 57980 16720
rect 57935 16680 57980 16708
rect 57974 16668 57980 16680
rect 58032 16668 58038 16720
rect 58158 16708 58164 16720
rect 58119 16680 58164 16708
rect 58158 16668 58164 16680
rect 58216 16668 58222 16720
rect 56781 16643 56839 16649
rect 56781 16640 56793 16643
rect 55876 16612 56793 16640
rect 55876 16572 55904 16612
rect 56781 16609 56793 16612
rect 56827 16609 56839 16643
rect 56781 16603 56839 16609
rect 56965 16643 57023 16649
rect 56965 16609 56977 16643
rect 57011 16609 57023 16643
rect 56965 16603 57023 16609
rect 57425 16643 57483 16649
rect 57425 16609 57437 16643
rect 57471 16640 57483 16643
rect 57471 16612 58020 16640
rect 57471 16609 57483 16612
rect 57425 16603 57483 16609
rect 57992 16584 58020 16612
rect 55600 16544 55904 16572
rect 57974 16532 57980 16584
rect 58032 16532 58038 16584
rect 1104 16346 58880 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 58880 16346
rect 1104 16272 58880 16294
rect 56594 16192 56600 16244
rect 56652 16232 56658 16244
rect 56965 16235 57023 16241
rect 56965 16232 56977 16235
rect 56652 16204 56977 16232
rect 56652 16192 56658 16204
rect 56965 16201 56977 16204
rect 57011 16201 57023 16235
rect 56965 16195 57023 16201
rect 55677 16167 55735 16173
rect 55677 16133 55689 16167
rect 55723 16164 55735 16167
rect 57514 16164 57520 16176
rect 55723 16136 57520 16164
rect 55723 16133 55735 16136
rect 55677 16127 55735 16133
rect 57514 16124 57520 16136
rect 57572 16124 57578 16176
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 4706 16056 4712 16108
rect 4764 16096 4770 16108
rect 4982 16096 4988 16108
rect 4764 16068 4988 16096
rect 4764 16056 4770 16068
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 16028 1915 16031
rect 5810 16028 5816 16040
rect 1903 16000 5816 16028
rect 1903 15997 1915 16000
rect 1857 15991 1915 15997
rect 5810 15988 5816 16000
rect 5868 15988 5874 16040
rect 14734 16028 14740 16040
rect 14695 16000 14740 16028
rect 14734 15988 14740 16000
rect 14792 15988 14798 16040
rect 54849 16031 54907 16037
rect 54849 15997 54861 16031
rect 54895 16028 54907 16031
rect 55582 16028 55588 16040
rect 54895 16000 55588 16028
rect 54895 15997 54907 16000
rect 54849 15991 54907 15997
rect 55582 15988 55588 16000
rect 55640 15988 55646 16040
rect 56137 16031 56195 16037
rect 56137 15997 56149 16031
rect 56183 16028 56195 16031
rect 56318 16028 56324 16040
rect 56183 16000 56324 16028
rect 56183 15997 56195 16000
rect 56137 15991 56195 15997
rect 56318 15988 56324 16000
rect 56376 15988 56382 16040
rect 15010 15960 15016 15972
rect 14971 15932 15016 15960
rect 15010 15920 15016 15932
rect 15068 15920 15074 15972
rect 56873 15963 56931 15969
rect 56873 15929 56885 15963
rect 56919 15960 56931 15963
rect 57054 15960 57060 15972
rect 56919 15932 57060 15960
rect 56919 15929 56931 15932
rect 56873 15923 56931 15929
rect 57054 15920 57060 15932
rect 57112 15920 57118 15972
rect 57977 15963 58035 15969
rect 57977 15929 57989 15963
rect 58023 15960 58035 15963
rect 58158 15960 58164 15972
rect 58023 15932 58164 15960
rect 58023 15929 58035 15932
rect 57977 15923 58035 15929
rect 58158 15920 58164 15932
rect 58216 15920 58222 15972
rect 56318 15892 56324 15904
rect 56279 15864 56324 15892
rect 56318 15852 56324 15864
rect 56376 15852 56382 15904
rect 58066 15892 58072 15904
rect 58027 15864 58072 15892
rect 58066 15852 58072 15864
rect 58124 15852 58130 15904
rect 1104 15802 58880 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 50326 15802
rect 50378 15750 50390 15802
rect 50442 15750 50454 15802
rect 50506 15750 50518 15802
rect 50570 15750 58880 15802
rect 1104 15728 58880 15750
rect 58158 15688 58164 15700
rect 58119 15660 58164 15688
rect 58158 15648 58164 15660
rect 58216 15648 58222 15700
rect 55769 15555 55827 15561
rect 55769 15521 55781 15555
rect 55815 15552 55827 15555
rect 56318 15552 56324 15564
rect 55815 15524 56324 15552
rect 55815 15521 55827 15524
rect 55769 15515 55827 15521
rect 56318 15512 56324 15524
rect 56376 15552 56382 15564
rect 56686 15552 56692 15564
rect 56376 15524 56692 15552
rect 56376 15512 56382 15524
rect 56686 15512 56692 15524
rect 56744 15512 56750 15564
rect 56870 15552 56876 15564
rect 56831 15524 56876 15552
rect 56870 15512 56876 15524
rect 56928 15512 56934 15564
rect 55125 15487 55183 15493
rect 55125 15453 55137 15487
rect 55171 15484 55183 15487
rect 57517 15487 57575 15493
rect 57517 15484 57529 15487
rect 55171 15456 57529 15484
rect 55171 15453 55183 15456
rect 55125 15447 55183 15453
rect 57517 15453 57529 15456
rect 57563 15453 57575 15487
rect 57517 15447 57575 15453
rect 57701 15487 57759 15493
rect 57701 15453 57713 15487
rect 57747 15453 57759 15487
rect 57701 15447 57759 15453
rect 55585 15419 55643 15425
rect 55585 15385 55597 15419
rect 55631 15416 55643 15419
rect 57716 15416 57744 15447
rect 55631 15388 57744 15416
rect 55631 15385 55643 15388
rect 55585 15379 55643 15385
rect 56962 15348 56968 15360
rect 56923 15320 56968 15348
rect 56962 15308 56968 15320
rect 57020 15308 57026 15360
rect 1104 15258 58880 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 58880 15258
rect 1104 15184 58880 15206
rect 1946 15144 1952 15156
rect 1907 15116 1952 15144
rect 1946 15104 1952 15116
rect 2004 15104 2010 15156
rect 55214 15104 55220 15156
rect 55272 15144 55278 15156
rect 56321 15147 56379 15153
rect 56321 15144 56333 15147
rect 55272 15116 56333 15144
rect 55272 15104 55278 15116
rect 56321 15113 56333 15116
rect 56367 15144 56379 15147
rect 56413 15147 56471 15153
rect 56413 15144 56425 15147
rect 56367 15116 56425 15144
rect 56367 15113 56379 15116
rect 56321 15107 56379 15113
rect 56413 15113 56425 15116
rect 56459 15113 56471 15147
rect 56413 15107 56471 15113
rect 56870 15104 56876 15156
rect 56928 15144 56934 15156
rect 56965 15147 57023 15153
rect 56965 15144 56977 15147
rect 56928 15116 56977 15144
rect 56928 15104 56934 15116
rect 56965 15113 56977 15116
rect 57011 15113 57023 15147
rect 56965 15107 57023 15113
rect 55953 15079 56011 15085
rect 55953 15045 55965 15079
rect 55999 15045 56011 15079
rect 55953 15039 56011 15045
rect 58161 15079 58219 15085
rect 58161 15045 58173 15079
rect 58207 15076 58219 15079
rect 58250 15076 58256 15088
rect 58207 15048 58256 15076
rect 58207 15045 58219 15048
rect 58161 15039 58219 15045
rect 55968 15008 55996 15039
rect 58250 15036 58256 15048
rect 58308 15036 58314 15088
rect 56781 15011 56839 15017
rect 56781 15008 56793 15011
rect 55968 14980 56793 15008
rect 56781 14977 56793 14980
rect 56827 14977 56839 15011
rect 56781 14971 56839 14977
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 7374 14940 7380 14952
rect 1903 14912 7380 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 55766 14900 55772 14952
rect 55824 14940 55830 14952
rect 56134 14940 56140 14952
rect 55824 14912 56140 14940
rect 55824 14900 55830 14912
rect 56134 14900 56140 14912
rect 56192 14900 56198 14952
rect 56321 14943 56379 14949
rect 56321 14909 56333 14943
rect 56367 14940 56379 14943
rect 56597 14943 56655 14949
rect 56597 14940 56609 14943
rect 56367 14912 56609 14940
rect 56367 14909 56379 14912
rect 56321 14903 56379 14909
rect 56597 14909 56609 14912
rect 56643 14909 56655 14943
rect 57974 14940 57980 14952
rect 57935 14912 57980 14940
rect 56597 14903 56655 14909
rect 57974 14900 57980 14912
rect 58032 14900 58038 14952
rect 1104 14714 58880 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 50326 14714
rect 50378 14662 50390 14714
rect 50442 14662 50454 14714
rect 50506 14662 50518 14714
rect 50570 14662 58880 14714
rect 1104 14640 58880 14662
rect 56781 14603 56839 14609
rect 56781 14569 56793 14603
rect 56827 14600 56839 14603
rect 56827 14572 57652 14600
rect 56827 14569 56839 14572
rect 56781 14563 56839 14569
rect 1857 14535 1915 14541
rect 1857 14501 1869 14535
rect 1903 14532 1915 14535
rect 7558 14532 7564 14544
rect 1903 14504 7564 14532
rect 1903 14501 1915 14504
rect 1857 14495 1915 14501
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 57624 14541 57652 14572
rect 57609 14535 57667 14541
rect 57609 14501 57621 14535
rect 57655 14501 57667 14535
rect 57609 14495 57667 14501
rect 55582 14464 55588 14476
rect 55543 14436 55588 14464
rect 55582 14424 55588 14436
rect 55640 14424 55646 14476
rect 56594 14424 56600 14476
rect 56652 14464 56658 14476
rect 56965 14467 57023 14473
rect 56965 14464 56977 14467
rect 56652 14436 56977 14464
rect 56652 14424 56658 14436
rect 56965 14433 56977 14436
rect 57011 14433 57023 14467
rect 56965 14427 57023 14433
rect 55766 14356 55772 14408
rect 55824 14396 55830 14408
rect 57517 14399 57575 14405
rect 57517 14396 57529 14399
rect 55824 14368 57529 14396
rect 55824 14356 55830 14368
rect 57517 14365 57529 14368
rect 57563 14365 57575 14399
rect 57517 14359 57575 14365
rect 57793 14399 57851 14405
rect 57793 14365 57805 14399
rect 57839 14365 57851 14399
rect 57793 14359 57851 14365
rect 53834 14288 53840 14340
rect 53892 14328 53898 14340
rect 57808 14328 57836 14359
rect 53892 14300 57836 14328
rect 53892 14288 53898 14300
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 1104 14170 58880 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 58880 14170
rect 1104 14096 58880 14118
rect 55766 14056 55772 14068
rect 55727 14028 55772 14056
rect 55766 14016 55772 14028
rect 55824 14016 55830 14068
rect 56229 13991 56287 13997
rect 56229 13957 56241 13991
rect 56275 13988 56287 13991
rect 56778 13988 56784 14000
rect 56275 13960 56784 13988
rect 56275 13957 56287 13960
rect 56229 13951 56287 13957
rect 56778 13948 56784 13960
rect 56836 13948 56842 14000
rect 56873 13991 56931 13997
rect 56873 13957 56885 13991
rect 56919 13957 56931 13991
rect 56873 13951 56931 13957
rect 56888 13920 56916 13951
rect 57701 13923 57759 13929
rect 57701 13920 57713 13923
rect 56888 13892 57713 13920
rect 57701 13889 57713 13892
rect 57747 13889 57759 13923
rect 57701 13883 57759 13889
rect 56134 13812 56140 13864
rect 56192 13852 56198 13864
rect 56413 13855 56471 13861
rect 56413 13852 56425 13855
rect 56192 13824 56425 13852
rect 56192 13812 56198 13824
rect 56413 13821 56425 13824
rect 56459 13821 56471 13855
rect 56413 13815 56471 13821
rect 56686 13812 56692 13864
rect 56744 13852 56750 13864
rect 57057 13855 57115 13861
rect 57057 13852 57069 13855
rect 56744 13824 57069 13852
rect 56744 13812 56750 13824
rect 57057 13821 57069 13824
rect 57103 13852 57115 13855
rect 57146 13852 57152 13864
rect 57103 13824 57152 13852
rect 57103 13821 57115 13824
rect 57057 13815 57115 13821
rect 57146 13812 57152 13824
rect 57204 13812 57210 13864
rect 57514 13852 57520 13864
rect 57475 13824 57520 13852
rect 57514 13812 57520 13824
rect 57572 13812 57578 13864
rect 58158 13716 58164 13728
rect 58119 13688 58164 13716
rect 58158 13676 58164 13688
rect 58216 13676 58222 13728
rect 1104 13626 58880 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 50326 13626
rect 50378 13574 50390 13626
rect 50442 13574 50454 13626
rect 50506 13574 50518 13626
rect 50570 13574 58880 13626
rect 1104 13552 58880 13574
rect 58066 13512 58072 13524
rect 58027 13484 58072 13512
rect 58066 13472 58072 13484
rect 58124 13472 58130 13524
rect 1857 13447 1915 13453
rect 1857 13413 1869 13447
rect 1903 13444 1915 13447
rect 7466 13444 7472 13456
rect 1903 13416 7472 13444
rect 1903 13413 1915 13416
rect 1857 13407 1915 13413
rect 7466 13404 7472 13416
rect 7524 13404 7530 13456
rect 57514 13444 57520 13456
rect 55784 13416 57520 13444
rect 55784 13385 55812 13416
rect 57514 13404 57520 13416
rect 57572 13404 57578 13456
rect 57977 13447 58035 13453
rect 57977 13413 57989 13447
rect 58023 13444 58035 13447
rect 58158 13444 58164 13456
rect 58023 13416 58164 13444
rect 58023 13413 58035 13416
rect 57977 13407 58035 13413
rect 58158 13404 58164 13416
rect 58216 13404 58222 13456
rect 55769 13379 55827 13385
rect 55769 13345 55781 13379
rect 55815 13345 55827 13379
rect 55769 13339 55827 13345
rect 56778 13336 56784 13388
rect 56836 13376 56842 13388
rect 56873 13379 56931 13385
rect 56873 13376 56885 13379
rect 56836 13348 56885 13376
rect 56836 13336 56842 13348
rect 56873 13345 56885 13348
rect 56919 13345 56931 13379
rect 56873 13339 56931 13345
rect 56689 13311 56747 13317
rect 56689 13277 56701 13311
rect 56735 13277 56747 13311
rect 56689 13271 56747 13277
rect 2038 13240 2044 13252
rect 1999 13212 2044 13240
rect 2038 13200 2044 13212
rect 2096 13200 2102 13252
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 56597 13243 56655 13249
rect 56597 13240 56609 13243
rect 23440 13212 56609 13240
rect 23440 13200 23446 13212
rect 56597 13209 56609 13212
rect 56643 13240 56655 13243
rect 56704 13240 56732 13271
rect 56643 13212 56732 13240
rect 56643 13209 56655 13212
rect 56597 13203 56655 13209
rect 57238 13172 57244 13184
rect 57199 13144 57244 13172
rect 57238 13132 57244 13144
rect 57296 13132 57302 13184
rect 1104 13082 58880 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 58880 13082
rect 1104 13008 58880 13030
rect 56134 12928 56140 12980
rect 56192 12968 56198 12980
rect 56229 12971 56287 12977
rect 56229 12968 56241 12971
rect 56192 12940 56241 12968
rect 56192 12928 56198 12940
rect 56229 12937 56241 12940
rect 56275 12937 56287 12971
rect 57330 12968 57336 12980
rect 57291 12940 57336 12968
rect 56229 12931 56287 12937
rect 57330 12928 57336 12940
rect 57388 12928 57394 12980
rect 55398 12764 55404 12776
rect 55359 12736 55404 12764
rect 55398 12724 55404 12736
rect 55456 12724 55462 12776
rect 56042 12764 56048 12776
rect 56003 12736 56048 12764
rect 56042 12724 56048 12736
rect 56100 12724 56106 12776
rect 57238 12764 57244 12776
rect 57199 12736 57244 12764
rect 57238 12724 57244 12736
rect 57296 12724 57302 12776
rect 57974 12696 57980 12708
rect 57935 12668 57980 12696
rect 57974 12656 57980 12668
rect 58032 12656 58038 12708
rect 57882 12588 57888 12640
rect 57940 12628 57946 12640
rect 58069 12631 58127 12637
rect 58069 12628 58081 12631
rect 57940 12600 58081 12628
rect 57940 12588 57946 12600
rect 58069 12597 58081 12600
rect 58115 12597 58127 12631
rect 58069 12591 58127 12597
rect 1104 12538 58880 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 50326 12538
rect 50378 12486 50390 12538
rect 50442 12486 50454 12538
rect 50506 12486 50518 12538
rect 50570 12486 58880 12538
rect 1104 12464 58880 12486
rect 1946 12424 1952 12436
rect 1907 12396 1952 12424
rect 1946 12384 1952 12396
rect 2004 12384 2010 12436
rect 57974 12384 57980 12436
rect 58032 12424 58038 12436
rect 58161 12427 58219 12433
rect 58161 12424 58173 12427
rect 58032 12396 58173 12424
rect 58032 12384 58038 12396
rect 58161 12393 58173 12396
rect 58207 12393 58219 12427
rect 58161 12387 58219 12393
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 4890 12356 4896 12368
rect 1903 12328 4896 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 4890 12316 4896 12328
rect 4948 12316 4954 12368
rect 56870 12288 56876 12300
rect 56831 12260 56876 12288
rect 56870 12248 56876 12260
rect 56928 12248 56934 12300
rect 55582 12180 55588 12232
rect 55640 12220 55646 12232
rect 57517 12223 57575 12229
rect 57517 12220 57529 12223
rect 55640 12192 57529 12220
rect 55640 12180 55646 12192
rect 57517 12189 57529 12192
rect 57563 12189 57575 12223
rect 57698 12220 57704 12232
rect 57659 12192 57704 12220
rect 57517 12183 57575 12189
rect 57698 12180 57704 12192
rect 57756 12180 57762 12232
rect 56502 12044 56508 12096
rect 56560 12084 56566 12096
rect 56965 12087 57023 12093
rect 56965 12084 56977 12087
rect 56560 12056 56977 12084
rect 56560 12044 56566 12056
rect 56965 12053 56977 12056
rect 57011 12053 57023 12087
rect 56965 12047 57023 12053
rect 1104 11994 58880 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 58880 11994
rect 1104 11920 58880 11942
rect 55582 11880 55588 11892
rect 55543 11852 55588 11880
rect 55582 11840 55588 11852
rect 55640 11840 55646 11892
rect 56870 11840 56876 11892
rect 56928 11880 56934 11892
rect 57701 11883 57759 11889
rect 57701 11880 57713 11883
rect 56928 11852 57713 11880
rect 56928 11840 56934 11852
rect 57701 11849 57713 11852
rect 57747 11849 57759 11883
rect 57701 11843 57759 11849
rect 56689 11815 56747 11821
rect 56689 11781 56701 11815
rect 56735 11812 56747 11815
rect 56735 11784 57560 11812
rect 56735 11781 56747 11784
rect 56689 11775 56747 11781
rect 57532 11753 57560 11784
rect 56229 11747 56287 11753
rect 56229 11713 56241 11747
rect 56275 11744 56287 11747
rect 57333 11747 57391 11753
rect 57333 11744 57345 11747
rect 56275 11716 57345 11744
rect 56275 11713 56287 11716
rect 56229 11707 56287 11713
rect 57333 11713 57345 11716
rect 57379 11713 57391 11747
rect 57333 11707 57391 11713
rect 57517 11747 57575 11753
rect 57517 11713 57529 11747
rect 57563 11713 57575 11747
rect 57517 11707 57575 11713
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 4798 11676 4804 11688
rect 1903 11648 4804 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 56134 11636 56140 11688
rect 56192 11676 56198 11688
rect 56873 11679 56931 11685
rect 56873 11676 56885 11679
rect 56192 11648 56885 11676
rect 56192 11636 56198 11648
rect 56873 11645 56885 11648
rect 56919 11645 56931 11679
rect 56873 11639 56931 11645
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 1104 11450 58880 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 50326 11450
rect 50378 11398 50390 11450
rect 50442 11398 50454 11450
rect 50506 11398 50518 11450
rect 50570 11398 58880 11450
rect 1104 11376 58880 11398
rect 57241 11339 57299 11345
rect 57241 11305 57253 11339
rect 57287 11336 57299 11339
rect 57698 11336 57704 11348
rect 57287 11308 57704 11336
rect 57287 11305 57299 11308
rect 57241 11299 57299 11305
rect 57698 11296 57704 11308
rect 57756 11296 57762 11348
rect 55582 11200 55588 11212
rect 55543 11172 55588 11200
rect 55582 11160 55588 11172
rect 55640 11160 55646 11212
rect 57146 11160 57152 11212
rect 57204 11200 57210 11212
rect 57425 11203 57483 11209
rect 57425 11200 57437 11203
rect 57204 11172 57437 11200
rect 57204 11160 57210 11172
rect 57425 11169 57437 11172
rect 57471 11169 57483 11203
rect 57974 11200 57980 11212
rect 57935 11172 57980 11200
rect 57425 11163 57483 11169
rect 57974 11160 57980 11172
rect 58032 11160 58038 11212
rect 57882 11024 57888 11076
rect 57940 11064 57946 11076
rect 58161 11067 58219 11073
rect 58161 11064 58173 11067
rect 57940 11036 58173 11064
rect 57940 11024 57946 11036
rect 58161 11033 58173 11036
rect 58207 11033 58219 11067
rect 58161 11027 58219 11033
rect 1104 10906 58880 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 58880 10906
rect 1104 10832 58880 10854
rect 57974 10792 57980 10804
rect 57935 10764 57980 10792
rect 57974 10752 57980 10764
rect 58032 10752 58038 10804
rect 56413 10659 56471 10665
rect 56413 10625 56425 10659
rect 56459 10656 56471 10659
rect 57517 10659 57575 10665
rect 57517 10656 57529 10659
rect 56459 10628 57529 10656
rect 56459 10625 56471 10628
rect 56413 10619 56471 10625
rect 57517 10625 57529 10628
rect 57563 10625 57575 10659
rect 57517 10619 57575 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10588 1915 10591
rect 3602 10588 3608 10600
rect 1903 10560 3608 10588
rect 1903 10557 1915 10560
rect 1857 10551 1915 10557
rect 3602 10548 3608 10560
rect 3660 10548 3666 10600
rect 57057 10591 57115 10597
rect 57057 10557 57069 10591
rect 57103 10588 57115 10591
rect 57146 10588 57152 10600
rect 57103 10560 57152 10588
rect 57103 10557 57115 10560
rect 57057 10551 57115 10557
rect 57146 10548 57152 10560
rect 57204 10548 57210 10600
rect 57238 10548 57244 10600
rect 57296 10588 57302 10600
rect 57701 10591 57759 10597
rect 57701 10588 57713 10591
rect 57296 10560 57713 10588
rect 57296 10548 57302 10560
rect 57701 10557 57713 10560
rect 57747 10557 57759 10591
rect 57701 10551 57759 10557
rect 2038 10520 2044 10532
rect 1999 10492 2044 10520
rect 2038 10480 2044 10492
rect 2096 10480 2102 10532
rect 56873 10455 56931 10461
rect 56873 10421 56885 10455
rect 56919 10452 56931 10455
rect 57698 10452 57704 10464
rect 56919 10424 57704 10452
rect 56919 10421 56931 10424
rect 56873 10415 56931 10421
rect 57698 10412 57704 10424
rect 57756 10412 57762 10464
rect 1104 10362 58880 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 50326 10362
rect 50378 10310 50390 10362
rect 50442 10310 50454 10362
rect 50506 10310 50518 10362
rect 50570 10310 58880 10362
rect 1104 10288 58880 10310
rect 57238 10248 57244 10260
rect 57199 10220 57244 10248
rect 57238 10208 57244 10220
rect 57296 10208 57302 10260
rect 55582 10112 55588 10124
rect 55543 10084 55588 10112
rect 55582 10072 55588 10084
rect 55640 10072 55646 10124
rect 57146 10072 57152 10124
rect 57204 10112 57210 10124
rect 57425 10115 57483 10121
rect 57425 10112 57437 10115
rect 57204 10084 57437 10112
rect 57204 10072 57210 10084
rect 57425 10081 57437 10084
rect 57471 10081 57483 10115
rect 57425 10075 57483 10081
rect 57606 10072 57612 10124
rect 57664 10112 57670 10124
rect 57977 10115 58035 10121
rect 57977 10112 57989 10115
rect 57664 10084 57989 10112
rect 57664 10072 57670 10084
rect 57977 10081 57989 10084
rect 58023 10081 58035 10115
rect 57977 10075 58035 10081
rect 58158 9976 58164 9988
rect 58119 9948 58164 9976
rect 58158 9936 58164 9948
rect 58216 9936 58222 9988
rect 1104 9818 58880 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 58880 9818
rect 1104 9744 58880 9766
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 57606 9636 57612 9648
rect 57567 9608 57612 9636
rect 57606 9596 57612 9608
rect 57664 9596 57670 9648
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9500 1915 9503
rect 4062 9500 4068 9512
rect 1903 9472 4068 9500
rect 1903 9469 1915 9472
rect 1857 9463 1915 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 55674 9500 55680 9512
rect 55635 9472 55680 9500
rect 55674 9460 55680 9472
rect 55732 9460 55738 9512
rect 56505 9503 56563 9509
rect 56505 9469 56517 9503
rect 56551 9500 56563 9503
rect 56778 9500 56784 9512
rect 56551 9472 56784 9500
rect 56551 9469 56563 9472
rect 56505 9463 56563 9469
rect 56778 9460 56784 9472
rect 56836 9460 56842 9512
rect 56962 9500 56968 9512
rect 56923 9472 56968 9500
rect 56962 9460 56968 9472
rect 57020 9460 57026 9512
rect 57146 9500 57152 9512
rect 57107 9472 57152 9500
rect 57146 9460 57152 9472
rect 57204 9460 57210 9512
rect 1104 9274 58880 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 50326 9274
rect 50378 9222 50390 9274
rect 50442 9222 50454 9274
rect 50506 9222 50518 9274
rect 50570 9222 58880 9274
rect 1104 9200 58880 9222
rect 56873 9163 56931 9169
rect 56873 9129 56885 9163
rect 56919 9160 56931 9163
rect 57146 9160 57152 9172
rect 56919 9132 57152 9160
rect 56919 9129 56931 9132
rect 56873 9123 56931 9129
rect 57146 9120 57152 9132
rect 57204 9120 57210 9172
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 2958 9092 2964 9104
rect 1903 9064 2964 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 56134 9052 56140 9104
rect 56192 9092 56198 9104
rect 56192 9064 57100 9092
rect 56192 9052 56198 9064
rect 55769 9027 55827 9033
rect 55769 8993 55781 9027
rect 55815 9024 55827 9027
rect 56962 9024 56968 9036
rect 55815 8996 56968 9024
rect 55815 8993 55827 8996
rect 55769 8987 55827 8993
rect 56962 8984 56968 8996
rect 57020 8984 57026 9036
rect 57072 9033 57100 9064
rect 57057 9027 57115 9033
rect 57057 8993 57069 9027
rect 57103 8993 57115 9027
rect 57698 9024 57704 9036
rect 57659 8996 57704 9024
rect 57057 8987 57115 8993
rect 57698 8984 57704 8996
rect 57756 8984 57762 9036
rect 55125 8959 55183 8965
rect 55125 8925 55137 8959
rect 55171 8956 55183 8959
rect 57517 8959 57575 8965
rect 57517 8956 57529 8959
rect 55171 8928 57529 8956
rect 55171 8925 55183 8928
rect 55125 8919 55183 8925
rect 57517 8925 57529 8928
rect 57563 8925 57575 8959
rect 57517 8919 57575 8925
rect 1946 8820 1952 8832
rect 1907 8792 1952 8820
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 57974 8820 57980 8832
rect 57935 8792 57980 8820
rect 57974 8780 57980 8792
rect 58032 8780 58038 8832
rect 1104 8730 58880 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 58880 8730
rect 1104 8656 58880 8678
rect 56134 8616 56140 8628
rect 56095 8588 56140 8616
rect 56134 8576 56140 8588
rect 56192 8576 56198 8628
rect 55309 8551 55367 8557
rect 55309 8517 55321 8551
rect 55355 8548 55367 8551
rect 57330 8548 57336 8560
rect 55355 8520 57336 8548
rect 55355 8517 55367 8520
rect 55309 8511 55367 8517
rect 57330 8508 57336 8520
rect 57388 8508 57394 8560
rect 58158 8548 58164 8560
rect 58119 8520 58164 8548
rect 58158 8508 58164 8520
rect 58216 8508 58222 8560
rect 54849 8483 54907 8489
rect 54849 8449 54861 8483
rect 54895 8480 54907 8483
rect 56410 8480 56416 8492
rect 54895 8452 56416 8480
rect 54895 8449 54907 8452
rect 54849 8443 54907 8449
rect 56410 8440 56416 8452
rect 56468 8440 56474 8492
rect 57422 8480 57428 8492
rect 57383 8452 57428 8480
rect 57422 8440 57428 8452
rect 57480 8440 57486 8492
rect 55493 8415 55551 8421
rect 55493 8381 55505 8415
rect 55539 8381 55551 8415
rect 55493 8375 55551 8381
rect 55953 8415 56011 8421
rect 55953 8381 55965 8415
rect 55999 8412 56011 8415
rect 56042 8412 56048 8424
rect 55999 8384 56048 8412
rect 55999 8381 56011 8384
rect 55953 8375 56011 8381
rect 55508 8344 55536 8375
rect 56042 8372 56048 8384
rect 56100 8372 56106 8424
rect 57974 8412 57980 8424
rect 57935 8384 57980 8412
rect 57974 8372 57980 8384
rect 58032 8372 58038 8424
rect 55766 8344 55772 8356
rect 55508 8316 55772 8344
rect 55766 8304 55772 8316
rect 55824 8344 55830 8356
rect 56134 8344 56140 8356
rect 55824 8316 56140 8344
rect 55824 8304 55830 8316
rect 56134 8304 56140 8316
rect 56192 8304 56198 8356
rect 57241 8347 57299 8353
rect 57241 8313 57253 8347
rect 57287 8344 57299 8347
rect 57514 8344 57520 8356
rect 57287 8316 57520 8344
rect 57287 8313 57299 8316
rect 57241 8307 57299 8313
rect 57514 8304 57520 8316
rect 57572 8304 57578 8356
rect 1104 8186 58880 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 50326 8186
rect 50378 8134 50390 8186
rect 50442 8134 50454 8186
rect 50506 8134 50518 8186
rect 50570 8134 58880 8186
rect 1104 8112 58880 8134
rect 1854 8004 1860 8016
rect 1815 7976 1860 8004
rect 1854 7964 1860 7976
rect 1912 7964 1918 8016
rect 53653 7939 53711 7945
rect 53653 7905 53665 7939
rect 53699 7936 53711 7939
rect 55122 7936 55128 7948
rect 53699 7908 55128 7936
rect 53699 7905 53711 7908
rect 53653 7899 53711 7905
rect 55122 7896 55128 7908
rect 55180 7896 55186 7948
rect 56778 7896 56784 7948
rect 56836 7936 56842 7948
rect 57149 7939 57207 7945
rect 57149 7936 57161 7939
rect 56836 7908 57161 7936
rect 56836 7896 56842 7908
rect 57149 7905 57161 7908
rect 57195 7905 57207 7939
rect 57330 7936 57336 7948
rect 57291 7908 57336 7936
rect 57149 7899 57207 7905
rect 57330 7896 57336 7908
rect 57388 7896 57394 7948
rect 2038 7800 2044 7812
rect 1999 7772 2044 7800
rect 2038 7760 2044 7772
rect 2096 7760 2102 7812
rect 54481 7803 54539 7809
rect 54481 7769 54493 7803
rect 54527 7800 54539 7803
rect 57330 7800 57336 7812
rect 54527 7772 57336 7800
rect 54527 7769 54539 7772
rect 54481 7763 54539 7769
rect 57330 7760 57336 7772
rect 57388 7760 57394 7812
rect 57514 7800 57520 7812
rect 57475 7772 57520 7800
rect 57514 7760 57520 7772
rect 57572 7760 57578 7812
rect 55125 7735 55183 7741
rect 55125 7701 55137 7735
rect 55171 7732 55183 7735
rect 55674 7732 55680 7744
rect 55171 7704 55680 7732
rect 55171 7701 55183 7704
rect 55125 7695 55183 7701
rect 55674 7692 55680 7704
rect 55732 7692 55738 7744
rect 55769 7735 55827 7741
rect 55769 7701 55781 7735
rect 55815 7732 55827 7735
rect 56226 7732 56232 7744
rect 55815 7704 56232 7732
rect 55815 7701 55827 7704
rect 55769 7695 55827 7701
rect 56226 7692 56232 7704
rect 56284 7692 56290 7744
rect 1104 7642 58880 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 58880 7642
rect 1104 7568 58880 7590
rect 52546 7488 52552 7540
rect 52604 7528 52610 7540
rect 52604 7500 57560 7528
rect 52604 7488 52610 7500
rect 55769 7463 55827 7469
rect 55769 7429 55781 7463
rect 55815 7429 55827 7463
rect 55769 7423 55827 7429
rect 55214 7392 55220 7404
rect 52932 7364 55220 7392
rect 52932 7333 52960 7364
rect 55214 7352 55220 7364
rect 55272 7352 55278 7404
rect 55784 7392 55812 7423
rect 57532 7401 57560 7500
rect 56597 7395 56655 7401
rect 56597 7392 56609 7395
rect 55784 7364 56609 7392
rect 56597 7361 56609 7364
rect 56643 7361 56655 7395
rect 56597 7355 56655 7361
rect 57517 7395 57575 7401
rect 57517 7361 57529 7395
rect 57563 7361 57575 7395
rect 57517 7355 57575 7361
rect 52917 7327 52975 7333
rect 52917 7293 52929 7327
rect 52963 7293 52975 7327
rect 52917 7287 52975 7293
rect 54665 7327 54723 7333
rect 54665 7293 54677 7327
rect 54711 7293 54723 7327
rect 54665 7287 54723 7293
rect 55309 7327 55367 7333
rect 55309 7293 55321 7327
rect 55355 7324 55367 7327
rect 55398 7324 55404 7336
rect 55355 7296 55404 7324
rect 55355 7293 55367 7296
rect 55309 7287 55367 7293
rect 54680 7256 54708 7287
rect 55398 7284 55404 7296
rect 55456 7284 55462 7336
rect 55582 7284 55588 7336
rect 55640 7324 55646 7336
rect 55953 7327 56011 7333
rect 55953 7324 55965 7327
rect 55640 7296 55965 7324
rect 55640 7284 55646 7296
rect 55953 7293 55965 7296
rect 55999 7324 56011 7327
rect 56410 7324 56416 7336
rect 55999 7296 56272 7324
rect 56371 7296 56416 7324
rect 55999 7293 56011 7296
rect 55953 7287 56011 7293
rect 56042 7256 56048 7268
rect 54680 7228 56048 7256
rect 56042 7216 56048 7228
rect 56100 7216 56106 7268
rect 56244 7256 56272 7296
rect 56410 7284 56416 7296
rect 56468 7284 56474 7336
rect 57698 7324 57704 7336
rect 57659 7296 57704 7324
rect 57698 7284 57704 7296
rect 57756 7284 57762 7336
rect 57238 7256 57244 7268
rect 56244 7228 57244 7256
rect 57238 7216 57244 7228
rect 57296 7216 57302 7268
rect 55674 7148 55680 7200
rect 55732 7188 55738 7200
rect 56502 7188 56508 7200
rect 55732 7160 56508 7188
rect 55732 7148 55738 7160
rect 56502 7148 56508 7160
rect 56560 7148 56566 7200
rect 57057 7191 57115 7197
rect 57057 7157 57069 7191
rect 57103 7188 57115 7191
rect 57974 7188 57980 7200
rect 57103 7160 57980 7188
rect 57103 7157 57115 7160
rect 57057 7151 57115 7157
rect 57974 7148 57980 7160
rect 58032 7148 58038 7200
rect 58066 7148 58072 7200
rect 58124 7188 58130 7200
rect 58161 7191 58219 7197
rect 58161 7188 58173 7191
rect 58124 7160 58173 7188
rect 58124 7148 58130 7160
rect 58161 7157 58173 7160
rect 58207 7157 58219 7191
rect 58161 7151 58219 7157
rect 1104 7098 58880 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 50326 7098
rect 50378 7046 50390 7098
rect 50442 7046 50454 7098
rect 50506 7046 50518 7098
rect 50570 7046 58880 7098
rect 1104 7024 58880 7046
rect 57054 6984 57060 6996
rect 55232 6956 57060 6984
rect 53742 6876 53748 6928
rect 53800 6916 53806 6928
rect 55232 6916 55260 6956
rect 57054 6944 57060 6956
rect 57112 6944 57118 6996
rect 53800 6888 55260 6916
rect 53800 6876 53806 6888
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 14642 6848 14648 6860
rect 1903 6820 14648 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 51721 6851 51779 6857
rect 51721 6817 51733 6851
rect 51767 6817 51779 6851
rect 52546 6848 52552 6860
rect 52507 6820 52552 6848
rect 51721 6811 51779 6817
rect 2038 6780 2044 6792
rect 1999 6752 2044 6780
rect 2038 6740 2044 6752
rect 2096 6740 2102 6792
rect 51736 6712 51764 6811
rect 52546 6808 52552 6820
rect 52604 6808 52610 6860
rect 55148 6857 55176 6888
rect 55125 6851 55183 6857
rect 55125 6817 55137 6851
rect 55171 6817 55183 6851
rect 55766 6848 55772 6860
rect 55727 6820 55772 6848
rect 55125 6811 55183 6817
rect 55766 6808 55772 6820
rect 55824 6808 55830 6860
rect 57974 6848 57980 6860
rect 57935 6820 57980 6848
rect 57974 6808 57980 6820
rect 58032 6808 58038 6860
rect 58158 6848 58164 6860
rect 58119 6820 58164 6848
rect 58158 6808 58164 6820
rect 58216 6808 58222 6860
rect 53193 6783 53251 6789
rect 53193 6749 53205 6783
rect 53239 6780 53251 6783
rect 56781 6783 56839 6789
rect 56781 6780 56793 6783
rect 53239 6752 56793 6780
rect 53239 6749 53251 6752
rect 53193 6743 53251 6749
rect 56781 6749 56793 6752
rect 56827 6749 56839 6783
rect 56781 6743 56839 6749
rect 56965 6783 57023 6789
rect 56965 6749 56977 6783
rect 57011 6749 57023 6783
rect 56965 6743 57023 6749
rect 55490 6712 55496 6724
rect 51736 6684 55496 6712
rect 55490 6672 55496 6684
rect 55548 6672 55554 6724
rect 55585 6715 55643 6721
rect 55585 6681 55597 6715
rect 55631 6712 55643 6715
rect 56980 6712 57008 6743
rect 55631 6684 57008 6712
rect 55631 6681 55643 6684
rect 55585 6675 55643 6681
rect 53837 6647 53895 6653
rect 53837 6613 53849 6647
rect 53883 6644 53895 6647
rect 54294 6644 54300 6656
rect 53883 6616 54300 6644
rect 53883 6613 53895 6616
rect 53837 6607 53895 6613
rect 54294 6604 54300 6616
rect 54352 6604 54358 6656
rect 54478 6644 54484 6656
rect 54439 6616 54484 6644
rect 54478 6604 54484 6616
rect 54536 6604 54542 6656
rect 54941 6647 54999 6653
rect 54941 6613 54953 6647
rect 54987 6644 54999 6647
rect 55858 6644 55864 6656
rect 54987 6616 55864 6644
rect 54987 6613 54999 6616
rect 54941 6607 54999 6613
rect 55858 6604 55864 6616
rect 55916 6604 55922 6656
rect 56134 6604 56140 6656
rect 56192 6644 56198 6656
rect 57149 6647 57207 6653
rect 57149 6644 57161 6647
rect 56192 6616 57161 6644
rect 56192 6604 56198 6616
rect 57149 6613 57161 6616
rect 57195 6613 57207 6647
rect 57149 6607 57207 6613
rect 1104 6554 58880 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 58880 6554
rect 1104 6480 58880 6502
rect 55401 6443 55459 6449
rect 55401 6409 55413 6443
rect 55447 6440 55459 6443
rect 57698 6440 57704 6452
rect 55447 6412 57704 6440
rect 55447 6409 55459 6412
rect 55401 6403 55459 6409
rect 57698 6400 57704 6412
rect 57756 6400 57762 6452
rect 52454 6332 52460 6384
rect 52512 6372 52518 6384
rect 56321 6375 56379 6381
rect 52512 6344 56180 6372
rect 52512 6332 52518 6344
rect 55490 6304 55496 6316
rect 52472 6276 55496 6304
rect 51629 6239 51687 6245
rect 51629 6205 51641 6239
rect 51675 6236 51687 6239
rect 52362 6236 52368 6248
rect 51675 6208 52368 6236
rect 51675 6205 51687 6208
rect 51629 6199 51687 6205
rect 52362 6196 52368 6208
rect 52420 6196 52426 6248
rect 52472 6245 52500 6276
rect 55490 6264 55496 6276
rect 55548 6264 55554 6316
rect 56152 6304 56180 6344
rect 56321 6341 56333 6375
rect 56367 6372 56379 6375
rect 56410 6372 56416 6384
rect 56367 6344 56416 6372
rect 56367 6341 56379 6344
rect 56321 6335 56379 6341
rect 56410 6332 56416 6344
rect 56468 6332 56474 6384
rect 56594 6332 56600 6384
rect 56652 6372 56658 6384
rect 57422 6372 57428 6384
rect 56652 6344 57428 6372
rect 56652 6332 56658 6344
rect 57422 6332 57428 6344
rect 57480 6332 57486 6384
rect 56152 6276 56456 6304
rect 52457 6239 52515 6245
rect 52457 6205 52469 6239
rect 52503 6205 52515 6239
rect 52457 6199 52515 6205
rect 53101 6239 53159 6245
rect 53101 6205 53113 6239
rect 53147 6205 53159 6239
rect 53101 6199 53159 6205
rect 53116 6168 53144 6199
rect 54018 6196 54024 6248
rect 54076 6236 54082 6248
rect 54205 6239 54263 6245
rect 54205 6236 54217 6239
rect 54076 6208 54217 6236
rect 54076 6196 54082 6208
rect 54205 6205 54217 6208
rect 54251 6205 54263 6239
rect 54938 6236 54944 6248
rect 54899 6208 54944 6236
rect 54205 6199 54263 6205
rect 54938 6196 54944 6208
rect 54996 6196 55002 6248
rect 55582 6236 55588 6248
rect 55543 6208 55588 6236
rect 55582 6196 55588 6208
rect 55640 6196 55646 6248
rect 56134 6236 56140 6248
rect 56095 6208 56140 6236
rect 56134 6196 56140 6208
rect 56192 6196 56198 6248
rect 56428 6236 56456 6276
rect 56502 6264 56508 6316
rect 56560 6304 56566 6316
rect 56781 6307 56839 6313
rect 56781 6304 56793 6307
rect 56560 6276 56793 6304
rect 56560 6264 56566 6276
rect 56781 6273 56793 6276
rect 56827 6273 56839 6307
rect 56781 6267 56839 6273
rect 56962 6236 56968 6248
rect 56428 6208 56824 6236
rect 56923 6208 56968 6236
rect 56686 6168 56692 6180
rect 53116 6140 56692 6168
rect 56686 6128 56692 6140
rect 56744 6128 56750 6180
rect 56796 6168 56824 6208
rect 56962 6196 56968 6208
rect 57020 6196 57026 6248
rect 57146 6168 57152 6180
rect 56796 6140 57152 6168
rect 57146 6128 57152 6140
rect 57204 6128 57210 6180
rect 57425 6171 57483 6177
rect 57425 6137 57437 6171
rect 57471 6168 57483 6171
rect 57977 6171 58035 6177
rect 57977 6168 57989 6171
rect 57471 6140 57989 6168
rect 57471 6137 57483 6140
rect 57425 6131 57483 6137
rect 57977 6137 57989 6140
rect 58023 6137 58035 6171
rect 57977 6131 58035 6137
rect 54754 6100 54760 6112
rect 54715 6072 54760 6100
rect 54754 6060 54760 6072
rect 54812 6060 54818 6112
rect 55858 6060 55864 6112
rect 55916 6100 55922 6112
rect 57238 6100 57244 6112
rect 55916 6072 57244 6100
rect 55916 6060 55922 6072
rect 57238 6060 57244 6072
rect 57296 6060 57302 6112
rect 57882 6060 57888 6112
rect 57940 6100 57946 6112
rect 58069 6103 58127 6109
rect 58069 6100 58081 6103
rect 57940 6072 58081 6100
rect 57940 6060 57946 6072
rect 58069 6069 58081 6072
rect 58115 6069 58127 6103
rect 58069 6063 58127 6069
rect 1104 6010 58880 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 50326 6010
rect 50378 5958 50390 6010
rect 50442 5958 50454 6010
rect 50506 5958 50518 6010
rect 50570 5958 58880 6010
rect 1104 5936 58880 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 54849 5899 54907 5905
rect 54849 5865 54861 5899
rect 54895 5896 54907 5899
rect 56962 5896 56968 5908
rect 54895 5868 56968 5896
rect 54895 5865 54907 5868
rect 54849 5859 54907 5865
rect 56962 5856 56968 5868
rect 57020 5856 57026 5908
rect 1854 5828 1860 5840
rect 1815 5800 1860 5828
rect 1854 5788 1860 5800
rect 1912 5788 1918 5840
rect 55674 5828 55680 5840
rect 48286 5800 53788 5828
rect 29546 5720 29552 5772
rect 29604 5760 29610 5772
rect 48286 5760 48314 5800
rect 53760 5772 53788 5800
rect 55048 5800 55680 5828
rect 52454 5760 52460 5772
rect 29604 5732 48314 5760
rect 52415 5732 52460 5760
rect 29604 5720 29610 5732
rect 52454 5720 52460 5732
rect 52512 5720 52518 5772
rect 53742 5760 53748 5772
rect 53703 5732 53748 5760
rect 53742 5720 53748 5732
rect 53800 5720 53806 5772
rect 55048 5769 55076 5800
rect 55674 5788 55680 5800
rect 55732 5788 55738 5840
rect 55769 5831 55827 5837
rect 55769 5797 55781 5831
rect 55815 5828 55827 5831
rect 57606 5828 57612 5840
rect 55815 5800 57612 5828
rect 55815 5797 55827 5800
rect 55769 5791 55827 5797
rect 57606 5788 57612 5800
rect 57664 5788 57670 5840
rect 58158 5828 58164 5840
rect 58119 5800 58164 5828
rect 58158 5788 58164 5800
rect 58216 5788 58222 5840
rect 54389 5763 54447 5769
rect 54389 5729 54401 5763
rect 54435 5760 54447 5763
rect 55033 5763 55091 5769
rect 55033 5760 55045 5763
rect 54435 5732 55045 5760
rect 54435 5729 54447 5732
rect 54389 5723 54447 5729
rect 55033 5729 55045 5732
rect 55079 5729 55091 5763
rect 55033 5723 55091 5729
rect 55585 5763 55643 5769
rect 55585 5729 55597 5763
rect 55631 5760 55643 5763
rect 56502 5760 56508 5772
rect 55631 5732 56508 5760
rect 55631 5729 55643 5732
rect 55585 5723 55643 5729
rect 56502 5720 56508 5732
rect 56560 5720 56566 5772
rect 56686 5760 56692 5772
rect 56647 5732 56692 5760
rect 56686 5720 56692 5732
rect 56744 5720 56750 5772
rect 57977 5763 58035 5769
rect 57977 5729 57989 5763
rect 58023 5760 58035 5763
rect 58066 5760 58072 5772
rect 58023 5732 58072 5760
rect 58023 5729 58035 5732
rect 57977 5723 58035 5729
rect 58066 5720 58072 5732
rect 58124 5720 58130 5772
rect 51813 5695 51871 5701
rect 51813 5661 51825 5695
rect 51859 5692 51871 5695
rect 56778 5692 56784 5704
rect 51859 5664 56784 5692
rect 51859 5661 51871 5664
rect 51813 5655 51871 5661
rect 56778 5652 56784 5664
rect 56836 5652 56842 5704
rect 56873 5695 56931 5701
rect 56873 5661 56885 5695
rect 56919 5661 56931 5695
rect 56873 5655 56931 5661
rect 54205 5627 54263 5633
rect 54205 5593 54217 5627
rect 54251 5624 54263 5627
rect 56888 5624 56916 5655
rect 54251 5596 56916 5624
rect 54251 5593 54263 5596
rect 54205 5587 54263 5593
rect 14734 5516 14740 5568
rect 14792 5556 14798 5568
rect 15010 5556 15016 5568
rect 14792 5528 15016 5556
rect 14792 5516 14798 5528
rect 15010 5516 15016 5528
rect 15068 5556 15074 5568
rect 29546 5556 29552 5568
rect 15068 5528 29552 5556
rect 15068 5516 15074 5528
rect 29546 5516 29552 5528
rect 29604 5516 29610 5568
rect 53098 5556 53104 5568
rect 53059 5528 53104 5556
rect 53098 5516 53104 5528
rect 53156 5516 53162 5568
rect 53561 5559 53619 5565
rect 53561 5525 53573 5559
rect 53607 5556 53619 5559
rect 56870 5556 56876 5568
rect 53607 5528 56876 5556
rect 53607 5525 53619 5528
rect 53561 5519 53619 5525
rect 56870 5516 56876 5528
rect 56928 5516 56934 5568
rect 57054 5556 57060 5568
rect 57015 5528 57060 5556
rect 57054 5516 57060 5528
rect 57112 5516 57118 5568
rect 1104 5466 58880 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 58880 5466
rect 1104 5392 58880 5414
rect 53190 5312 53196 5364
rect 53248 5352 53254 5364
rect 54205 5355 54263 5361
rect 54205 5352 54217 5355
rect 53248 5324 54217 5352
rect 53248 5312 53254 5324
rect 54205 5321 54217 5324
rect 54251 5352 54263 5355
rect 54938 5352 54944 5364
rect 54251 5324 54944 5352
rect 54251 5321 54263 5324
rect 54205 5315 54263 5321
rect 54938 5312 54944 5324
rect 54996 5312 55002 5364
rect 50982 5176 50988 5228
rect 51040 5216 51046 5228
rect 54941 5219 54999 5225
rect 51040 5188 54800 5216
rect 51040 5176 51046 5188
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 2130 5148 2136 5160
rect 1903 5120 2136 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 49789 5151 49847 5157
rect 49789 5117 49801 5151
rect 49835 5148 49847 5151
rect 49970 5148 49976 5160
rect 49835 5120 49976 5148
rect 49835 5117 49847 5120
rect 49789 5111 49847 5117
rect 49970 5108 49976 5120
rect 50028 5108 50034 5160
rect 50614 5148 50620 5160
rect 50575 5120 50620 5148
rect 50614 5108 50620 5120
rect 50672 5108 50678 5160
rect 51626 5148 51632 5160
rect 51587 5120 51632 5148
rect 51626 5108 51632 5120
rect 51684 5108 51690 5160
rect 52454 5148 52460 5160
rect 52415 5120 52460 5148
rect 52454 5108 52460 5120
rect 52512 5108 52518 5160
rect 54772 5157 54800 5188
rect 54941 5185 54953 5219
rect 54987 5216 54999 5219
rect 55950 5216 55956 5228
rect 54987 5188 55956 5216
rect 54987 5185 54999 5188
rect 54941 5179 54999 5185
rect 53101 5151 53159 5157
rect 53101 5117 53113 5151
rect 53147 5117 53159 5151
rect 53101 5111 53159 5117
rect 54021 5151 54079 5157
rect 54021 5117 54033 5151
rect 54067 5117 54079 5151
rect 54021 5111 54079 5117
rect 54757 5151 54815 5157
rect 54757 5117 54769 5151
rect 54803 5117 54815 5151
rect 54757 5111 54815 5117
rect 51902 5040 51908 5092
rect 51960 5080 51966 5092
rect 53116 5080 53144 5111
rect 51960 5052 53144 5080
rect 54036 5080 54064 5111
rect 54956 5080 54984 5179
rect 55950 5176 55956 5188
rect 56008 5176 56014 5228
rect 57330 5176 57336 5228
rect 57388 5216 57394 5228
rect 57517 5219 57575 5225
rect 57517 5216 57529 5219
rect 57388 5188 57529 5216
rect 57388 5176 57394 5188
rect 57517 5185 57529 5188
rect 57563 5185 57575 5219
rect 57517 5179 57575 5185
rect 56873 5151 56931 5157
rect 56873 5117 56885 5151
rect 56919 5148 56931 5151
rect 57054 5148 57060 5160
rect 56919 5120 57060 5148
rect 56919 5117 56931 5120
rect 56873 5111 56931 5117
rect 57054 5108 57060 5120
rect 57112 5108 57118 5160
rect 57698 5148 57704 5160
rect 57659 5120 57704 5148
rect 57698 5108 57704 5120
rect 57756 5108 57762 5160
rect 55858 5080 55864 5092
rect 54036 5052 54984 5080
rect 55819 5052 55864 5080
rect 51960 5040 51966 5052
rect 55858 5040 55864 5052
rect 55916 5040 55922 5092
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 52917 5015 52975 5021
rect 52917 4981 52929 5015
rect 52963 5012 52975 5015
rect 53282 5012 53288 5024
rect 52963 4984 53288 5012
rect 52963 4981 52975 4984
rect 52917 4975 52975 4981
rect 53282 4972 53288 4984
rect 53340 4972 53346 5024
rect 55766 4972 55772 5024
rect 55824 5012 55830 5024
rect 55953 5015 56011 5021
rect 55953 5012 55965 5015
rect 55824 4984 55965 5012
rect 55824 4972 55830 4984
rect 55953 4981 55965 4984
rect 55999 4981 56011 5015
rect 55953 4975 56011 4981
rect 56965 5015 57023 5021
rect 56965 4981 56977 5015
rect 57011 5012 57023 5015
rect 57054 5012 57060 5024
rect 57011 4984 57060 5012
rect 57011 4981 57023 4984
rect 56965 4975 57023 4981
rect 57054 4972 57060 4984
rect 57112 4972 57118 5024
rect 58158 5012 58164 5024
rect 58119 4984 58164 5012
rect 58158 4972 58164 4984
rect 58216 4972 58222 5024
rect 1104 4922 58880 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 50326 4922
rect 50378 4870 50390 4922
rect 50442 4870 50454 4922
rect 50506 4870 50518 4922
rect 50570 4870 58880 4922
rect 1104 4848 58880 4870
rect 56686 4808 56692 4820
rect 53760 4780 56692 4808
rect 53760 4749 53788 4780
rect 56686 4768 56692 4780
rect 56744 4768 56750 4820
rect 53745 4743 53803 4749
rect 53745 4709 53757 4743
rect 53791 4709 53803 4743
rect 53745 4703 53803 4709
rect 54481 4743 54539 4749
rect 54481 4709 54493 4743
rect 54527 4740 54539 4743
rect 56410 4740 56416 4752
rect 54527 4712 56416 4740
rect 54527 4709 54539 4712
rect 54481 4703 54539 4709
rect 56410 4700 56416 4712
rect 56468 4700 56474 4752
rect 56873 4743 56931 4749
rect 56873 4709 56885 4743
rect 56919 4740 56931 4743
rect 58158 4740 58164 4752
rect 56919 4712 58164 4740
rect 56919 4709 56931 4712
rect 56873 4703 56931 4709
rect 58158 4700 58164 4712
rect 58216 4700 58222 4752
rect 37366 4632 37372 4684
rect 37424 4672 37430 4684
rect 37921 4675 37979 4681
rect 37921 4672 37933 4675
rect 37424 4644 37933 4672
rect 37424 4632 37430 4644
rect 37921 4641 37933 4644
rect 37967 4641 37979 4675
rect 37921 4635 37979 4641
rect 48961 4675 49019 4681
rect 48961 4641 48973 4675
rect 49007 4672 49019 4675
rect 49142 4672 49148 4684
rect 49007 4644 49148 4672
rect 49007 4641 49019 4644
rect 48961 4635 49019 4641
rect 49142 4632 49148 4644
rect 49200 4632 49206 4684
rect 51902 4672 51908 4684
rect 51863 4644 51908 4672
rect 51902 4632 51908 4644
rect 51960 4632 51966 4684
rect 52549 4675 52607 4681
rect 52549 4641 52561 4675
rect 52595 4672 52607 4675
rect 53190 4672 53196 4684
rect 52595 4644 53196 4672
rect 52595 4641 52607 4644
rect 52549 4635 52607 4641
rect 53190 4632 53196 4644
rect 53248 4632 53254 4684
rect 54570 4632 54576 4684
rect 54628 4672 54634 4684
rect 55309 4675 55367 4681
rect 55309 4672 55321 4675
rect 54628 4644 55321 4672
rect 54628 4632 54634 4644
rect 55309 4641 55321 4644
rect 55355 4641 55367 4675
rect 55309 4635 55367 4641
rect 56594 4632 56600 4684
rect 56652 4672 56658 4684
rect 57701 4675 57759 4681
rect 57701 4672 57713 4675
rect 56652 4644 57713 4672
rect 56652 4632 56658 4644
rect 57701 4641 57713 4644
rect 57747 4641 57759 4675
rect 57701 4635 57759 4641
rect 54294 4564 54300 4616
rect 54352 4604 54358 4616
rect 55125 4607 55183 4613
rect 55125 4604 55137 4607
rect 54352 4576 55137 4604
rect 54352 4564 54358 4576
rect 55125 4573 55137 4576
rect 55171 4573 55183 4607
rect 55125 4567 55183 4573
rect 56778 4564 56784 4616
rect 56836 4604 56842 4616
rect 57517 4607 57575 4613
rect 57517 4604 57529 4607
rect 56836 4576 57529 4604
rect 56836 4564 56842 4576
rect 57517 4573 57529 4576
rect 57563 4573 57575 4607
rect 57517 4567 57575 4573
rect 46385 4539 46443 4545
rect 46385 4505 46397 4539
rect 46431 4536 46443 4539
rect 46934 4536 46940 4548
rect 46431 4508 46940 4536
rect 46431 4505 46443 4508
rect 46385 4499 46443 4505
rect 46934 4496 46940 4508
rect 46992 4496 46998 4548
rect 53009 4539 53067 4545
rect 53009 4505 53021 4539
rect 53055 4536 53067 4539
rect 55030 4536 55036 4548
rect 53055 4508 55036 4536
rect 53055 4505 53067 4508
rect 53009 4499 53067 4505
rect 55030 4496 55036 4508
rect 55088 4496 55094 4548
rect 32953 4471 33011 4477
rect 32953 4437 32965 4471
rect 32999 4468 33011 4471
rect 33594 4468 33600 4480
rect 32999 4440 33600 4468
rect 32999 4437 33011 4440
rect 32953 4431 33011 4437
rect 33594 4428 33600 4440
rect 33652 4428 33658 4480
rect 36081 4471 36139 4477
rect 36081 4437 36093 4471
rect 36127 4468 36139 4471
rect 36262 4468 36268 4480
rect 36127 4440 36268 4468
rect 36127 4437 36139 4440
rect 36081 4431 36139 4437
rect 36262 4428 36268 4440
rect 36320 4428 36326 4480
rect 37001 4471 37059 4477
rect 37001 4437 37013 4471
rect 37047 4468 37059 4471
rect 37274 4468 37280 4480
rect 37047 4440 37280 4468
rect 37047 4437 37059 4440
rect 37001 4431 37059 4437
rect 37274 4428 37280 4440
rect 37332 4428 37338 4480
rect 37737 4471 37795 4477
rect 37737 4437 37749 4471
rect 37783 4468 37795 4471
rect 38378 4468 38384 4480
rect 37783 4440 38384 4468
rect 37783 4437 37795 4440
rect 37737 4431 37795 4437
rect 38378 4428 38384 4440
rect 38436 4428 38442 4480
rect 38562 4468 38568 4480
rect 38523 4440 38568 4468
rect 38562 4428 38568 4440
rect 38620 4428 38626 4480
rect 39209 4471 39267 4477
rect 39209 4437 39221 4471
rect 39255 4468 39267 4471
rect 39390 4468 39396 4480
rect 39255 4440 39396 4468
rect 39255 4437 39267 4440
rect 39209 4431 39267 4437
rect 39390 4428 39396 4440
rect 39448 4428 39454 4480
rect 39482 4428 39488 4480
rect 39540 4468 39546 4480
rect 39853 4471 39911 4477
rect 39853 4468 39865 4471
rect 39540 4440 39865 4468
rect 39540 4428 39546 4440
rect 39853 4437 39865 4440
rect 39899 4437 39911 4471
rect 41506 4468 41512 4480
rect 41467 4440 41512 4468
rect 39853 4431 39911 4437
rect 41506 4428 41512 4440
rect 41564 4428 41570 4480
rect 42334 4468 42340 4480
rect 42295 4440 42340 4468
rect 42334 4428 42340 4440
rect 42392 4428 42398 4480
rect 43438 4468 43444 4480
rect 43399 4440 43444 4468
rect 43438 4428 43444 4440
rect 43496 4428 43502 4480
rect 47026 4468 47032 4480
rect 46987 4440 47032 4468
rect 47026 4428 47032 4440
rect 47084 4428 47090 4480
rect 48038 4468 48044 4480
rect 47999 4440 48044 4468
rect 48038 4428 48044 4440
rect 48096 4428 48102 4480
rect 48777 4471 48835 4477
rect 48777 4437 48789 4471
rect 48823 4468 48835 4471
rect 48958 4468 48964 4480
rect 48823 4440 48964 4468
rect 48823 4437 48835 4440
rect 48777 4431 48835 4437
rect 48958 4428 48964 4440
rect 49016 4428 49022 4480
rect 49050 4428 49056 4480
rect 49108 4468 49114 4480
rect 49605 4471 49663 4477
rect 49605 4468 49617 4471
rect 49108 4440 49617 4468
rect 49108 4428 49114 4440
rect 49605 4437 49617 4440
rect 49651 4437 49663 4471
rect 49605 4431 49663 4437
rect 49694 4428 49700 4480
rect 49752 4468 49758 4480
rect 50249 4471 50307 4477
rect 50249 4468 50261 4471
rect 49752 4440 50261 4468
rect 49752 4428 49758 4440
rect 50249 4437 50261 4440
rect 50295 4437 50307 4471
rect 51718 4468 51724 4480
rect 51679 4440 51724 4468
rect 50249 4431 50307 4437
rect 51718 4428 51724 4440
rect 51776 4428 51782 4480
rect 52365 4471 52423 4477
rect 52365 4437 52377 4471
rect 52411 4468 52423 4471
rect 53742 4468 53748 4480
rect 52411 4440 53748 4468
rect 52411 4437 52423 4440
rect 52365 4431 52423 4437
rect 53742 4428 53748 4440
rect 53800 4428 53806 4480
rect 53837 4471 53895 4477
rect 53837 4437 53849 4471
rect 53883 4468 53895 4471
rect 54386 4468 54392 4480
rect 53883 4440 54392 4468
rect 53883 4437 53895 4440
rect 53837 4431 53895 4437
rect 54386 4428 54392 4440
rect 54444 4428 54450 4480
rect 54573 4471 54631 4477
rect 54573 4437 54585 4471
rect 54619 4468 54631 4471
rect 55306 4468 55312 4480
rect 54619 4440 55312 4468
rect 54619 4437 54631 4440
rect 54573 4431 54631 4437
rect 55306 4428 55312 4440
rect 55364 4428 55370 4480
rect 55582 4468 55588 4480
rect 55543 4440 55588 4468
rect 55582 4428 55588 4440
rect 55640 4428 55646 4480
rect 56962 4468 56968 4480
rect 56923 4440 56968 4468
rect 56962 4428 56968 4440
rect 57020 4428 57026 4480
rect 57974 4468 57980 4480
rect 57935 4440 57980 4468
rect 57974 4428 57980 4440
rect 58032 4428 58038 4480
rect 1104 4378 58880 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 58880 4378
rect 1104 4304 58880 4326
rect 34790 4196 34796 4208
rect 34751 4168 34796 4196
rect 34790 4156 34796 4168
rect 34848 4156 34854 4208
rect 44266 4156 44272 4208
rect 44324 4196 44330 4208
rect 45097 4199 45155 4205
rect 45097 4196 45109 4199
rect 44324 4168 45109 4196
rect 44324 4156 44330 4168
rect 45097 4165 45109 4168
rect 45143 4165 45155 4199
rect 45738 4196 45744 4208
rect 45699 4168 45744 4196
rect 45097 4159 45155 4165
rect 45738 4156 45744 4168
rect 45796 4156 45802 4208
rect 54386 4156 54392 4208
rect 54444 4196 54450 4208
rect 54444 4168 57008 4196
rect 54444 4156 54450 4168
rect 2038 4128 2044 4140
rect 1999 4100 2044 4128
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 49881 4131 49939 4137
rect 49881 4128 49893 4131
rect 47688 4100 49893 4128
rect 47688 4072 47716 4100
rect 49881 4097 49893 4100
rect 49927 4128 49939 4131
rect 49927 4100 50384 4128
rect 49927 4097 49939 4100
rect 49881 4091 49939 4097
rect 30006 4020 30012 4072
rect 30064 4060 30070 4072
rect 30285 4063 30343 4069
rect 30285 4060 30297 4063
rect 30064 4032 30297 4060
rect 30064 4020 30070 4032
rect 30285 4029 30297 4032
rect 30331 4029 30343 4063
rect 30285 4023 30343 4029
rect 32125 4063 32183 4069
rect 32125 4029 32137 4063
rect 32171 4060 32183 4063
rect 33042 4060 33048 4072
rect 32171 4032 33048 4060
rect 32171 4029 32183 4032
rect 32125 4023 32183 4029
rect 33042 4020 33048 4032
rect 33100 4020 33106 4072
rect 33229 4063 33287 4069
rect 33229 4029 33241 4063
rect 33275 4060 33287 4063
rect 34149 4063 34207 4069
rect 34149 4060 34161 4063
rect 33275 4032 34161 4060
rect 33275 4029 33287 4032
rect 33229 4023 33287 4029
rect 34149 4029 34161 4032
rect 34195 4060 34207 4063
rect 34195 4032 34928 4060
rect 34195 4029 34207 4032
rect 34149 4023 34207 4029
rect 1857 3995 1915 4001
rect 1857 3961 1869 3995
rect 1903 3992 1915 3995
rect 13170 3992 13176 4004
rect 1903 3964 13176 3992
rect 1903 3961 1915 3964
rect 1857 3955 1915 3961
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 34900 3936 34928 4032
rect 35250 4020 35256 4072
rect 35308 4060 35314 4072
rect 35437 4063 35495 4069
rect 35437 4060 35449 4063
rect 35308 4032 35449 4060
rect 35308 4020 35314 4032
rect 35437 4029 35449 4032
rect 35483 4029 35495 4063
rect 36078 4060 36084 4072
rect 36039 4032 36084 4060
rect 35437 4023 35495 4029
rect 36078 4020 36084 4032
rect 36136 4020 36142 4072
rect 37366 4060 37372 4072
rect 37327 4032 37372 4060
rect 37366 4020 37372 4032
rect 37424 4060 37430 4072
rect 38841 4063 38899 4069
rect 38841 4060 38853 4063
rect 37424 4032 38853 4060
rect 37424 4020 37430 4032
rect 38841 4029 38853 4032
rect 38887 4060 38899 4063
rect 39945 4063 40003 4069
rect 39945 4060 39957 4063
rect 38887 4032 39957 4060
rect 38887 4029 38899 4032
rect 38841 4023 38899 4029
rect 39945 4029 39957 4032
rect 39991 4060 40003 4063
rect 40589 4063 40647 4069
rect 40589 4060 40601 4063
rect 39991 4032 40601 4060
rect 39991 4029 40003 4032
rect 39945 4023 40003 4029
rect 40589 4029 40601 4032
rect 40635 4029 40647 4063
rect 41230 4060 41236 4072
rect 41191 4032 41236 4060
rect 40589 4023 40647 4029
rect 41230 4020 41236 4032
rect 41288 4020 41294 4072
rect 42061 4063 42119 4069
rect 42061 4029 42073 4063
rect 42107 4060 42119 4063
rect 42426 4060 42432 4072
rect 42107 4032 42432 4060
rect 42107 4029 42119 4032
rect 42061 4023 42119 4029
rect 42426 4020 42432 4032
rect 42484 4060 42490 4072
rect 43717 4063 43775 4069
rect 43717 4060 43729 4063
rect 42484 4032 43729 4060
rect 42484 4020 42490 4032
rect 43717 4029 43729 4032
rect 43763 4060 43775 4063
rect 43898 4060 43904 4072
rect 43763 4032 43904 4060
rect 43763 4029 43775 4032
rect 43717 4023 43775 4029
rect 43898 4020 43904 4032
rect 43956 4060 43962 4072
rect 44453 4063 44511 4069
rect 44453 4060 44465 4063
rect 43956 4032 44465 4060
rect 43956 4020 43962 4032
rect 44453 4029 44465 4032
rect 44499 4029 44511 4063
rect 44453 4023 44511 4029
rect 46937 4063 46995 4069
rect 46937 4029 46949 4063
rect 46983 4029 46995 4063
rect 47670 4060 47676 4072
rect 47631 4032 47676 4060
rect 46937 4023 46995 4029
rect 46952 3992 46980 4023
rect 47670 4020 47676 4032
rect 47728 4020 47734 4072
rect 49142 4060 49148 4072
rect 49103 4032 49148 4060
rect 49142 4020 49148 4032
rect 49200 4020 49206 4072
rect 49786 4060 49792 4072
rect 49620 4032 49792 4060
rect 47210 3992 47216 4004
rect 46952 3964 47216 3992
rect 47210 3952 47216 3964
rect 47268 3992 47274 4004
rect 49160 3992 49188 4020
rect 47268 3964 49188 3992
rect 47268 3952 47274 3964
rect 33045 3927 33103 3933
rect 33045 3893 33057 3927
rect 33091 3924 33103 3927
rect 33778 3924 33784 3936
rect 33091 3896 33784 3924
rect 33091 3893 33103 3896
rect 33045 3887 33103 3893
rect 33778 3884 33784 3896
rect 33836 3884 33842 3936
rect 33965 3927 34023 3933
rect 33965 3893 33977 3927
rect 34011 3924 34023 3927
rect 34514 3924 34520 3936
rect 34011 3896 34520 3924
rect 34011 3893 34023 3896
rect 33965 3887 34023 3893
rect 34514 3884 34520 3896
rect 34572 3884 34578 3936
rect 34882 3884 34888 3936
rect 34940 3924 34946 3936
rect 36265 3927 36323 3933
rect 36265 3924 36277 3927
rect 34940 3896 36277 3924
rect 34940 3884 34946 3896
rect 36265 3893 36277 3896
rect 36311 3893 36323 3927
rect 36265 3887 36323 3893
rect 37185 3927 37243 3933
rect 37185 3893 37197 3927
rect 37231 3924 37243 3927
rect 37550 3924 37556 3936
rect 37231 3896 37556 3924
rect 37231 3893 37243 3896
rect 37185 3887 37243 3893
rect 37550 3884 37556 3896
rect 37608 3884 37614 3936
rect 38657 3927 38715 3933
rect 38657 3893 38669 3927
rect 38703 3924 38715 3927
rect 39574 3924 39580 3936
rect 38703 3896 39580 3924
rect 38703 3893 38715 3896
rect 38657 3887 38715 3893
rect 39574 3884 39580 3896
rect 39632 3884 39638 3936
rect 39758 3924 39764 3936
rect 39719 3896 39764 3924
rect 39758 3884 39764 3896
rect 39816 3884 39822 3936
rect 40402 3924 40408 3936
rect 40363 3896 40408 3924
rect 40402 3884 40408 3896
rect 40460 3884 40466 3936
rect 41874 3924 41880 3936
rect 41835 3896 41880 3924
rect 41874 3884 41880 3896
rect 41932 3884 41938 3936
rect 43533 3927 43591 3933
rect 43533 3893 43545 3927
rect 43579 3924 43591 3927
rect 43714 3924 43720 3936
rect 43579 3896 43720 3924
rect 43579 3893 43591 3896
rect 43533 3887 43591 3893
rect 43714 3884 43720 3896
rect 43772 3884 43778 3936
rect 44269 3927 44327 3933
rect 44269 3893 44281 3927
rect 44315 3924 44327 3927
rect 44450 3924 44456 3936
rect 44315 3896 44456 3924
rect 44315 3893 44327 3896
rect 44269 3887 44327 3893
rect 44450 3884 44456 3896
rect 44508 3884 44514 3936
rect 46753 3927 46811 3933
rect 46753 3893 46765 3927
rect 46799 3924 46811 3927
rect 47118 3924 47124 3936
rect 46799 3896 47124 3924
rect 46799 3893 46811 3896
rect 46753 3887 46811 3893
rect 47118 3884 47124 3896
rect 47176 3884 47182 3936
rect 47872 3933 47900 3964
rect 47857 3927 47915 3933
rect 47857 3893 47869 3927
rect 47903 3893 47915 3927
rect 47857 3887 47915 3893
rect 48961 3927 49019 3933
rect 48961 3893 48973 3927
rect 49007 3924 49019 3927
rect 49620 3924 49648 4032
rect 49786 4020 49792 4032
rect 49844 4020 49850 4072
rect 50356 4069 50384 4100
rect 55030 4088 55036 4140
rect 55088 4128 55094 4140
rect 56413 4131 56471 4137
rect 56413 4128 56425 4131
rect 55088 4100 56425 4128
rect 55088 4088 55094 4100
rect 56413 4097 56425 4100
rect 56459 4097 56471 4131
rect 56413 4091 56471 4097
rect 56502 4088 56508 4140
rect 56560 4128 56566 4140
rect 56873 4131 56931 4137
rect 56873 4128 56885 4131
rect 56560 4100 56885 4128
rect 56560 4088 56566 4100
rect 56873 4097 56885 4100
rect 56919 4097 56931 4131
rect 56980 4128 57008 4168
rect 58526 4128 58532 4140
rect 56980 4100 58532 4128
rect 56873 4091 56931 4097
rect 58526 4088 58532 4100
rect 58584 4088 58590 4140
rect 50341 4063 50399 4069
rect 50341 4029 50353 4063
rect 50387 4029 50399 4063
rect 50982 4060 50988 4072
rect 50341 4023 50399 4029
rect 50448 4032 50988 4060
rect 49697 3995 49755 4001
rect 49697 3961 49709 3995
rect 49743 3992 49755 3995
rect 50448 3992 50476 4032
rect 50982 4020 50988 4032
rect 51040 4020 51046 4072
rect 51169 4063 51227 4069
rect 51169 4029 51181 4063
rect 51215 4060 51227 4063
rect 51813 4063 51871 4069
rect 51813 4060 51825 4063
rect 51215 4032 51825 4060
rect 51215 4029 51227 4032
rect 51169 4023 51227 4029
rect 51813 4029 51825 4032
rect 51859 4060 51871 4063
rect 51902 4060 51908 4072
rect 51859 4032 51908 4060
rect 51859 4029 51871 4032
rect 51813 4023 51871 4029
rect 51184 3992 51212 4023
rect 51902 4020 51908 4032
rect 51960 4020 51966 4072
rect 52457 4063 52515 4069
rect 52457 4029 52469 4063
rect 52503 4060 52515 4063
rect 53101 4063 53159 4069
rect 53101 4060 53113 4063
rect 52503 4032 53113 4060
rect 52503 4029 52515 4032
rect 52457 4023 52515 4029
rect 53101 4029 53113 4032
rect 53147 4060 53159 4063
rect 53190 4060 53196 4072
rect 53147 4032 53196 4060
rect 53147 4029 53159 4032
rect 53101 4023 53159 4029
rect 53190 4020 53196 4032
rect 53248 4020 53254 4072
rect 54570 4060 54576 4072
rect 53944 4032 54576 4060
rect 53944 3992 53972 4032
rect 54570 4020 54576 4032
rect 54628 4020 54634 4072
rect 55674 4020 55680 4072
rect 55732 4060 55738 4072
rect 55769 4063 55827 4069
rect 55769 4060 55781 4063
rect 55732 4032 55781 4060
rect 55732 4020 55738 4032
rect 55769 4029 55781 4032
rect 55815 4029 55827 4063
rect 56226 4060 56232 4072
rect 56187 4032 56232 4060
rect 55769 4023 55827 4029
rect 56226 4020 56232 4032
rect 56284 4020 56290 4072
rect 57974 4060 57980 4072
rect 57935 4032 57980 4060
rect 57974 4020 57980 4032
rect 58032 4020 58038 4072
rect 54110 3992 54116 4004
rect 49743 3964 50476 3992
rect 50540 3964 51212 3992
rect 52932 3964 53972 3992
rect 54071 3964 54116 3992
rect 49743 3961 49755 3964
rect 49697 3955 49755 3961
rect 49007 3896 49648 3924
rect 49007 3893 49019 3896
rect 48961 3887 49019 3893
rect 49878 3884 49884 3936
rect 49936 3924 49942 3936
rect 50540 3933 50568 3964
rect 50525 3927 50583 3933
rect 50525 3924 50537 3927
rect 49936 3896 50537 3924
rect 49936 3884 49942 3896
rect 50525 3893 50537 3896
rect 50571 3893 50583 3927
rect 50525 3887 50583 3893
rect 50985 3927 51043 3933
rect 50985 3893 50997 3927
rect 51031 3924 51043 3927
rect 51534 3924 51540 3936
rect 51031 3896 51540 3924
rect 51031 3893 51043 3896
rect 50985 3887 51043 3893
rect 51534 3884 51540 3896
rect 51592 3884 51598 3936
rect 51629 3927 51687 3933
rect 51629 3893 51641 3927
rect 51675 3924 51687 3927
rect 51994 3924 52000 3936
rect 51675 3896 52000 3924
rect 51675 3893 51687 3896
rect 51629 3887 51687 3893
rect 51994 3884 52000 3896
rect 52052 3884 52058 3936
rect 52273 3927 52331 3933
rect 52273 3893 52285 3927
rect 52319 3924 52331 3927
rect 52822 3924 52828 3936
rect 52319 3896 52828 3924
rect 52319 3893 52331 3896
rect 52273 3887 52331 3893
rect 52822 3884 52828 3896
rect 52880 3884 52886 3936
rect 52932 3933 52960 3964
rect 54110 3952 54116 3964
rect 54168 3952 54174 4004
rect 54662 3952 54668 4004
rect 54720 3992 54726 4004
rect 54941 3995 54999 4001
rect 54941 3992 54953 3995
rect 54720 3964 54953 3992
rect 54720 3952 54726 3964
rect 54941 3961 54953 3964
rect 54987 3961 54999 3995
rect 58158 3992 58164 4004
rect 58119 3964 58164 3992
rect 54941 3955 54999 3961
rect 58158 3952 58164 3964
rect 58216 3952 58222 4004
rect 52917 3927 52975 3933
rect 52917 3893 52929 3927
rect 52963 3893 52975 3927
rect 52917 3887 52975 3893
rect 53926 3884 53932 3936
rect 53984 3924 53990 3936
rect 54205 3927 54263 3933
rect 54205 3924 54217 3927
rect 53984 3896 54217 3924
rect 53984 3884 53990 3896
rect 54205 3893 54217 3896
rect 54251 3893 54263 3927
rect 54205 3887 54263 3893
rect 54846 3884 54852 3936
rect 54904 3924 54910 3936
rect 55033 3927 55091 3933
rect 55033 3924 55045 3927
rect 54904 3896 55045 3924
rect 54904 3884 54910 3896
rect 55033 3893 55045 3896
rect 55079 3893 55091 3927
rect 55033 3887 55091 3893
rect 55585 3927 55643 3933
rect 55585 3893 55597 3927
rect 55631 3924 55643 3927
rect 56594 3924 56600 3936
rect 55631 3896 56600 3924
rect 55631 3893 55643 3896
rect 55585 3887 55643 3893
rect 56594 3884 56600 3896
rect 56652 3884 56658 3936
rect 1104 3834 58880 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 50326 3834
rect 50378 3782 50390 3834
rect 50442 3782 50454 3834
rect 50506 3782 50518 3834
rect 50570 3782 58880 3834
rect 1104 3760 58880 3782
rect 12345 3723 12403 3729
rect 12345 3720 12357 3723
rect 11348 3692 12357 3720
rect 1857 3655 1915 3661
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 7834 3652 7840 3664
rect 1903 3624 7840 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 11238 3652 11244 3664
rect 11199 3624 11244 3652
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 11348 3661 11376 3692
rect 12345 3689 12357 3692
rect 12391 3689 12403 3723
rect 12345 3683 12403 3689
rect 36909 3723 36967 3729
rect 36909 3689 36921 3723
rect 36955 3720 36967 3723
rect 37366 3720 37372 3732
rect 36955 3692 37372 3720
rect 36955 3689 36967 3692
rect 36909 3683 36967 3689
rect 37366 3680 37372 3692
rect 37424 3680 37430 3732
rect 43898 3720 43904 3732
rect 43859 3692 43904 3720
rect 43898 3680 43904 3692
rect 43956 3680 43962 3732
rect 53745 3723 53803 3729
rect 53745 3689 53757 3723
rect 53791 3720 53803 3723
rect 54110 3720 54116 3732
rect 53791 3692 54116 3720
rect 53791 3689 53803 3692
rect 53745 3683 53803 3689
rect 54110 3680 54116 3692
rect 54168 3680 54174 3732
rect 56689 3723 56747 3729
rect 56689 3689 56701 3723
rect 56735 3720 56747 3723
rect 57698 3720 57704 3732
rect 56735 3692 57704 3720
rect 56735 3689 56747 3692
rect 56689 3683 56747 3689
rect 57698 3680 57704 3692
rect 57756 3680 57762 3732
rect 11333 3655 11391 3661
rect 11333 3621 11345 3655
rect 11379 3621 11391 3655
rect 11333 3615 11391 3621
rect 32324 3624 34376 3652
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2372 3556 2881 3584
rect 2372 3544 2378 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3584 12587 3587
rect 14734 3584 14740 3596
rect 12575 3556 14740 3584
rect 12575 3553 12587 3556
rect 12529 3547 12587 3553
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 30650 3584 30656 3596
rect 30611 3556 30656 3584
rect 30650 3544 30656 3556
rect 30708 3544 30714 3596
rect 32324 3593 32352 3624
rect 34348 3596 34376 3624
rect 32309 3587 32367 3593
rect 32309 3553 32321 3587
rect 32355 3553 32367 3587
rect 32309 3547 32367 3553
rect 32861 3587 32919 3593
rect 32861 3553 32873 3587
rect 32907 3584 32919 3587
rect 33410 3584 33416 3596
rect 32907 3556 33416 3584
rect 32907 3553 32919 3556
rect 32861 3547 32919 3553
rect 33410 3544 33416 3556
rect 33468 3544 33474 3596
rect 33781 3587 33839 3593
rect 33781 3553 33793 3587
rect 33827 3584 33839 3587
rect 33962 3584 33968 3596
rect 33827 3556 33968 3584
rect 33827 3553 33839 3556
rect 33781 3547 33839 3553
rect 33962 3544 33968 3556
rect 34020 3544 34026 3596
rect 34330 3544 34336 3596
rect 34388 3584 34394 3596
rect 34793 3587 34851 3593
rect 34793 3584 34805 3587
rect 34388 3556 34805 3584
rect 34388 3544 34394 3556
rect 34793 3553 34805 3556
rect 34839 3584 34851 3587
rect 34882 3584 34888 3596
rect 34839 3556 34888 3584
rect 34839 3553 34851 3556
rect 34793 3547 34851 3553
rect 34882 3544 34888 3556
rect 34940 3544 34946 3596
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 35805 3587 35863 3593
rect 35805 3584 35817 3587
rect 35492 3556 35817 3584
rect 35492 3544 35498 3556
rect 35805 3553 35817 3556
rect 35851 3553 35863 3587
rect 35805 3547 35863 3553
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 36725 3587 36783 3593
rect 36725 3584 36737 3587
rect 36136 3556 36737 3584
rect 36136 3544 36142 3556
rect 36725 3553 36737 3556
rect 36771 3553 36783 3587
rect 36725 3547 36783 3553
rect 37461 3587 37519 3593
rect 37461 3553 37473 3587
rect 37507 3584 37519 3587
rect 37734 3584 37740 3596
rect 37507 3556 37740 3584
rect 37507 3553 37519 3556
rect 37461 3547 37519 3553
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11517 3519 11575 3525
rect 11517 3516 11529 3519
rect 11112 3488 11529 3516
rect 11112 3476 11118 3488
rect 11517 3485 11529 3488
rect 11563 3485 11575 3519
rect 36740 3516 36768 3547
rect 37734 3544 37740 3556
rect 37792 3544 37798 3596
rect 38381 3587 38439 3593
rect 38381 3553 38393 3587
rect 38427 3584 38439 3587
rect 38654 3584 38660 3596
rect 38427 3556 38660 3584
rect 38427 3553 38439 3556
rect 38381 3547 38439 3553
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 39298 3584 39304 3596
rect 39259 3556 39304 3584
rect 39298 3544 39304 3556
rect 39356 3544 39362 3596
rect 41046 3584 41052 3596
rect 41007 3556 41052 3584
rect 41046 3544 41052 3556
rect 41104 3544 41110 3596
rect 42426 3584 42432 3596
rect 42387 3556 42432 3584
rect 42426 3544 42432 3556
rect 42484 3544 42490 3596
rect 42981 3587 43039 3593
rect 42981 3553 42993 3587
rect 43027 3584 43039 3587
rect 43070 3584 43076 3596
rect 43027 3556 43076 3584
rect 43027 3553 43039 3556
rect 42981 3547 43039 3553
rect 43070 3544 43076 3556
rect 43128 3544 43134 3596
rect 43717 3587 43775 3593
rect 43717 3553 43729 3587
rect 43763 3553 43775 3587
rect 43916 3584 43944 3680
rect 55582 3652 55588 3664
rect 55543 3624 55588 3652
rect 55582 3612 55588 3624
rect 55640 3612 55646 3664
rect 55674 3612 55680 3664
rect 55732 3652 55738 3664
rect 55732 3624 56916 3652
rect 55732 3612 55738 3624
rect 44729 3587 44787 3593
rect 44729 3584 44741 3587
rect 43916 3556 44741 3584
rect 43717 3547 43775 3553
rect 44729 3553 44741 3556
rect 44775 3553 44787 3587
rect 44729 3547 44787 3553
rect 46385 3587 46443 3593
rect 46385 3553 46397 3587
rect 46431 3584 46443 3587
rect 47029 3587 47087 3593
rect 47029 3584 47041 3587
rect 46431 3556 47041 3584
rect 46431 3553 46443 3556
rect 46385 3547 46443 3553
rect 47029 3553 47041 3556
rect 47075 3584 47087 3587
rect 47210 3584 47216 3596
rect 47075 3556 47216 3584
rect 47075 3553 47087 3556
rect 47029 3547 47087 3553
rect 43732 3516 43760 3547
rect 47210 3544 47216 3556
rect 47268 3544 47274 3596
rect 47578 3584 47584 3596
rect 47539 3556 47584 3584
rect 47578 3544 47584 3556
rect 47636 3544 47642 3596
rect 48498 3584 48504 3596
rect 48459 3556 48504 3584
rect 48498 3544 48504 3556
rect 48556 3544 48562 3596
rect 49789 3587 49847 3593
rect 49789 3553 49801 3587
rect 49835 3584 49847 3587
rect 49878 3584 49884 3596
rect 49835 3556 49884 3584
rect 49835 3553 49847 3556
rect 49789 3547 49847 3553
rect 49878 3544 49884 3556
rect 49936 3544 49942 3596
rect 50154 3544 50160 3596
rect 50212 3584 50218 3596
rect 50341 3587 50399 3593
rect 50341 3584 50353 3587
rect 50212 3556 50353 3584
rect 50212 3544 50218 3556
rect 50341 3553 50353 3556
rect 50387 3553 50399 3587
rect 50341 3547 50399 3553
rect 51442 3544 51448 3596
rect 51500 3584 51506 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 51500 3556 51549 3584
rect 51500 3544 51506 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 52273 3587 52331 3593
rect 52273 3553 52285 3587
rect 52319 3584 52331 3587
rect 52638 3584 52644 3596
rect 52319 3556 52644 3584
rect 52319 3553 52331 3556
rect 52273 3547 52331 3553
rect 52638 3544 52644 3556
rect 52696 3544 52702 3596
rect 53098 3584 53104 3596
rect 53059 3556 53104 3584
rect 53098 3544 53104 3556
rect 53156 3544 53162 3596
rect 53282 3584 53288 3596
rect 53243 3556 53288 3584
rect 53282 3544 53288 3556
rect 53340 3544 53346 3596
rect 54294 3584 54300 3596
rect 54255 3556 54300 3584
rect 54294 3544 54300 3556
rect 54352 3544 54358 3596
rect 55306 3544 55312 3596
rect 55364 3584 55370 3596
rect 56778 3584 56784 3596
rect 55364 3556 56784 3584
rect 55364 3544 55370 3556
rect 56778 3544 56784 3556
rect 56836 3544 56842 3596
rect 56888 3593 56916 3624
rect 56873 3587 56931 3593
rect 56873 3553 56885 3587
rect 56919 3553 56931 3587
rect 56873 3547 56931 3553
rect 56962 3544 56968 3596
rect 57020 3584 57026 3596
rect 57517 3587 57575 3593
rect 57517 3584 57529 3587
rect 57020 3556 57529 3584
rect 57020 3544 57026 3556
rect 57517 3553 57529 3556
rect 57563 3553 57575 3587
rect 57517 3547 57575 3553
rect 47670 3516 47676 3528
rect 36740 3488 47676 3516
rect 11517 3479 11575 3485
rect 47670 3476 47676 3488
rect 47728 3476 47734 3528
rect 57333 3519 57391 3525
rect 57333 3485 57345 3519
rect 57379 3516 57391 3519
rect 57422 3516 57428 3528
rect 57379 3488 57428 3516
rect 57379 3485 57391 3488
rect 57333 3479 57391 3485
rect 57422 3476 57428 3488
rect 57480 3476 57486 3528
rect 46201 3451 46259 3457
rect 46201 3417 46213 3451
rect 46247 3448 46259 3451
rect 47210 3448 47216 3460
rect 46247 3420 47216 3448
rect 46247 3417 46259 3420
rect 46201 3411 46259 3417
rect 47210 3408 47216 3420
rect 47268 3408 47274 3460
rect 55769 3451 55827 3457
rect 55769 3417 55781 3451
rect 55815 3448 55827 3451
rect 55950 3448 55956 3460
rect 55815 3420 55956 3448
rect 55815 3417 55827 3420
rect 55769 3411 55827 3417
rect 55950 3408 55956 3420
rect 56008 3408 56014 3460
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 8294 3380 8300 3392
rect 2096 3352 8300 3380
rect 2096 3340 2102 3352
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 29457 3383 29515 3389
rect 29457 3380 29469 3383
rect 29144 3352 29469 3380
rect 29144 3340 29150 3352
rect 29457 3349 29469 3352
rect 29503 3349 29515 3383
rect 29457 3343 29515 3349
rect 30190 3340 30196 3392
rect 30248 3380 30254 3392
rect 30469 3383 30527 3389
rect 30469 3380 30481 3383
rect 30248 3352 30481 3380
rect 30248 3340 30254 3352
rect 30469 3349 30481 3352
rect 30515 3349 30527 3383
rect 30469 3343 30527 3349
rect 30926 3340 30932 3392
rect 30984 3380 30990 3392
rect 31297 3383 31355 3389
rect 31297 3380 31309 3383
rect 30984 3352 31309 3380
rect 30984 3340 30990 3352
rect 31297 3349 31309 3352
rect 31343 3349 31355 3383
rect 32122 3380 32128 3392
rect 32083 3352 32128 3380
rect 31297 3343 31355 3349
rect 32122 3340 32128 3352
rect 32180 3340 32186 3392
rect 32766 3340 32772 3392
rect 32824 3380 32830 3392
rect 32953 3383 33011 3389
rect 32953 3380 32965 3383
rect 32824 3352 32965 3380
rect 32824 3340 32830 3352
rect 32953 3349 32965 3352
rect 32999 3349 33011 3383
rect 32953 3343 33011 3349
rect 33686 3340 33692 3392
rect 33744 3380 33750 3392
rect 33873 3383 33931 3389
rect 33873 3380 33885 3383
rect 33744 3352 33885 3380
rect 33744 3340 33750 3352
rect 33873 3349 33885 3352
rect 33919 3349 33931 3383
rect 34606 3380 34612 3392
rect 34567 3352 34612 3380
rect 33873 3343 33931 3349
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 35526 3340 35532 3392
rect 35584 3380 35590 3392
rect 35897 3383 35955 3389
rect 35897 3380 35909 3383
rect 35584 3352 35909 3380
rect 35584 3340 35590 3352
rect 35897 3349 35909 3352
rect 35943 3349 35955 3383
rect 35897 3343 35955 3349
rect 37366 3340 37372 3392
rect 37424 3380 37430 3392
rect 37553 3383 37611 3389
rect 37553 3380 37565 3383
rect 37424 3352 37565 3380
rect 37424 3340 37430 3352
rect 37553 3349 37565 3352
rect 37599 3349 37611 3383
rect 37553 3343 37611 3349
rect 38286 3340 38292 3392
rect 38344 3380 38350 3392
rect 38473 3383 38531 3389
rect 38473 3380 38485 3383
rect 38344 3352 38485 3380
rect 38344 3340 38350 3352
rect 38473 3349 38485 3352
rect 38519 3349 38531 3383
rect 38473 3343 38531 3349
rect 39206 3340 39212 3392
rect 39264 3380 39270 3392
rect 39393 3383 39451 3389
rect 39393 3380 39405 3383
rect 39264 3352 39405 3380
rect 39264 3340 39270 3352
rect 39393 3349 39405 3352
rect 39439 3349 39451 3383
rect 39393 3343 39451 3349
rect 40126 3340 40132 3392
rect 40184 3380 40190 3392
rect 41141 3383 41199 3389
rect 41141 3380 41153 3383
rect 40184 3352 41153 3380
rect 40184 3340 40190 3352
rect 41141 3349 41153 3352
rect 41187 3349 41199 3383
rect 41141 3343 41199 3349
rect 42245 3383 42303 3389
rect 42245 3349 42257 3383
rect 42291 3380 42303 3383
rect 42794 3380 42800 3392
rect 42291 3352 42800 3380
rect 42291 3349 42303 3352
rect 42245 3343 42303 3349
rect 42794 3340 42800 3352
rect 42852 3340 42858 3392
rect 42886 3340 42892 3392
rect 42944 3380 42950 3392
rect 43073 3383 43131 3389
rect 43073 3380 43085 3383
rect 42944 3352 43085 3380
rect 42944 3340 42950 3352
rect 43073 3349 43085 3352
rect 43119 3349 43131 3383
rect 43073 3343 43131 3349
rect 44545 3383 44603 3389
rect 44545 3349 44557 3383
rect 44591 3380 44603 3383
rect 45554 3380 45560 3392
rect 44591 3352 45560 3380
rect 44591 3349 44603 3352
rect 44545 3343 44603 3349
rect 45554 3340 45560 3352
rect 45612 3340 45618 3392
rect 46845 3383 46903 3389
rect 46845 3349 46857 3383
rect 46891 3380 46903 3383
rect 47394 3380 47400 3392
rect 46891 3352 47400 3380
rect 46891 3349 46903 3352
rect 46845 3343 46903 3349
rect 47394 3340 47400 3352
rect 47452 3340 47458 3392
rect 47486 3340 47492 3392
rect 47544 3380 47550 3392
rect 47673 3383 47731 3389
rect 47673 3380 47685 3383
rect 47544 3352 47685 3380
rect 47544 3340 47550 3352
rect 47673 3349 47685 3352
rect 47719 3349 47731 3383
rect 47673 3343 47731 3349
rect 48406 3340 48412 3392
rect 48464 3380 48470 3392
rect 48593 3383 48651 3389
rect 48593 3380 48605 3383
rect 48464 3352 48605 3380
rect 48464 3340 48470 3352
rect 48593 3349 48605 3352
rect 48639 3349 48651 3383
rect 49602 3380 49608 3392
rect 49563 3352 49608 3380
rect 48593 3343 48651 3349
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 50062 3340 50068 3392
rect 50120 3380 50126 3392
rect 50433 3383 50491 3389
rect 50433 3380 50445 3383
rect 50120 3352 50445 3380
rect 50120 3340 50126 3352
rect 50433 3349 50445 3352
rect 50479 3349 50491 3383
rect 50433 3343 50491 3349
rect 51166 3340 51172 3392
rect 51224 3380 51230 3392
rect 51629 3383 51687 3389
rect 51629 3380 51641 3383
rect 51224 3352 51641 3380
rect 51224 3340 51230 3352
rect 51629 3349 51641 3352
rect 51675 3349 51687 3383
rect 51629 3343 51687 3349
rect 52086 3340 52092 3392
rect 52144 3380 52150 3392
rect 52365 3383 52423 3389
rect 52365 3380 52377 3383
rect 52144 3352 52377 3380
rect 52144 3340 52150 3352
rect 52365 3349 52377 3352
rect 52411 3349 52423 3383
rect 52365 3343 52423 3349
rect 53006 3340 53012 3392
rect 53064 3380 53070 3392
rect 54389 3383 54447 3389
rect 54389 3380 54401 3383
rect 53064 3352 54401 3380
rect 53064 3340 53070 3352
rect 54389 3349 54401 3352
rect 54435 3349 54447 3383
rect 57974 3380 57980 3392
rect 57935 3352 57980 3380
rect 54389 3343 54447 3349
rect 57974 3340 57980 3352
rect 58032 3340 58038 3392
rect 1104 3290 58880 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 58880 3290
rect 1104 3216 58880 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1670 3176 1676 3188
rect 1627 3148 1676 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1670 3136 1676 3148
rect 1728 3176 1734 3188
rect 2038 3176 2044 3188
rect 1728 3148 2044 3176
rect 1728 3136 1734 3148
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3050 3176 3056 3188
rect 3011 3148 3056 3176
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 33410 3176 33416 3188
rect 33371 3148 33416 3176
rect 33410 3136 33416 3148
rect 33468 3136 33474 3188
rect 35434 3176 35440 3188
rect 35395 3148 35440 3176
rect 35434 3136 35440 3148
rect 35492 3136 35498 3188
rect 38654 3176 38660 3188
rect 38615 3148 38660 3176
rect 38654 3136 38660 3148
rect 38712 3136 38718 3188
rect 39298 3136 39304 3188
rect 39356 3176 39362 3188
rect 39761 3179 39819 3185
rect 39761 3176 39773 3179
rect 39356 3148 39773 3176
rect 39356 3136 39362 3148
rect 39761 3145 39773 3148
rect 39807 3145 39819 3179
rect 47578 3176 47584 3188
rect 47539 3148 47584 3176
rect 39761 3139 39819 3145
rect 47578 3136 47584 3148
rect 47636 3136 47642 3188
rect 51442 3176 51448 3188
rect 51403 3148 51448 3176
rect 51442 3136 51448 3148
rect 51500 3136 51506 3188
rect 52825 3179 52883 3185
rect 52825 3145 52837 3179
rect 52871 3176 52883 3179
rect 54294 3176 54300 3188
rect 52871 3148 54300 3176
rect 52871 3145 52883 3148
rect 52825 3139 52883 3145
rect 54294 3136 54300 3148
rect 54352 3136 54358 3188
rect 54662 3176 54668 3188
rect 54623 3148 54668 3176
rect 54662 3136 54668 3148
rect 54720 3136 54726 3188
rect 55769 3179 55827 3185
rect 55769 3145 55781 3179
rect 55815 3176 55827 3179
rect 55858 3176 55864 3188
rect 55815 3148 55864 3176
rect 55815 3145 55827 3148
rect 55769 3139 55827 3145
rect 55858 3136 55864 3148
rect 55916 3136 55922 3188
rect 56410 3136 56416 3188
rect 56468 3176 56474 3188
rect 56689 3179 56747 3185
rect 56689 3176 56701 3179
rect 56468 3148 56701 3176
rect 56468 3136 56474 3148
rect 56689 3145 56701 3148
rect 56735 3145 56747 3179
rect 56689 3139 56747 3145
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 30650 3108 30656 3120
rect 4764 3080 30656 3108
rect 4764 3068 4770 3080
rect 30650 3068 30656 3080
rect 30708 3068 30714 3120
rect 49602 3068 49608 3120
rect 49660 3108 49666 3120
rect 49660 3080 51028 3108
rect 49660 3068 49666 3080
rect 8938 3040 8944 3052
rect 2240 3012 8944 3040
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 2240 2981 2268 3012
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 30006 3040 30012 3052
rect 29967 3012 30012 3040
rect 30006 3000 30012 3012
rect 30064 3000 30070 3052
rect 30190 3040 30196 3052
rect 30151 3012 30196 3040
rect 30190 3000 30196 3012
rect 30248 3000 30254 3052
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 532 2944 1409 2972
rect 532 2932 538 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2941 2283 2975
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 2225 2935 2283 2941
rect 2884 2944 3617 2972
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 2774 2904 2780 2916
rect 2455 2876 2780 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 2884 2836 2912 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 4249 2975 4307 2981
rect 4249 2941 4261 2975
rect 4295 2941 4307 2975
rect 28074 2972 28080 2984
rect 28035 2944 28080 2972
rect 4249 2935 4307 2941
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2873 3019 2907
rect 2961 2867 3019 2873
rect 1452 2808 2912 2836
rect 2976 2836 3004 2867
rect 3234 2864 3240 2916
rect 3292 2904 3298 2916
rect 4264 2904 4292 2935
rect 28074 2932 28080 2944
rect 28132 2932 28138 2984
rect 28721 2975 28779 2981
rect 28721 2941 28733 2975
rect 28767 2972 28779 2975
rect 28994 2972 29000 2984
rect 28767 2944 29000 2972
rect 28767 2941 28779 2944
rect 28721 2935 28779 2941
rect 28994 2932 29000 2944
rect 29052 2932 29058 2984
rect 29546 2972 29552 2984
rect 29507 2944 29552 2972
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 30668 2972 30696 3068
rect 32122 3000 32128 3052
rect 32180 3040 32186 3052
rect 33229 3043 33287 3049
rect 33229 3040 33241 3043
rect 32180 3012 33241 3040
rect 32180 3000 32186 3012
rect 33229 3009 33241 3012
rect 33275 3009 33287 3043
rect 33229 3003 33287 3009
rect 34606 3000 34612 3052
rect 34664 3040 34670 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34664 3012 34989 3040
rect 34664 3000 34670 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 34977 3003 35035 3009
rect 38289 3043 38347 3049
rect 38289 3009 38301 3043
rect 38335 3040 38347 3043
rect 38562 3040 38568 3052
rect 38335 3012 38568 3040
rect 38335 3009 38347 3012
rect 38289 3003 38347 3009
rect 38562 3000 38568 3012
rect 38620 3000 38626 3052
rect 39390 3040 39396 3052
rect 39351 3012 39396 3040
rect 39390 3000 39396 3012
rect 39448 3000 39454 3052
rect 39574 3040 39580 3052
rect 39535 3012 39580 3040
rect 39574 3000 39580 3012
rect 39632 3000 39638 3052
rect 39758 3000 39764 3052
rect 39816 3040 39822 3052
rect 40681 3043 40739 3049
rect 40681 3040 40693 3043
rect 39816 3012 40693 3040
rect 39816 3000 39822 3012
rect 40681 3009 40693 3012
rect 40727 3009 40739 3043
rect 40681 3003 40739 3009
rect 43438 3000 43444 3052
rect 43496 3040 43502 3052
rect 43533 3043 43591 3049
rect 43533 3040 43545 3043
rect 43496 3012 43545 3040
rect 43496 3000 43502 3012
rect 43533 3009 43545 3012
rect 43579 3009 43591 3043
rect 43714 3040 43720 3052
rect 43675 3012 43720 3040
rect 43533 3003 43591 3009
rect 43714 3000 43720 3012
rect 43772 3000 43778 3052
rect 44726 3000 44732 3052
rect 44784 3040 44790 3052
rect 45649 3043 45707 3049
rect 45649 3040 45661 3043
rect 44784 3012 45661 3040
rect 44784 3000 44790 3012
rect 45649 3009 45661 3012
rect 45695 3009 45707 3043
rect 47118 3040 47124 3052
rect 47079 3012 47124 3040
rect 45649 3003 45707 3009
rect 47118 3000 47124 3012
rect 47176 3000 47182 3052
rect 48958 3040 48964 3052
rect 48919 3012 48964 3040
rect 48958 3000 48964 3012
rect 49016 3000 49022 3052
rect 50614 3000 50620 3052
rect 50672 3040 50678 3052
rect 51000 3049 51028 3080
rect 51994 3068 52000 3120
rect 52052 3108 52058 3120
rect 52052 3080 54248 3108
rect 52052 3068 52058 3080
rect 50801 3043 50859 3049
rect 50801 3040 50813 3043
rect 50672 3012 50813 3040
rect 50672 3000 50678 3012
rect 50801 3009 50813 3012
rect 50847 3009 50859 3043
rect 50801 3003 50859 3009
rect 50985 3043 51043 3049
rect 50985 3009 50997 3043
rect 51031 3009 51043 3043
rect 50985 3003 51043 3009
rect 52181 3043 52239 3049
rect 52181 3009 52193 3043
rect 52227 3040 52239 3043
rect 52454 3040 52460 3052
rect 52227 3012 52460 3040
rect 52227 3009 52239 3012
rect 52181 3003 52239 3009
rect 52454 3000 52460 3012
rect 52512 3000 52518 3052
rect 54018 3040 54024 3052
rect 53979 3012 54024 3040
rect 54018 3000 54024 3012
rect 54076 3000 54082 3052
rect 54220 3049 54248 3080
rect 54754 3068 54760 3120
rect 54812 3108 54818 3120
rect 54812 3080 56456 3108
rect 54812 3068 54818 3080
rect 54205 3043 54263 3049
rect 54205 3009 54217 3043
rect 54251 3009 54263 3043
rect 54205 3003 54263 3009
rect 54478 3000 54484 3052
rect 54536 3040 54542 3052
rect 55125 3043 55183 3049
rect 55125 3040 55137 3043
rect 54536 3012 55137 3040
rect 54536 3000 54542 3012
rect 55125 3009 55137 3012
rect 55171 3009 55183 3043
rect 55125 3003 55183 3009
rect 55398 3000 55404 3052
rect 55456 3040 55462 3052
rect 56428 3049 56456 3080
rect 56594 3068 56600 3120
rect 56652 3108 56658 3120
rect 57885 3111 57943 3117
rect 57885 3108 57897 3111
rect 56652 3080 57897 3108
rect 56652 3068 56658 3080
rect 57885 3077 57897 3080
rect 57931 3077 57943 3111
rect 57885 3071 57943 3077
rect 56229 3043 56287 3049
rect 56229 3040 56241 3043
rect 55456 3012 56241 3040
rect 55456 3000 55462 3012
rect 56229 3009 56241 3012
rect 56275 3009 56287 3043
rect 56229 3003 56287 3009
rect 56413 3043 56471 3049
rect 56413 3009 56425 3043
rect 56459 3009 56471 3043
rect 56413 3003 56471 3009
rect 57238 3000 57244 3052
rect 57296 3040 57302 3052
rect 57701 3043 57759 3049
rect 57701 3040 57713 3043
rect 57296 3012 57713 3040
rect 57296 3000 57302 3012
rect 57701 3009 57713 3012
rect 57747 3009 57759 3043
rect 57701 3003 57759 3009
rect 31297 2975 31355 2981
rect 31297 2972 31309 2975
rect 30668 2944 31309 2972
rect 31297 2941 31309 2944
rect 31343 2941 31355 2975
rect 33042 2972 33048 2984
rect 33003 2944 33048 2972
rect 31297 2935 31355 2941
rect 33042 2932 33048 2944
rect 33100 2932 33106 2984
rect 34330 2972 34336 2984
rect 34291 2944 34336 2972
rect 34330 2932 34336 2944
rect 34388 2932 34394 2984
rect 34793 2975 34851 2981
rect 34793 2941 34805 2975
rect 34839 2972 34851 2975
rect 35250 2972 35256 2984
rect 34839 2944 35256 2972
rect 34839 2941 34851 2944
rect 34793 2935 34851 2941
rect 35250 2932 35256 2944
rect 35308 2932 35314 2984
rect 36173 2975 36231 2981
rect 36173 2972 36185 2975
rect 35866 2944 36185 2972
rect 3292 2876 4292 2904
rect 30653 2907 30711 2913
rect 3292 2864 3298 2876
rect 30653 2873 30665 2907
rect 30699 2904 30711 2907
rect 31754 2904 31760 2916
rect 30699 2876 31760 2904
rect 30699 2873 30711 2876
rect 30653 2867 30711 2873
rect 31754 2864 31760 2876
rect 31812 2864 31818 2916
rect 31938 2904 31944 2916
rect 31899 2876 31944 2904
rect 31938 2864 31944 2876
rect 31996 2864 32002 2916
rect 34606 2864 34612 2916
rect 34664 2904 34670 2916
rect 35866 2904 35894 2944
rect 36173 2941 36185 2944
rect 36219 2941 36231 2975
rect 36173 2935 36231 2941
rect 38378 2932 38384 2984
rect 38436 2972 38442 2984
rect 38473 2975 38531 2981
rect 38473 2972 38485 2975
rect 38436 2944 38485 2972
rect 38436 2932 38442 2944
rect 38473 2941 38485 2944
rect 38519 2941 38531 2975
rect 38473 2935 38531 2941
rect 40497 2975 40555 2981
rect 40497 2941 40509 2975
rect 40543 2972 40555 2975
rect 41230 2972 41236 2984
rect 40543 2944 41236 2972
rect 40543 2941 40555 2944
rect 40497 2935 40555 2941
rect 41230 2932 41236 2944
rect 41288 2932 41294 2984
rect 46937 2975 46995 2981
rect 46937 2941 46949 2975
rect 46983 2972 46995 2975
rect 47026 2972 47032 2984
rect 46983 2944 47032 2972
rect 46983 2941 46995 2944
rect 46937 2935 46995 2941
rect 47026 2932 47032 2944
rect 47084 2932 47090 2984
rect 48777 2975 48835 2981
rect 48777 2941 48789 2975
rect 48823 2972 48835 2975
rect 49050 2972 49056 2984
rect 48823 2944 49056 2972
rect 48823 2941 48835 2944
rect 48777 2935 48835 2941
rect 49050 2932 49056 2944
rect 49108 2932 49114 2984
rect 51718 2932 51724 2984
rect 51776 2972 51782 2984
rect 52365 2975 52423 2981
rect 52365 2972 52377 2975
rect 51776 2944 52377 2972
rect 51776 2932 51782 2944
rect 52365 2941 52377 2944
rect 52411 2941 52423 2975
rect 52365 2935 52423 2941
rect 53742 2932 53748 2984
rect 53800 2972 53806 2984
rect 55309 2975 55367 2981
rect 55309 2972 55321 2975
rect 53800 2944 55321 2972
rect 53800 2932 53806 2944
rect 55309 2941 55321 2944
rect 55355 2941 55367 2975
rect 55309 2935 55367 2941
rect 57146 2932 57152 2984
rect 57204 2972 57210 2984
rect 57517 2975 57575 2981
rect 57517 2972 57529 2975
rect 57204 2944 57529 2972
rect 57204 2932 57210 2944
rect 57517 2941 57529 2944
rect 57563 2941 57575 2975
rect 57517 2935 57575 2941
rect 35986 2904 35992 2916
rect 34664 2876 35894 2904
rect 35947 2876 35992 2904
rect 34664 2864 34670 2876
rect 35986 2864 35992 2876
rect 36044 2864 36050 2916
rect 36722 2904 36728 2916
rect 36683 2876 36728 2904
rect 36722 2864 36728 2876
rect 36780 2864 36786 2916
rect 41141 2907 41199 2913
rect 41141 2873 41153 2907
rect 41187 2904 41199 2907
rect 41693 2907 41751 2913
rect 41693 2904 41705 2907
rect 41187 2876 41705 2904
rect 41187 2873 41199 2876
rect 41141 2867 41199 2873
rect 41693 2873 41705 2876
rect 41739 2873 41751 2907
rect 42426 2904 42432 2916
rect 42387 2876 42432 2904
rect 41693 2867 41751 2873
rect 42426 2864 42432 2876
rect 42484 2864 42490 2916
rect 44177 2907 44235 2913
rect 44177 2873 44189 2907
rect 44223 2904 44235 2907
rect 44729 2907 44787 2913
rect 44729 2904 44741 2907
rect 44223 2876 44741 2904
rect 44223 2873 44235 2876
rect 44177 2867 44235 2873
rect 44729 2873 44741 2876
rect 44775 2873 44787 2907
rect 45462 2904 45468 2916
rect 45423 2876 45468 2904
rect 44729 2867 44787 2873
rect 45462 2864 45468 2876
rect 45520 2864 45526 2916
rect 46198 2904 46204 2916
rect 46159 2876 46204 2904
rect 46198 2864 46204 2876
rect 46256 2864 46262 2916
rect 49421 2907 49479 2913
rect 49421 2873 49433 2907
rect 49467 2904 49479 2907
rect 49973 2907 50031 2913
rect 49973 2904 49985 2907
rect 49467 2876 49985 2904
rect 49467 2873 49479 2876
rect 49421 2867 49479 2873
rect 49973 2873 49985 2876
rect 50019 2873 50031 2907
rect 49973 2867 50031 2873
rect 55214 2864 55220 2916
rect 55272 2904 55278 2916
rect 59446 2904 59452 2916
rect 55272 2876 59452 2904
rect 55272 2864 55278 2876
rect 59446 2864 59452 2876
rect 59504 2864 59510 2916
rect 6454 2836 6460 2848
rect 2976 2808 6460 2836
rect 1452 2796 1458 2808
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 29362 2836 29368 2848
rect 29323 2808 29368 2836
rect 29362 2796 29368 2808
rect 29420 2796 29426 2848
rect 31110 2836 31116 2848
rect 31071 2808 31116 2836
rect 31110 2796 31116 2808
rect 31168 2796 31174 2848
rect 31846 2796 31852 2848
rect 31904 2836 31910 2848
rect 32033 2839 32091 2845
rect 32033 2836 32045 2839
rect 31904 2808 32045 2836
rect 31904 2796 31910 2808
rect 32033 2805 32045 2808
rect 32079 2805 32091 2839
rect 32033 2799 32091 2805
rect 34149 2839 34207 2845
rect 34149 2805 34161 2839
rect 34195 2836 34207 2839
rect 34974 2836 34980 2848
rect 34195 2808 34980 2836
rect 34195 2805 34207 2808
rect 34149 2799 34207 2805
rect 34974 2796 34980 2808
rect 35032 2796 35038 2848
rect 36446 2796 36452 2848
rect 36504 2836 36510 2848
rect 36817 2839 36875 2845
rect 36817 2836 36829 2839
rect 36504 2808 36829 2836
rect 36504 2796 36510 2808
rect 36817 2805 36829 2808
rect 36863 2805 36875 2839
rect 36817 2799 36875 2805
rect 40954 2796 40960 2848
rect 41012 2836 41018 2848
rect 41785 2839 41843 2845
rect 41785 2836 41797 2839
rect 41012 2808 41797 2836
rect 41012 2796 41018 2808
rect 41785 2805 41797 2808
rect 41831 2805 41843 2839
rect 41785 2799 41843 2805
rect 41966 2796 41972 2848
rect 42024 2836 42030 2848
rect 42521 2839 42579 2845
rect 42521 2836 42533 2839
rect 42024 2808 42533 2836
rect 42024 2796 42030 2808
rect 42521 2805 42533 2808
rect 42567 2805 42579 2839
rect 42521 2799 42579 2805
rect 43806 2796 43812 2848
rect 43864 2836 43870 2848
rect 44821 2839 44879 2845
rect 44821 2836 44833 2839
rect 43864 2808 44833 2836
rect 43864 2796 43870 2808
rect 44821 2805 44833 2808
rect 44867 2805 44879 2839
rect 44821 2799 44879 2805
rect 45646 2796 45652 2848
rect 45704 2836 45710 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45704 2808 46305 2836
rect 45704 2796 45710 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50065 2839 50123 2845
rect 50065 2836 50077 2839
rect 49384 2808 50077 2836
rect 49384 2796 49390 2808
rect 50065 2805 50077 2808
rect 50111 2805 50123 2839
rect 50065 2799 50123 2805
rect 1104 2746 58880 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 50326 2746
rect 50378 2694 50390 2746
rect 50442 2694 50454 2746
rect 50506 2694 50518 2746
rect 50570 2694 58880 2746
rect 1104 2672 58880 2694
rect 31573 2635 31631 2641
rect 31573 2601 31585 2635
rect 31619 2632 31631 2635
rect 31938 2632 31944 2644
rect 31619 2604 31944 2632
rect 31619 2601 31631 2604
rect 31573 2595 31631 2601
rect 31938 2592 31944 2604
rect 31996 2592 32002 2644
rect 35345 2635 35403 2641
rect 35345 2601 35357 2635
rect 35391 2632 35403 2635
rect 35986 2632 35992 2644
rect 35391 2604 35992 2632
rect 35391 2601 35403 2604
rect 35345 2595 35403 2601
rect 35986 2592 35992 2604
rect 36044 2592 36050 2644
rect 36722 2592 36728 2644
rect 36780 2632 36786 2644
rect 36909 2635 36967 2641
rect 36909 2632 36921 2635
rect 36780 2604 36921 2632
rect 36780 2592 36786 2604
rect 36909 2601 36921 2604
rect 36955 2601 36967 2635
rect 36909 2595 36967 2601
rect 40129 2635 40187 2641
rect 40129 2601 40141 2635
rect 40175 2632 40187 2635
rect 41046 2632 41052 2644
rect 40175 2604 41052 2632
rect 40175 2601 40187 2604
rect 40129 2595 40187 2601
rect 41046 2592 41052 2604
rect 41104 2592 41110 2644
rect 42245 2635 42303 2641
rect 42245 2601 42257 2635
rect 42291 2632 42303 2635
rect 42426 2632 42432 2644
rect 42291 2604 42432 2632
rect 42291 2601 42303 2604
rect 42245 2595 42303 2601
rect 42426 2592 42432 2604
rect 42484 2592 42490 2644
rect 44913 2635 44971 2641
rect 44913 2601 44925 2635
rect 44959 2632 44971 2635
rect 45462 2632 45468 2644
rect 44959 2604 45468 2632
rect 44959 2601 44971 2604
rect 44913 2595 44971 2601
rect 45462 2592 45468 2604
rect 45520 2592 45526 2644
rect 46017 2635 46075 2641
rect 46017 2601 46029 2635
rect 46063 2632 46075 2635
rect 46198 2632 46204 2644
rect 46063 2604 46204 2632
rect 46063 2601 46075 2604
rect 46017 2595 46075 2601
rect 46198 2592 46204 2604
rect 46256 2592 46262 2644
rect 48498 2592 48504 2644
rect 48556 2632 48562 2644
rect 48685 2635 48743 2641
rect 48685 2632 48697 2635
rect 48556 2604 48697 2632
rect 48556 2592 48562 2604
rect 48685 2601 48697 2604
rect 48731 2601 48743 2635
rect 48685 2595 48743 2601
rect 50154 2592 50160 2644
rect 50212 2632 50218 2644
rect 50249 2635 50307 2641
rect 50249 2632 50261 2635
rect 50212 2604 50261 2632
rect 50212 2592 50218 2604
rect 50249 2601 50261 2604
rect 50295 2601 50307 2635
rect 56686 2632 56692 2644
rect 56647 2604 56692 2632
rect 50249 2595 50307 2601
rect 56686 2592 56692 2604
rect 56744 2592 56750 2644
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 11054 2564 11060 2576
rect 2823 2536 11060 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 11054 2524 11060 2536
rect 11112 2524 11118 2576
rect 28445 2567 28503 2573
rect 28445 2533 28457 2567
rect 28491 2564 28503 2567
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 28491 2536 29745 2564
rect 28491 2533 28503 2536
rect 28445 2527 28503 2533
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 31754 2524 31760 2576
rect 31812 2564 31818 2576
rect 32125 2567 32183 2573
rect 32125 2564 32137 2567
rect 31812 2536 32137 2564
rect 31812 2524 31818 2536
rect 32125 2533 32137 2536
rect 32171 2533 32183 2567
rect 32125 2527 32183 2533
rect 47581 2567 47639 2573
rect 47581 2533 47593 2567
rect 47627 2564 47639 2567
rect 50801 2567 50859 2573
rect 50801 2564 50813 2567
rect 47627 2536 50813 2564
rect 47627 2533 47639 2536
rect 47581 2527 47639 2533
rect 50801 2533 50813 2536
rect 50847 2533 50859 2567
rect 53834 2564 53840 2576
rect 53795 2536 53840 2564
rect 50801 2527 50859 2533
rect 53834 2524 53840 2536
rect 53892 2524 53898 2576
rect 54021 2567 54079 2573
rect 54021 2533 54033 2567
rect 54067 2564 54079 2567
rect 55214 2564 55220 2576
rect 54067 2536 55220 2564
rect 54067 2533 54079 2536
rect 54021 2527 54079 2533
rect 55214 2524 55220 2536
rect 55272 2524 55278 2576
rect 55401 2567 55459 2573
rect 55401 2533 55413 2567
rect 55447 2564 55459 2567
rect 56594 2564 56600 2576
rect 55447 2536 56600 2564
rect 55447 2533 55459 2536
rect 55401 2527 55459 2533
rect 56594 2524 56600 2536
rect 56652 2524 56658 2576
rect 57974 2564 57980 2576
rect 57935 2536 57980 2564
rect 57974 2524 57980 2536
rect 58032 2524 58038 2576
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4249 2499 4307 2505
rect 4249 2496 4261 2499
rect 4212 2468 4261 2496
rect 4212 2456 4218 2468
rect 4249 2465 4261 2468
rect 4295 2465 4307 2499
rect 5074 2496 5080 2508
rect 5035 2468 5080 2496
rect 4249 2459 4307 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 5994 2496 6000 2508
rect 5859 2468 6000 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 7834 2496 7840 2508
rect 6972 2468 7017 2496
rect 7795 2468 7840 2496
rect 6972 2456 6978 2468
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 8754 2496 8760 2508
rect 8527 2468 8760 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9674 2496 9680 2508
rect 9635 2468 9680 2496
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10594 2496 10600 2508
rect 10555 2468 10600 2496
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 12253 2499 12311 2505
rect 12253 2496 12265 2499
rect 11572 2468 12265 2496
rect 11572 2456 11578 2468
rect 12253 2465 12265 2468
rect 12299 2465 12311 2499
rect 12253 2459 12311 2465
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12492 2468 12909 2496
rect 12492 2456 12498 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 13541 2499 13599 2505
rect 13541 2496 13553 2499
rect 13412 2468 13553 2496
rect 13412 2456 13418 2468
rect 13541 2465 13553 2468
rect 13587 2465 13599 2499
rect 13541 2459 13599 2465
rect 14274 2456 14280 2508
rect 14332 2496 14338 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14332 2468 14933 2496
rect 14332 2456 14338 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15252 2468 15577 2496
rect 15252 2456 15258 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 16172 2468 16221 2496
rect 16172 2456 16178 2468
rect 16209 2465 16221 2468
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 17034 2456 17040 2508
rect 17092 2496 17098 2508
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 17092 2468 17601 2496
rect 17092 2456 17098 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18233 2499 18291 2505
rect 18233 2496 18245 2499
rect 18012 2468 18245 2496
rect 18012 2456 18018 2468
rect 18233 2465 18245 2468
rect 18279 2465 18291 2499
rect 18874 2496 18880 2508
rect 18835 2468 18880 2496
rect 18233 2459 18291 2465
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 19852 2468 20269 2496
rect 19852 2456 19858 2468
rect 20257 2465 20269 2468
rect 20303 2465 20315 2499
rect 20257 2459 20315 2465
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 20772 2468 20913 2496
rect 20772 2456 20778 2468
rect 20901 2465 20913 2468
rect 20947 2465 20959 2499
rect 21634 2496 21640 2508
rect 21595 2468 21640 2496
rect 20901 2459 20959 2465
rect 21634 2456 21640 2468
rect 21692 2456 21698 2508
rect 22554 2456 22560 2508
rect 22612 2496 22618 2508
rect 22925 2499 22983 2505
rect 22925 2496 22937 2499
rect 22612 2468 22937 2496
rect 22612 2456 22618 2468
rect 22925 2465 22937 2468
rect 22971 2465 22983 2499
rect 22925 2459 22983 2465
rect 23474 2456 23480 2508
rect 23532 2496 23538 2508
rect 23569 2499 23627 2505
rect 23569 2496 23581 2499
rect 23532 2468 23581 2496
rect 23532 2456 23538 2468
rect 23569 2465 23581 2468
rect 23615 2465 23627 2499
rect 24394 2496 24400 2508
rect 24355 2468 24400 2496
rect 23569 2459 23627 2465
rect 24394 2456 24400 2468
rect 24452 2456 24458 2508
rect 25314 2456 25320 2508
rect 25372 2496 25378 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 25372 2468 25605 2496
rect 25372 2456 25378 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 26234 2456 26240 2508
rect 26292 2496 26298 2508
rect 27154 2496 27160 2508
rect 26292 2468 26337 2496
rect 27115 2468 27160 2496
rect 26292 2456 26298 2468
rect 27154 2456 27160 2468
rect 27212 2456 27218 2508
rect 29086 2496 29092 2508
rect 29047 2468 29092 2496
rect 29086 2456 29092 2468
rect 29144 2456 29150 2508
rect 29273 2499 29331 2505
rect 29273 2465 29285 2499
rect 29319 2496 29331 2499
rect 29362 2496 29368 2508
rect 29319 2468 29368 2496
rect 29319 2465 29331 2468
rect 29273 2459 29331 2465
rect 29362 2456 29368 2468
rect 29420 2456 29426 2508
rect 30926 2496 30932 2508
rect 30887 2468 30932 2496
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 31110 2496 31116 2508
rect 31071 2468 31116 2496
rect 31110 2456 31116 2468
rect 31168 2456 31174 2508
rect 33594 2496 33600 2508
rect 33555 2468 33600 2496
rect 33594 2456 33600 2468
rect 33652 2456 33658 2508
rect 33778 2496 33784 2508
rect 33739 2468 33784 2496
rect 33778 2456 33784 2468
rect 33836 2456 33842 2508
rect 34701 2499 34759 2505
rect 34701 2465 34713 2499
rect 34747 2496 34759 2499
rect 34790 2496 34796 2508
rect 34747 2468 34796 2496
rect 34747 2465 34759 2468
rect 34701 2459 34759 2465
rect 34790 2456 34796 2468
rect 34848 2456 34854 2508
rect 34974 2456 34980 2508
rect 35032 2496 35038 2508
rect 36449 2499 36507 2505
rect 36449 2496 36461 2499
rect 35032 2468 36461 2496
rect 35032 2456 35038 2468
rect 36449 2465 36461 2468
rect 36495 2465 36507 2499
rect 36449 2459 36507 2465
rect 37274 2456 37280 2508
rect 37332 2496 37338 2508
rect 37369 2499 37427 2505
rect 37369 2496 37381 2499
rect 37332 2468 37381 2496
rect 37332 2456 37338 2468
rect 37369 2465 37381 2468
rect 37415 2465 37427 2499
rect 37550 2496 37556 2508
rect 37511 2468 37556 2496
rect 37369 2459 37427 2465
rect 37550 2456 37556 2468
rect 37608 2456 37614 2508
rect 39482 2496 39488 2508
rect 39443 2468 39488 2496
rect 39482 2456 39488 2468
rect 39540 2456 39546 2508
rect 39669 2499 39727 2505
rect 39669 2465 39681 2499
rect 39715 2496 39727 2499
rect 40402 2496 40408 2508
rect 39715 2468 40408 2496
rect 39715 2465 39727 2468
rect 39669 2459 39727 2465
rect 40402 2456 40408 2468
rect 40460 2456 40466 2508
rect 41506 2456 41512 2508
rect 41564 2496 41570 2508
rect 41601 2499 41659 2505
rect 41601 2496 41613 2499
rect 41564 2468 41613 2496
rect 41564 2456 41570 2468
rect 41601 2465 41613 2468
rect 41647 2465 41659 2499
rect 41601 2459 41659 2465
rect 41785 2499 41843 2505
rect 41785 2465 41797 2499
rect 41831 2496 41843 2499
rect 41874 2496 41880 2508
rect 41831 2468 41880 2496
rect 41831 2465 41843 2468
rect 41785 2459 41843 2465
rect 41874 2456 41880 2468
rect 41932 2456 41938 2508
rect 42334 2456 42340 2508
rect 42392 2496 42398 2508
rect 42705 2499 42763 2505
rect 42705 2496 42717 2499
rect 42392 2468 42717 2496
rect 42392 2456 42398 2468
rect 42705 2465 42717 2468
rect 42751 2465 42763 2499
rect 42705 2459 42763 2465
rect 42794 2456 42800 2508
rect 42852 2496 42858 2508
rect 42889 2499 42947 2505
rect 42889 2496 42901 2499
rect 42852 2468 42901 2496
rect 42852 2456 42858 2468
rect 42889 2465 42901 2468
rect 42935 2465 42947 2499
rect 44266 2496 44272 2508
rect 44227 2468 44272 2496
rect 42889 2459 42947 2465
rect 44266 2456 44272 2468
rect 44324 2456 44330 2508
rect 44450 2496 44456 2508
rect 44411 2468 44456 2496
rect 44450 2456 44456 2468
rect 44508 2456 44514 2508
rect 45373 2499 45431 2505
rect 45373 2465 45385 2499
rect 45419 2496 45431 2499
rect 45738 2496 45744 2508
rect 45419 2468 45744 2496
rect 45419 2465 45431 2468
rect 45373 2459 45431 2465
rect 45738 2456 45744 2468
rect 45796 2456 45802 2508
rect 46934 2496 46940 2508
rect 46895 2468 46940 2496
rect 46934 2456 46940 2468
rect 46992 2456 46998 2508
rect 47121 2499 47179 2505
rect 47121 2465 47133 2499
rect 47167 2496 47179 2499
rect 47210 2496 47216 2508
rect 47167 2468 47216 2496
rect 47167 2465 47179 2468
rect 47121 2459 47179 2465
rect 47210 2456 47216 2468
rect 47268 2456 47274 2508
rect 48038 2496 48044 2508
rect 47999 2468 48044 2496
rect 48038 2456 48044 2468
rect 48096 2456 48102 2508
rect 49786 2496 49792 2508
rect 49747 2468 49792 2496
rect 49786 2456 49792 2468
rect 49844 2456 49850 2508
rect 51626 2456 51632 2508
rect 51684 2496 51690 2508
rect 52273 2499 52331 2505
rect 52273 2496 52285 2499
rect 51684 2468 52285 2496
rect 51684 2456 51690 2468
rect 52273 2465 52285 2468
rect 52319 2465 52331 2499
rect 56042 2496 56048 2508
rect 56003 2468 56048 2496
rect 52273 2459 52331 2465
rect 56042 2456 56048 2468
rect 56100 2456 56106 2508
rect 34514 2388 34520 2440
rect 34572 2428 34578 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34572 2400 34897 2428
rect 34572 2388 34578 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36262 2428 36268 2440
rect 36223 2400 36268 2428
rect 34885 2391 34943 2397
rect 36262 2388 36268 2400
rect 36320 2388 36326 2440
rect 45554 2388 45560 2440
rect 45612 2428 45618 2440
rect 45612 2400 45657 2428
rect 45612 2388 45618 2400
rect 47394 2388 47400 2440
rect 47452 2428 47458 2440
rect 48225 2431 48283 2437
rect 48225 2428 48237 2431
rect 47452 2400 48237 2428
rect 47452 2388 47458 2400
rect 48225 2397 48237 2400
rect 48271 2397 48283 2431
rect 48225 2391 48283 2397
rect 49605 2431 49663 2437
rect 49605 2397 49617 2431
rect 49651 2428 49663 2431
rect 49694 2428 49700 2440
rect 49651 2400 49700 2428
rect 49651 2397 49663 2400
rect 49605 2391 49663 2397
rect 49694 2388 49700 2400
rect 49752 2388 49758 2440
rect 51534 2388 51540 2440
rect 51592 2428 51598 2440
rect 52457 2431 52515 2437
rect 52457 2428 52469 2431
rect 51592 2400 52469 2428
rect 51592 2388 51598 2400
rect 52457 2397 52469 2400
rect 52503 2397 52515 2431
rect 52457 2391 52515 2397
rect 52822 2388 52828 2440
rect 52880 2428 52886 2440
rect 56229 2431 56287 2437
rect 56229 2428 56241 2431
rect 52880 2400 56241 2428
rect 52880 2388 52886 2400
rect 56229 2397 56241 2400
rect 56275 2397 56287 2431
rect 56229 2391 56287 2397
rect 2225 2363 2283 2369
rect 2225 2329 2237 2363
rect 2271 2360 2283 2363
rect 28629 2363 28687 2369
rect 2271 2332 6914 2360
rect 2271 2329 2283 2332
rect 2225 2323 2283 2329
rect 2866 2292 2872 2304
rect 2827 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 6886 2292 6914 2332
rect 28629 2329 28641 2363
rect 28675 2360 28687 2363
rect 29914 2360 29920 2372
rect 28675 2332 29920 2360
rect 28675 2329 28687 2332
rect 28629 2323 28687 2329
rect 29914 2320 29920 2332
rect 29972 2320 29978 2372
rect 33962 2360 33968 2372
rect 33923 2332 33968 2360
rect 33962 2320 33968 2332
rect 34020 2320 34026 2372
rect 37734 2360 37740 2372
rect 37695 2332 37740 2360
rect 37734 2320 37740 2332
rect 37792 2320 37798 2372
rect 43070 2360 43076 2372
rect 43031 2332 43076 2360
rect 43070 2320 43076 2332
rect 43128 2320 43134 2372
rect 52638 2360 52644 2372
rect 52599 2332 52644 2360
rect 52638 2320 52644 2332
rect 52696 2320 52702 2372
rect 55582 2360 55588 2372
rect 55543 2332 55588 2360
rect 55582 2320 55588 2332
rect 55640 2320 55646 2372
rect 19426 2292 19432 2304
rect 6886 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 30926 2252 30932 2304
rect 30984 2292 30990 2304
rect 32217 2295 32275 2301
rect 32217 2292 32229 2295
rect 30984 2264 32229 2292
rect 30984 2252 30990 2264
rect 32217 2261 32229 2264
rect 32263 2261 32275 2295
rect 32217 2255 32275 2261
rect 46566 2252 46572 2304
rect 46624 2292 46630 2304
rect 50893 2295 50951 2301
rect 50893 2292 50905 2295
rect 46624 2264 50905 2292
rect 46624 2252 46630 2264
rect 50893 2261 50905 2264
rect 50939 2261 50951 2295
rect 50893 2255 50951 2261
rect 57882 2252 57888 2304
rect 57940 2292 57946 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 57940 2264 58081 2292
rect 57940 2252 57946 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 58880 2202
rect 1104 2128 58880 2150
rect 49970 1708 49976 1760
rect 50028 1748 50034 1760
rect 56502 1748 56508 1760
rect 50028 1720 56508 1748
rect 50028 1708 50034 1720
rect 56502 1708 56508 1720
rect 56560 1708 56566 1760
rect 52362 756 52368 808
rect 52420 796 52426 808
rect 56318 796 56324 808
rect 52420 768 56324 796
rect 52420 756 52426 768
rect 56318 756 56324 768
rect 56376 756 56382 808
<< via1 >>
rect 55312 58624 55364 58676
rect 56416 58624 56468 58676
rect 53748 58012 53800 58064
rect 56508 58012 56560 58064
rect 27252 57876 27304 57928
rect 34244 57876 34296 57928
rect 27988 57808 28040 57860
rect 29828 57808 29880 57860
rect 30380 57808 30432 57860
rect 37096 57808 37148 57860
rect 26424 57740 26476 57792
rect 32312 57740 32364 57792
rect 33508 57740 33560 57792
rect 36268 57740 36320 57792
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 4068 57536 4120 57588
rect 4620 57536 4672 57588
rect 2780 57468 2832 57520
rect 11980 57468 12032 57520
rect 12164 57468 12216 57520
rect 24032 57536 24084 57588
rect 6644 57400 6696 57452
rect 4252 57375 4304 57384
rect 4252 57341 4261 57375
rect 4261 57341 4295 57375
rect 4295 57341 4304 57375
rect 4252 57332 4304 57341
rect 4804 57332 4856 57384
rect 5080 57332 5132 57384
rect 5908 57332 5960 57384
rect 1860 57307 1912 57316
rect 1860 57273 1869 57307
rect 1869 57273 1903 57307
rect 1903 57273 1912 57307
rect 1860 57264 1912 57273
rect 7472 57264 7524 57316
rect 9036 57332 9088 57384
rect 9772 57332 9824 57384
rect 11428 57332 11480 57384
rect 12256 57375 12308 57384
rect 12256 57341 12265 57375
rect 12265 57341 12299 57375
rect 12299 57341 12308 57375
rect 12256 57332 12308 57341
rect 26148 57468 26200 57520
rect 26700 57468 26752 57520
rect 26884 57511 26936 57520
rect 26884 57477 26893 57511
rect 26893 57477 26927 57511
rect 26927 57477 26936 57511
rect 26884 57468 26936 57477
rect 27068 57536 27120 57588
rect 29920 57536 29972 57588
rect 14556 57400 14608 57452
rect 11796 57264 11848 57316
rect 13820 57332 13872 57384
rect 15384 57400 15436 57452
rect 20076 57400 20128 57452
rect 16948 57332 17000 57384
rect 17960 57332 18012 57384
rect 18512 57332 18564 57384
rect 19340 57332 19392 57384
rect 20904 57400 20956 57452
rect 24216 57400 24268 57452
rect 28356 57400 28408 57452
rect 22100 57332 22152 57384
rect 24308 57375 24360 57384
rect 24308 57341 24317 57375
rect 24317 57341 24351 57375
rect 24351 57341 24360 57375
rect 24308 57332 24360 57341
rect 24584 57375 24636 57384
rect 24584 57341 24593 57375
rect 24593 57341 24627 57375
rect 24627 57341 24636 57375
rect 25964 57375 26016 57384
rect 24584 57332 24636 57341
rect 25964 57341 25973 57375
rect 25973 57341 26007 57375
rect 26007 57341 26016 57375
rect 25964 57332 26016 57341
rect 26332 57332 26384 57384
rect 33416 57468 33468 57520
rect 46940 57468 46992 57520
rect 55128 57468 55180 57520
rect 55680 57468 55732 57520
rect 29644 57400 29696 57452
rect 29828 57400 29880 57452
rect 29276 57332 29328 57384
rect 32128 57332 32180 57384
rect 32312 57375 32364 57384
rect 32312 57341 32321 57375
rect 32321 57341 32355 57375
rect 32355 57341 32364 57375
rect 32312 57332 32364 57341
rect 32680 57332 32732 57384
rect 20168 57264 20220 57316
rect 5540 57239 5592 57248
rect 5540 57205 5549 57239
rect 5549 57205 5583 57239
rect 5583 57205 5592 57239
rect 5540 57196 5592 57205
rect 11060 57196 11112 57248
rect 11244 57239 11296 57248
rect 11244 57205 11253 57239
rect 11253 57205 11287 57239
rect 11287 57205 11296 57239
rect 11244 57196 11296 57205
rect 12440 57239 12492 57248
rect 12440 57205 12449 57239
rect 12449 57205 12483 57239
rect 12483 57205 12492 57239
rect 12440 57196 12492 57205
rect 13636 57239 13688 57248
rect 13636 57205 13645 57239
rect 13645 57205 13679 57239
rect 13679 57205 13688 57239
rect 13636 57196 13688 57205
rect 15108 57196 15160 57248
rect 15568 57239 15620 57248
rect 15568 57205 15577 57239
rect 15577 57205 15611 57239
rect 15611 57205 15620 57239
rect 15568 57196 15620 57205
rect 15660 57196 15712 57248
rect 17960 57196 18012 57248
rect 18236 57239 18288 57248
rect 18236 57205 18245 57239
rect 18245 57205 18279 57239
rect 18279 57205 18288 57239
rect 18236 57196 18288 57205
rect 18880 57239 18932 57248
rect 18880 57205 18889 57239
rect 18889 57205 18923 57239
rect 18923 57205 18932 57239
rect 18880 57196 18932 57205
rect 20260 57239 20312 57248
rect 20260 57205 20269 57239
rect 20269 57205 20303 57239
rect 20303 57205 20312 57239
rect 20260 57196 20312 57205
rect 20352 57196 20404 57248
rect 21548 57239 21600 57248
rect 21548 57205 21557 57239
rect 21557 57205 21591 57239
rect 21591 57205 21600 57239
rect 21548 57196 21600 57205
rect 23020 57264 23072 57316
rect 26700 57264 26752 57316
rect 29000 57264 29052 57316
rect 29184 57264 29236 57316
rect 33784 57375 33836 57384
rect 33784 57341 33793 57375
rect 33793 57341 33827 57375
rect 33827 57341 33836 57375
rect 36636 57400 36688 57452
rect 33784 57332 33836 57341
rect 35256 57332 35308 57384
rect 36452 57375 36504 57384
rect 36452 57341 36461 57375
rect 36461 57341 36495 57375
rect 36495 57341 36504 57375
rect 36452 57332 36504 57341
rect 37096 57375 37148 57384
rect 37096 57341 37105 57375
rect 37105 57341 37139 57375
rect 37139 57341 37148 57375
rect 37096 57332 37148 57341
rect 39028 57400 39080 57452
rect 41420 57400 41472 57452
rect 24124 57239 24176 57248
rect 24124 57205 24133 57239
rect 24133 57205 24167 57239
rect 24167 57205 24176 57239
rect 24124 57196 24176 57205
rect 25872 57196 25924 57248
rect 26148 57196 26200 57248
rect 28264 57239 28316 57248
rect 28264 57205 28273 57239
rect 28273 57205 28307 57239
rect 28307 57205 28316 57239
rect 28264 57196 28316 57205
rect 31668 57196 31720 57248
rect 38200 57264 38252 57316
rect 40592 57332 40644 57384
rect 45376 57400 45428 57452
rect 42984 57375 43036 57384
rect 42984 57341 42993 57375
rect 42993 57341 43027 57375
rect 43027 57341 43036 57375
rect 42984 57332 43036 57341
rect 43720 57332 43772 57384
rect 44548 57332 44600 57384
rect 46112 57332 46164 57384
rect 49240 57400 49292 57452
rect 47676 57332 47728 57384
rect 48504 57332 48556 57384
rect 50068 57400 50120 57452
rect 56416 57400 56468 57452
rect 58164 57443 58216 57452
rect 58164 57409 58173 57443
rect 58173 57409 58207 57443
rect 58207 57409 58216 57443
rect 58164 57400 58216 57409
rect 53748 57332 53800 57384
rect 54116 57332 54168 57384
rect 56784 57332 56836 57384
rect 53104 57307 53156 57316
rect 53104 57273 53113 57307
rect 53113 57273 53147 57307
rect 53147 57273 53156 57307
rect 53104 57264 53156 57273
rect 34244 57239 34296 57248
rect 34244 57205 34253 57239
rect 34253 57205 34287 57239
rect 34287 57205 34296 57239
rect 34244 57196 34296 57205
rect 34612 57196 34664 57248
rect 36912 57239 36964 57248
rect 36912 57205 36921 57239
rect 36921 57205 36955 57239
rect 36955 57205 36964 57239
rect 36912 57196 36964 57205
rect 38936 57239 38988 57248
rect 38936 57205 38945 57239
rect 38945 57205 38979 57239
rect 38979 57205 38988 57239
rect 38936 57196 38988 57205
rect 39580 57239 39632 57248
rect 39580 57205 39589 57239
rect 39589 57205 39623 57239
rect 39623 57205 39632 57239
rect 39580 57196 39632 57205
rect 40408 57239 40460 57248
rect 40408 57205 40417 57239
rect 40417 57205 40451 57239
rect 40451 57205 40460 57239
rect 40408 57196 40460 57205
rect 57980 57307 58032 57316
rect 57980 57273 57989 57307
rect 57989 57273 58023 57307
rect 58023 57273 58032 57307
rect 57980 57264 58032 57273
rect 58348 57196 58400 57248
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 50326 57094 50378 57146
rect 50390 57094 50442 57146
rect 50454 57094 50506 57146
rect 50518 57094 50570 57146
rect 4252 56992 4304 57044
rect 8300 56924 8352 56976
rect 1400 56899 1452 56908
rect 1400 56865 1409 56899
rect 1409 56865 1443 56899
rect 1443 56865 1452 56899
rect 1400 56856 1452 56865
rect 2136 56899 2188 56908
rect 2136 56865 2145 56899
rect 2145 56865 2179 56899
rect 2179 56865 2188 56899
rect 2136 56856 2188 56865
rect 3148 56899 3200 56908
rect 3148 56865 3157 56899
rect 3157 56865 3191 56899
rect 3191 56865 3200 56899
rect 3148 56856 3200 56865
rect 3332 56856 3384 56908
rect 8208 56899 8260 56908
rect 8208 56865 8217 56899
rect 8217 56865 8251 56899
rect 8251 56865 8260 56899
rect 8208 56856 8260 56865
rect 10600 56856 10652 56908
rect 12256 56924 12308 56976
rect 12992 56924 13044 56976
rect 15568 56924 15620 56976
rect 11980 56899 12032 56908
rect 11980 56865 11989 56899
rect 11989 56865 12023 56899
rect 12023 56865 12032 56899
rect 11980 56856 12032 56865
rect 15660 56856 15712 56908
rect 16120 56856 16172 56908
rect 4620 56788 4672 56840
rect 11060 56788 11112 56840
rect 11796 56831 11848 56840
rect 11796 56797 11805 56831
rect 11805 56797 11839 56831
rect 11839 56797 11848 56831
rect 11796 56788 11848 56797
rect 12164 56831 12216 56840
rect 12164 56797 12173 56831
rect 12173 56797 12207 56831
rect 12207 56797 12216 56831
rect 12164 56788 12216 56797
rect 15108 56831 15160 56840
rect 15108 56797 15117 56831
rect 15117 56797 15151 56831
rect 15151 56797 15160 56831
rect 15108 56788 15160 56797
rect 13176 56720 13228 56772
rect 18236 56924 18288 56976
rect 21548 56924 21600 56976
rect 18880 56856 18932 56908
rect 17960 56831 18012 56840
rect 17960 56797 17969 56831
rect 17969 56797 18003 56831
rect 18003 56797 18012 56831
rect 17960 56788 18012 56797
rect 20168 56831 20220 56840
rect 20168 56797 20174 56831
rect 20174 56797 20220 56831
rect 20168 56788 20220 56797
rect 20352 56831 20404 56840
rect 20352 56797 20361 56831
rect 20361 56797 20395 56831
rect 20395 56797 20404 56831
rect 20352 56788 20404 56797
rect 26884 56992 26936 57044
rect 28264 56924 28316 56976
rect 22468 56856 22520 56908
rect 25872 56856 25924 56908
rect 26700 56899 26752 56908
rect 26700 56865 26709 56899
rect 26709 56865 26743 56899
rect 26743 56865 26752 56899
rect 26700 56856 26752 56865
rect 27252 56856 27304 56908
rect 27988 56899 28040 56908
rect 27988 56865 27997 56899
rect 27997 56865 28031 56899
rect 28031 56865 28040 56899
rect 27988 56856 28040 56865
rect 35900 56992 35952 57044
rect 29184 56924 29236 56976
rect 36912 56924 36964 56976
rect 23020 56788 23072 56840
rect 23388 56831 23440 56840
rect 23388 56797 23397 56831
rect 23397 56797 23431 56831
rect 23431 56797 23440 56831
rect 23388 56788 23440 56797
rect 26332 56788 26384 56840
rect 29920 56856 29972 56908
rect 31300 56899 31352 56908
rect 31300 56865 31334 56899
rect 31334 56865 31352 56899
rect 31300 56856 31352 56865
rect 35440 56856 35492 56908
rect 35900 56899 35952 56908
rect 35900 56865 35909 56899
rect 35909 56865 35943 56899
rect 35943 56865 35952 56899
rect 35900 56856 35952 56865
rect 53104 56992 53156 57044
rect 57980 56992 58032 57044
rect 57060 56967 57112 56976
rect 57060 56933 57069 56967
rect 57069 56933 57103 56967
rect 57103 56933 57112 56967
rect 57060 56924 57112 56933
rect 29184 56831 29236 56840
rect 29184 56797 29193 56831
rect 29193 56797 29227 56831
rect 29227 56797 29236 56831
rect 29184 56788 29236 56797
rect 29276 56831 29328 56840
rect 29276 56797 29285 56831
rect 29285 56797 29319 56831
rect 29319 56797 29328 56831
rect 29276 56788 29328 56797
rect 30748 56788 30800 56840
rect 33324 56831 33376 56840
rect 33324 56797 33333 56831
rect 33333 56797 33367 56831
rect 33367 56797 33376 56831
rect 33324 56788 33376 56797
rect 34428 56788 34480 56840
rect 37464 56856 37516 56908
rect 39764 56899 39816 56908
rect 39764 56865 39773 56899
rect 39773 56865 39807 56899
rect 39807 56865 39816 56899
rect 39764 56856 39816 56865
rect 42156 56899 42208 56908
rect 42156 56865 42165 56899
rect 42165 56865 42199 56899
rect 42199 56865 42208 56899
rect 42156 56856 42208 56865
rect 51080 56856 51132 56908
rect 51632 56856 51684 56908
rect 54116 56899 54168 56908
rect 54116 56865 54125 56899
rect 54125 56865 54159 56899
rect 54159 56865 54168 56899
rect 54116 56856 54168 56865
rect 57152 56856 57204 56908
rect 54576 56831 54628 56840
rect 54576 56797 54585 56831
rect 54585 56797 54619 56831
rect 54619 56797 54628 56831
rect 54576 56788 54628 56797
rect 54760 56831 54812 56840
rect 54760 56797 54769 56831
rect 54769 56797 54803 56831
rect 54803 56797 54812 56831
rect 54760 56788 54812 56797
rect 56600 56788 56652 56840
rect 3240 56695 3292 56704
rect 3240 56661 3249 56695
rect 3249 56661 3283 56695
rect 3283 56661 3292 56695
rect 3240 56652 3292 56661
rect 20260 56763 20312 56772
rect 20260 56729 20269 56763
rect 20269 56729 20303 56763
rect 20303 56729 20312 56763
rect 20260 56720 20312 56729
rect 29092 56763 29144 56772
rect 29092 56729 29101 56763
rect 29101 56729 29135 56763
rect 29135 56729 29144 56763
rect 29092 56720 29144 56729
rect 23112 56652 23164 56704
rect 25596 56695 25648 56704
rect 25596 56661 25605 56695
rect 25605 56661 25639 56695
rect 25639 56661 25648 56695
rect 25596 56652 25648 56661
rect 25964 56695 26016 56704
rect 25964 56661 25973 56695
rect 25973 56661 26007 56695
rect 26007 56661 26016 56695
rect 25964 56652 26016 56661
rect 27068 56652 27120 56704
rect 28908 56652 28960 56704
rect 29276 56652 29328 56704
rect 30288 56652 30340 56704
rect 32128 56720 32180 56772
rect 34336 56720 34388 56772
rect 55772 56720 55824 56772
rect 56416 56720 56468 56772
rect 32956 56652 33008 56704
rect 33140 56652 33192 56704
rect 34428 56652 34480 56704
rect 34796 56652 34848 56704
rect 35256 56652 35308 56704
rect 37648 56695 37700 56704
rect 37648 56661 37657 56695
rect 37657 56661 37691 56695
rect 37691 56661 37700 56695
rect 37648 56652 37700 56661
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 388 56448 440 56500
rect 1308 56448 1360 56500
rect 3240 56448 3292 56500
rect 4804 56491 4856 56500
rect 4804 56457 4813 56491
rect 4813 56457 4847 56491
rect 4847 56457 4856 56491
rect 4804 56448 4856 56457
rect 23388 56448 23440 56500
rect 24584 56448 24636 56500
rect 26332 56448 26384 56500
rect 26792 56448 26844 56500
rect 3332 56423 3384 56432
rect 3332 56389 3341 56423
rect 3341 56389 3375 56423
rect 3375 56389 3384 56423
rect 3332 56380 3384 56389
rect 4252 56380 4304 56432
rect 11796 56380 11848 56432
rect 31300 56448 31352 56500
rect 31944 56448 31996 56500
rect 33048 56448 33100 56500
rect 33232 56491 33284 56500
rect 33232 56457 33256 56491
rect 33256 56457 33284 56491
rect 33232 56448 33284 56457
rect 34704 56448 34756 56500
rect 35256 56448 35308 56500
rect 34428 56380 34480 56432
rect 38936 56448 38988 56500
rect 54760 56448 54812 56500
rect 56416 56448 56468 56500
rect 56508 56448 56560 56500
rect 59544 56448 59596 56500
rect 35624 56380 35676 56432
rect 53932 56380 53984 56432
rect 54668 56380 54720 56432
rect 56140 56380 56192 56432
rect 58072 56380 58124 56432
rect 1124 56312 1176 56364
rect 1216 56244 1268 56296
rect 4620 56312 4672 56364
rect 11980 56312 12032 56364
rect 33416 56355 33468 56364
rect 2688 56244 2740 56296
rect 5264 56244 5316 56296
rect 11244 56244 11296 56296
rect 12072 56287 12124 56296
rect 12072 56253 12081 56287
rect 12081 56253 12115 56287
rect 12115 56253 12124 56287
rect 12072 56244 12124 56253
rect 33416 56321 33425 56355
rect 33425 56321 33459 56355
rect 33459 56321 33468 56355
rect 33416 56312 33468 56321
rect 23204 56244 23256 56296
rect 23388 56244 23440 56296
rect 24124 56244 24176 56296
rect 25320 56287 25372 56296
rect 25320 56253 25329 56287
rect 25329 56253 25363 56287
rect 25363 56253 25372 56287
rect 25320 56244 25372 56253
rect 25596 56287 25648 56296
rect 25596 56253 25630 56287
rect 25630 56253 25648 56287
rect 25596 56244 25648 56253
rect 29092 56244 29144 56296
rect 31668 56287 31720 56296
rect 31668 56253 31677 56287
rect 31677 56253 31711 56287
rect 31711 56253 31720 56287
rect 31668 56244 31720 56253
rect 32128 56287 32180 56296
rect 32128 56253 32137 56287
rect 32137 56253 32171 56287
rect 32171 56253 32180 56287
rect 32128 56244 32180 56253
rect 32588 56244 32640 56296
rect 12716 56176 12768 56228
rect 27896 56176 27948 56228
rect 4160 56151 4212 56160
rect 4160 56117 4169 56151
rect 4169 56117 4203 56151
rect 4203 56117 4212 56151
rect 4160 56108 4212 56117
rect 27344 56108 27396 56160
rect 29000 56108 29052 56160
rect 30472 56176 30524 56228
rect 31392 56176 31444 56228
rect 30840 56108 30892 56160
rect 31576 56108 31628 56160
rect 32036 56176 32088 56228
rect 33048 56219 33100 56228
rect 33048 56185 33057 56219
rect 33057 56185 33091 56219
rect 33091 56185 33100 56219
rect 33048 56176 33100 56185
rect 33416 56176 33468 56228
rect 34428 56287 34480 56296
rect 34428 56253 34437 56287
rect 34437 56253 34471 56287
rect 34471 56253 34480 56287
rect 34428 56244 34480 56253
rect 34796 56287 34848 56296
rect 34520 56176 34572 56228
rect 34796 56253 34805 56287
rect 34805 56253 34839 56287
rect 34839 56253 34848 56287
rect 34796 56244 34848 56253
rect 55772 56355 55824 56364
rect 55772 56321 55781 56355
rect 55781 56321 55815 56355
rect 55815 56321 55824 56355
rect 55772 56312 55824 56321
rect 56232 56355 56284 56364
rect 56232 56321 56241 56355
rect 56241 56321 56275 56355
rect 56275 56321 56284 56355
rect 56232 56312 56284 56321
rect 36268 56287 36320 56296
rect 36268 56253 36277 56287
rect 36277 56253 36311 56287
rect 36311 56253 36320 56287
rect 36268 56244 36320 56253
rect 52460 56287 52512 56296
rect 34980 56108 35032 56160
rect 36084 56151 36136 56160
rect 36084 56117 36093 56151
rect 36093 56117 36127 56151
rect 36127 56117 36136 56151
rect 36084 56108 36136 56117
rect 52460 56253 52469 56287
rect 52469 56253 52503 56287
rect 52503 56253 52512 56287
rect 52460 56244 52512 56253
rect 54300 56244 54352 56296
rect 56692 56176 56744 56228
rect 58716 56108 58768 56160
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 50326 56006 50378 56058
rect 50390 56006 50442 56058
rect 50454 56006 50506 56058
rect 50518 56006 50570 56058
rect 3148 55904 3200 55956
rect 4160 55904 4212 55956
rect 13360 55904 13412 55956
rect 24308 55947 24360 55956
rect 24308 55913 24317 55947
rect 24317 55913 24351 55947
rect 24351 55913 24360 55947
rect 25964 55947 26016 55956
rect 24308 55904 24360 55913
rect 1400 55811 1452 55820
rect 1400 55777 1409 55811
rect 1409 55777 1443 55811
rect 1443 55777 1452 55811
rect 1400 55768 1452 55777
rect 1952 55768 2004 55820
rect 3516 55768 3568 55820
rect 24216 55768 24268 55820
rect 24584 55768 24636 55820
rect 25228 55811 25280 55820
rect 25228 55777 25237 55811
rect 25237 55777 25271 55811
rect 25271 55777 25280 55811
rect 25228 55768 25280 55777
rect 25964 55913 25973 55947
rect 25973 55913 26007 55947
rect 26007 55913 26016 55947
rect 25964 55904 26016 55913
rect 27896 55947 27948 55956
rect 27896 55913 27905 55947
rect 27905 55913 27939 55947
rect 27939 55913 27948 55947
rect 27896 55904 27948 55913
rect 30472 55947 30524 55956
rect 30472 55913 30481 55947
rect 30481 55913 30515 55947
rect 30515 55913 30524 55947
rect 30472 55904 30524 55913
rect 27896 55768 27948 55820
rect 27988 55768 28040 55820
rect 32128 55904 32180 55956
rect 33140 55904 33192 55956
rect 33232 55904 33284 55956
rect 56784 55947 56836 55956
rect 56784 55913 56793 55947
rect 56793 55913 56827 55947
rect 56827 55913 56836 55947
rect 56784 55904 56836 55913
rect 28264 55768 28316 55820
rect 29000 55811 29052 55820
rect 29000 55777 29009 55811
rect 29009 55777 29043 55811
rect 29043 55777 29052 55811
rect 29000 55768 29052 55777
rect 32036 55836 32088 55888
rect 31392 55811 31444 55820
rect 1860 55700 1912 55752
rect 4252 55675 4304 55684
rect 4252 55641 4261 55675
rect 4261 55641 4295 55675
rect 4295 55641 4304 55675
rect 4252 55632 4304 55641
rect 27436 55700 27488 55752
rect 30380 55700 30432 55752
rect 31392 55777 31401 55811
rect 31401 55777 31435 55811
rect 31435 55777 31444 55811
rect 31392 55768 31444 55777
rect 31576 55811 31628 55820
rect 31576 55777 31585 55811
rect 31585 55777 31619 55811
rect 31619 55777 31628 55811
rect 31576 55768 31628 55777
rect 34796 55836 34848 55888
rect 33692 55811 33744 55820
rect 33692 55777 33726 55811
rect 33726 55777 33744 55811
rect 33692 55768 33744 55777
rect 34152 55768 34204 55820
rect 57244 55836 57296 55888
rect 53196 55811 53248 55820
rect 53196 55777 53205 55811
rect 53205 55777 53239 55811
rect 53239 55777 53248 55811
rect 53196 55768 53248 55777
rect 54024 55768 54076 55820
rect 54576 55768 54628 55820
rect 56600 55768 56652 55820
rect 56692 55768 56744 55820
rect 33232 55700 33284 55752
rect 56048 55700 56100 55752
rect 57704 55743 57756 55752
rect 57704 55709 57713 55743
rect 57713 55709 57747 55743
rect 57747 55709 57756 55743
rect 57704 55700 57756 55709
rect 26516 55607 26568 55616
rect 26516 55573 26525 55607
rect 26525 55573 26559 55607
rect 26559 55573 26568 55607
rect 26516 55564 26568 55573
rect 26884 55607 26936 55616
rect 26884 55573 26893 55607
rect 26893 55573 26927 55607
rect 26927 55573 26936 55607
rect 26884 55564 26936 55573
rect 28264 55607 28316 55616
rect 28264 55573 28273 55607
rect 28273 55573 28307 55607
rect 28307 55573 28316 55607
rect 28264 55564 28316 55573
rect 28724 55564 28776 55616
rect 31944 55564 31996 55616
rect 32220 55607 32272 55616
rect 32220 55573 32229 55607
rect 32229 55573 32263 55607
rect 32263 55573 32272 55607
rect 32220 55564 32272 55573
rect 56232 55632 56284 55684
rect 34796 55607 34848 55616
rect 34796 55573 34805 55607
rect 34805 55573 34839 55607
rect 34839 55573 34848 55607
rect 34796 55564 34848 55573
rect 57980 55607 58032 55616
rect 57980 55573 57989 55607
rect 57989 55573 58023 55607
rect 58023 55573 58032 55607
rect 57980 55564 58032 55573
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 30840 55360 30892 55412
rect 56048 55403 56100 55412
rect 22836 55292 22888 55344
rect 23388 55292 23440 55344
rect 56048 55369 56057 55403
rect 56057 55369 56091 55403
rect 56091 55369 56100 55403
rect 56048 55360 56100 55369
rect 57336 55403 57388 55412
rect 57336 55369 57345 55403
rect 57345 55369 57379 55403
rect 57379 55369 57388 55403
rect 57336 55360 57388 55369
rect 33508 55292 33560 55344
rect 24768 55224 24820 55276
rect 32036 55267 32088 55276
rect 22928 55199 22980 55208
rect 22928 55165 22937 55199
rect 22937 55165 22971 55199
rect 22971 55165 22980 55199
rect 22928 55156 22980 55165
rect 23388 55156 23440 55208
rect 32036 55233 32045 55267
rect 32045 55233 32079 55267
rect 32079 55233 32088 55267
rect 32036 55224 32088 55233
rect 32864 55224 32916 55276
rect 33416 55267 33468 55276
rect 33416 55233 33425 55267
rect 33425 55233 33459 55267
rect 33459 55233 33468 55267
rect 33416 55224 33468 55233
rect 34520 55292 34572 55344
rect 57704 55292 57756 55344
rect 58164 55335 58216 55344
rect 58164 55301 58173 55335
rect 58173 55301 58207 55335
rect 58207 55301 58216 55335
rect 58164 55292 58216 55301
rect 33876 55267 33928 55276
rect 33876 55233 33885 55267
rect 33885 55233 33919 55267
rect 33919 55233 33928 55267
rect 33876 55224 33928 55233
rect 34060 55224 34112 55276
rect 25872 55156 25924 55208
rect 26884 55156 26936 55208
rect 23296 55088 23348 55140
rect 23848 55088 23900 55140
rect 27896 55131 27948 55140
rect 22560 55063 22612 55072
rect 22560 55029 22569 55063
rect 22569 55029 22603 55063
rect 22603 55029 22612 55063
rect 22560 55020 22612 55029
rect 23112 55020 23164 55072
rect 24308 55020 24360 55072
rect 27896 55097 27905 55131
rect 27905 55097 27939 55131
rect 27939 55097 27948 55131
rect 27896 55088 27948 55097
rect 27436 55020 27488 55072
rect 29000 55199 29052 55208
rect 29000 55165 29009 55199
rect 29009 55165 29043 55199
rect 29043 55165 29052 55199
rect 29000 55156 29052 55165
rect 32220 55156 32272 55208
rect 33508 55199 33560 55208
rect 29092 55088 29144 55140
rect 29552 55020 29604 55072
rect 32588 55088 32640 55140
rect 33508 55165 33517 55199
rect 33517 55165 33551 55199
rect 33551 55165 33560 55199
rect 33508 55156 33560 55165
rect 34704 55156 34756 55208
rect 53932 55156 53984 55208
rect 55220 55199 55272 55208
rect 55220 55165 55229 55199
rect 55229 55165 55263 55199
rect 55263 55165 55272 55199
rect 56692 55199 56744 55208
rect 55220 55156 55272 55165
rect 56692 55165 56701 55199
rect 56701 55165 56735 55199
rect 56735 55165 56744 55199
rect 56692 55156 56744 55165
rect 57980 55199 58032 55208
rect 57980 55165 57989 55199
rect 57989 55165 58023 55199
rect 58023 55165 58032 55199
rect 57980 55156 58032 55165
rect 34244 55088 34296 55140
rect 35256 55088 35308 55140
rect 58532 55088 58584 55140
rect 33416 55020 33468 55072
rect 36176 55063 36228 55072
rect 36176 55029 36185 55063
rect 36185 55029 36219 55063
rect 36219 55029 36228 55063
rect 36176 55020 36228 55029
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 50326 54918 50378 54970
rect 50390 54918 50442 54970
rect 50454 54918 50506 54970
rect 50518 54918 50570 54970
rect 23388 54859 23440 54868
rect 8300 54748 8352 54800
rect 22560 54748 22612 54800
rect 23388 54825 23397 54859
rect 23397 54825 23431 54859
rect 23431 54825 23440 54859
rect 23388 54816 23440 54825
rect 23848 54859 23900 54868
rect 23848 54825 23857 54859
rect 23857 54825 23891 54859
rect 23891 54825 23900 54859
rect 23848 54816 23900 54825
rect 27436 54859 27488 54868
rect 27436 54825 27445 54859
rect 27445 54825 27479 54859
rect 27479 54825 27488 54859
rect 27436 54816 27488 54825
rect 28264 54816 28316 54868
rect 32036 54816 32088 54868
rect 1400 54723 1452 54732
rect 1400 54689 1409 54723
rect 1409 54689 1443 54723
rect 1443 54689 1452 54723
rect 1400 54680 1452 54689
rect 22100 54680 22152 54732
rect 22836 54680 22888 54732
rect 24308 54723 24360 54732
rect 24308 54689 24317 54723
rect 24317 54689 24351 54723
rect 24351 54689 24360 54723
rect 24308 54680 24360 54689
rect 25320 54680 25372 54732
rect 26148 54680 26200 54732
rect 26516 54748 26568 54800
rect 27896 54723 27948 54732
rect 27896 54689 27905 54723
rect 27905 54689 27939 54723
rect 27939 54689 27948 54723
rect 27896 54680 27948 54689
rect 31760 54748 31812 54800
rect 33140 54816 33192 54868
rect 58348 54816 58400 54868
rect 32588 54723 32640 54732
rect 25228 54612 25280 54664
rect 32588 54689 32597 54723
rect 32597 54689 32631 54723
rect 32631 54689 32640 54723
rect 32588 54680 32640 54689
rect 29368 54612 29420 54664
rect 30748 54655 30800 54664
rect 30748 54621 30757 54655
rect 30757 54621 30791 54655
rect 30791 54621 30800 54655
rect 30748 54612 30800 54621
rect 32864 54723 32916 54732
rect 32864 54689 32873 54723
rect 32873 54689 32907 54723
rect 32907 54689 32916 54723
rect 32864 54680 32916 54689
rect 33048 54680 33100 54732
rect 37648 54748 37700 54800
rect 34152 54723 34204 54732
rect 34152 54689 34161 54723
rect 34161 54689 34195 54723
rect 34195 54689 34204 54723
rect 34152 54680 34204 54689
rect 36176 54680 36228 54732
rect 56140 54748 56192 54800
rect 55312 54680 55364 54732
rect 55588 54723 55640 54732
rect 55588 54689 55597 54723
rect 55597 54689 55631 54723
rect 55631 54689 55640 54723
rect 55588 54680 55640 54689
rect 34796 54612 34848 54664
rect 29920 54544 29972 54596
rect 23940 54476 23992 54528
rect 28540 54519 28592 54528
rect 28540 54485 28549 54519
rect 28549 54485 28583 54519
rect 28583 54485 28592 54519
rect 28540 54476 28592 54485
rect 28908 54519 28960 54528
rect 28908 54485 28917 54519
rect 28917 54485 28951 54519
rect 28951 54485 28960 54519
rect 28908 54476 28960 54485
rect 31760 54544 31812 54596
rect 33692 54544 33744 54596
rect 57704 54655 57756 54664
rect 57704 54621 57713 54655
rect 57713 54621 57747 54655
rect 57747 54621 57756 54655
rect 57704 54612 57756 54621
rect 35440 54544 35492 54596
rect 33232 54476 33284 54528
rect 33876 54476 33928 54528
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 22928 54272 22980 54324
rect 23296 54315 23348 54324
rect 23296 54281 23305 54315
rect 23305 54281 23339 54315
rect 23339 54281 23348 54315
rect 23296 54272 23348 54281
rect 23940 54315 23992 54324
rect 23940 54281 23949 54315
rect 23949 54281 23983 54315
rect 23983 54281 23992 54315
rect 23940 54272 23992 54281
rect 25228 54272 25280 54324
rect 29092 54272 29144 54324
rect 33692 54272 33744 54324
rect 35256 54315 35308 54324
rect 35256 54281 35265 54315
rect 35265 54281 35299 54315
rect 35299 54281 35308 54315
rect 35256 54272 35308 54281
rect 57704 54272 57756 54324
rect 1400 54111 1452 54120
rect 1400 54077 1409 54111
rect 1409 54077 1443 54111
rect 1443 54077 1452 54111
rect 1400 54068 1452 54077
rect 22192 54068 22244 54120
rect 23388 54111 23440 54120
rect 23388 54077 23397 54111
rect 23397 54077 23431 54111
rect 23431 54077 23440 54111
rect 23388 54068 23440 54077
rect 24308 54136 24360 54188
rect 24768 54068 24820 54120
rect 25412 54068 25464 54120
rect 27712 54136 27764 54188
rect 29184 54111 29236 54120
rect 29184 54077 29193 54111
rect 29193 54077 29227 54111
rect 29227 54077 29236 54111
rect 29184 54068 29236 54077
rect 29368 54111 29420 54120
rect 29368 54077 29377 54111
rect 29377 54077 29411 54111
rect 29411 54077 29420 54111
rect 29368 54068 29420 54077
rect 29552 54068 29604 54120
rect 29920 54068 29972 54120
rect 31484 54111 31536 54120
rect 31484 54077 31493 54111
rect 31493 54077 31527 54111
rect 31527 54077 31536 54111
rect 31484 54068 31536 54077
rect 33048 54111 33100 54120
rect 33048 54077 33057 54111
rect 33057 54077 33091 54111
rect 33091 54077 33100 54111
rect 33048 54068 33100 54077
rect 39580 54204 39632 54256
rect 58164 54247 58216 54256
rect 58164 54213 58173 54247
rect 58173 54213 58207 54247
rect 58207 54213 58216 54247
rect 58164 54204 58216 54213
rect 35900 54179 35952 54188
rect 35900 54145 35909 54179
rect 35909 54145 35943 54179
rect 35943 54145 35952 54179
rect 35900 54136 35952 54145
rect 33600 54111 33652 54120
rect 27896 54043 27948 54052
rect 27896 54009 27905 54043
rect 27905 54009 27939 54043
rect 27939 54009 27948 54043
rect 27896 54000 27948 54009
rect 28908 54000 28960 54052
rect 32864 54000 32916 54052
rect 33140 54000 33192 54052
rect 33600 54077 33609 54111
rect 33609 54077 33643 54111
rect 33643 54077 33652 54111
rect 33600 54068 33652 54077
rect 35440 54111 35492 54120
rect 35440 54077 35449 54111
rect 35449 54077 35483 54111
rect 35483 54077 35492 54111
rect 35440 54068 35492 54077
rect 36176 54068 36228 54120
rect 8300 53932 8352 53984
rect 8852 53932 8904 53984
rect 25596 53932 25648 53984
rect 26424 53975 26476 53984
rect 26424 53941 26433 53975
rect 26433 53941 26467 53975
rect 26467 53941 26476 53975
rect 26424 53932 26476 53941
rect 32956 53932 33008 53984
rect 33324 53932 33376 53984
rect 33508 54000 33560 54052
rect 33784 53975 33836 53984
rect 33784 53941 33793 53975
rect 33793 53941 33827 53975
rect 33827 53941 33836 53975
rect 33784 53932 33836 53941
rect 36084 54000 36136 54052
rect 36360 54111 36412 54120
rect 36360 54077 36369 54111
rect 36369 54077 36403 54111
rect 36403 54077 36412 54111
rect 36360 54068 36412 54077
rect 55680 54068 55732 54120
rect 57336 54068 57388 54120
rect 57428 54111 57480 54120
rect 57428 54077 57437 54111
rect 57437 54077 57471 54111
rect 57471 54077 57480 54111
rect 57428 54068 57480 54077
rect 57980 54043 58032 54052
rect 57980 54009 57989 54043
rect 57989 54009 58023 54043
rect 58023 54009 58032 54043
rect 57980 54000 58032 54009
rect 36360 53932 36412 53984
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 50326 53830 50378 53882
rect 50390 53830 50442 53882
rect 50454 53830 50506 53882
rect 50518 53830 50570 53882
rect 27712 53771 27764 53780
rect 27712 53737 27721 53771
rect 27721 53737 27755 53771
rect 27755 53737 27764 53771
rect 27712 53728 27764 53737
rect 29368 53728 29420 53780
rect 33600 53728 33652 53780
rect 56968 53771 57020 53780
rect 56968 53737 56977 53771
rect 56977 53737 57011 53771
rect 57011 53737 57020 53771
rect 56968 53728 57020 53737
rect 57980 53728 58032 53780
rect 22100 53660 22152 53712
rect 26424 53660 26476 53712
rect 28540 53660 28592 53712
rect 30656 53660 30708 53712
rect 21732 53592 21784 53644
rect 23572 53592 23624 53644
rect 24768 53592 24820 53644
rect 25412 53635 25464 53644
rect 25412 53601 25421 53635
rect 25421 53601 25455 53635
rect 25455 53601 25464 53635
rect 25412 53592 25464 53601
rect 25596 53635 25648 53644
rect 25596 53601 25605 53635
rect 25605 53601 25639 53635
rect 25639 53601 25648 53635
rect 25596 53592 25648 53601
rect 26148 53592 26200 53644
rect 26332 53635 26384 53644
rect 26332 53601 26341 53635
rect 26341 53601 26375 53635
rect 26375 53601 26384 53635
rect 26332 53592 26384 53601
rect 29000 53592 29052 53644
rect 30932 53635 30984 53644
rect 30932 53601 30966 53635
rect 30966 53601 30984 53635
rect 31300 53660 31352 53712
rect 30932 53592 30984 53601
rect 33232 53592 33284 53644
rect 33784 53660 33836 53712
rect 57796 53660 57848 53712
rect 34612 53592 34664 53644
rect 35900 53635 35952 53644
rect 35900 53601 35909 53635
rect 35909 53601 35943 53635
rect 35943 53601 35952 53635
rect 35900 53592 35952 53601
rect 36176 53635 36228 53644
rect 36176 53601 36185 53635
rect 36185 53601 36219 53635
rect 36219 53601 36228 53635
rect 36176 53592 36228 53601
rect 56508 53592 56560 53644
rect 57336 53592 57388 53644
rect 23940 53567 23992 53576
rect 23940 53533 23949 53567
rect 23949 53533 23983 53567
rect 23983 53533 23992 53567
rect 23940 53524 23992 53533
rect 26056 53524 26108 53576
rect 30012 53524 30064 53576
rect 57704 53567 57756 53576
rect 57704 53533 57713 53567
rect 57713 53533 57747 53567
rect 57747 53533 57756 53567
rect 57704 53524 57756 53533
rect 31760 53456 31812 53508
rect 22560 53431 22612 53440
rect 22560 53397 22569 53431
rect 22569 53397 22603 53431
rect 22603 53397 22612 53431
rect 22560 53388 22612 53397
rect 23480 53431 23532 53440
rect 23480 53397 23489 53431
rect 23489 53397 23523 53431
rect 23523 53397 23532 53431
rect 23480 53388 23532 53397
rect 23664 53388 23716 53440
rect 25228 53431 25280 53440
rect 25228 53397 25237 53431
rect 25237 53397 25271 53431
rect 25271 53397 25280 53431
rect 25228 53388 25280 53397
rect 32036 53431 32088 53440
rect 32036 53397 32045 53431
rect 32045 53397 32079 53431
rect 32079 53397 32088 53431
rect 32036 53388 32088 53397
rect 32220 53388 32272 53440
rect 33876 53388 33928 53440
rect 35716 53431 35768 53440
rect 35716 53397 35725 53431
rect 35725 53397 35759 53431
rect 35759 53397 35768 53431
rect 35716 53388 35768 53397
rect 36360 53388 36412 53440
rect 36728 53388 36780 53440
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 11888 53184 11940 53236
rect 22192 53116 22244 53168
rect 26056 53159 26108 53168
rect 26056 53125 26065 53159
rect 26065 53125 26099 53159
rect 26099 53125 26108 53159
rect 26056 53116 26108 53125
rect 29184 53184 29236 53236
rect 29920 53227 29972 53236
rect 29920 53193 29929 53227
rect 29929 53193 29963 53227
rect 29963 53193 29972 53227
rect 29920 53184 29972 53193
rect 30932 53184 30984 53236
rect 34152 53184 34204 53236
rect 33048 53116 33100 53168
rect 36176 53184 36228 53236
rect 57704 53184 57756 53236
rect 22100 53048 22152 53100
rect 22836 53091 22888 53100
rect 22836 53057 22845 53091
rect 22845 53057 22879 53091
rect 22879 53057 22888 53091
rect 22836 53048 22888 53057
rect 1400 53023 1452 53032
rect 1400 52989 1409 53023
rect 1409 52989 1443 53023
rect 1443 52989 1452 53023
rect 1400 52980 1452 52989
rect 21456 53023 21508 53032
rect 21456 52989 21465 53023
rect 21465 52989 21499 53023
rect 21499 52989 21508 53023
rect 21456 52980 21508 52989
rect 22560 52980 22612 53032
rect 23480 52980 23532 53032
rect 25228 52980 25280 53032
rect 25688 52980 25740 53032
rect 29368 53048 29420 53100
rect 27896 53023 27948 53032
rect 27896 52989 27905 53023
rect 27905 52989 27939 53023
rect 27939 52989 27948 53023
rect 27896 52980 27948 52989
rect 29552 52980 29604 53032
rect 30748 53048 30800 53100
rect 30656 53023 30708 53032
rect 30656 52989 30663 53023
rect 30663 52989 30708 53023
rect 25320 52912 25372 52964
rect 25412 52912 25464 52964
rect 28908 52912 28960 52964
rect 30656 52980 30708 52989
rect 32036 53048 32088 53100
rect 31668 52980 31720 53032
rect 23112 52844 23164 52896
rect 23940 52844 23992 52896
rect 30656 52844 30708 52896
rect 31300 52912 31352 52964
rect 31944 52980 31996 53032
rect 33048 53023 33100 53032
rect 33048 52989 33057 53023
rect 33057 52989 33091 53023
rect 33091 52989 33100 53023
rect 33048 52980 33100 52989
rect 40408 53116 40460 53168
rect 32220 52912 32272 52964
rect 33140 52912 33192 52964
rect 32128 52844 32180 52896
rect 33324 52844 33376 52896
rect 33508 52980 33560 53032
rect 34704 53023 34756 53032
rect 34704 52989 34713 53023
rect 34713 52989 34747 53023
rect 34747 52989 34756 53023
rect 34704 52980 34756 52989
rect 35716 52980 35768 53032
rect 56508 52980 56560 53032
rect 57520 52980 57572 53032
rect 57980 52955 58032 52964
rect 57980 52921 57989 52955
rect 57989 52921 58023 52955
rect 58023 52921 58032 52955
rect 57980 52912 58032 52921
rect 58164 52955 58216 52964
rect 58164 52921 58173 52955
rect 58173 52921 58207 52955
rect 58207 52921 58216 52955
rect 58164 52912 58216 52921
rect 33784 52887 33836 52896
rect 33784 52853 33793 52887
rect 33793 52853 33827 52887
rect 33827 52853 33836 52887
rect 33784 52844 33836 52853
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 50326 52742 50378 52794
rect 50390 52742 50442 52794
rect 50454 52742 50506 52794
rect 50518 52742 50570 52794
rect 21732 52683 21784 52692
rect 21732 52649 21741 52683
rect 21741 52649 21775 52683
rect 21775 52649 21784 52683
rect 21732 52640 21784 52649
rect 22192 52640 22244 52692
rect 23480 52640 23532 52692
rect 23664 52683 23716 52692
rect 23664 52649 23673 52683
rect 23673 52649 23707 52683
rect 23707 52649 23716 52683
rect 23664 52640 23716 52649
rect 31484 52640 31536 52692
rect 20904 52504 20956 52556
rect 22560 52504 22612 52556
rect 29092 52572 29144 52624
rect 30380 52572 30432 52624
rect 23112 52547 23164 52556
rect 23112 52513 23121 52547
rect 23121 52513 23155 52547
rect 23155 52513 23164 52547
rect 23112 52504 23164 52513
rect 23756 52504 23808 52556
rect 21456 52436 21508 52488
rect 26148 52504 26200 52556
rect 30012 52504 30064 52556
rect 30656 52547 30708 52556
rect 30656 52513 30665 52547
rect 30665 52513 30699 52547
rect 30699 52513 30708 52547
rect 30656 52504 30708 52513
rect 32036 52547 32088 52556
rect 32036 52513 32045 52547
rect 32045 52513 32079 52547
rect 32079 52513 32088 52547
rect 32036 52504 32088 52513
rect 32588 52504 32640 52556
rect 33232 52640 33284 52692
rect 36728 52683 36780 52692
rect 36728 52649 36737 52683
rect 36737 52649 36771 52683
rect 36771 52649 36780 52683
rect 36728 52640 36780 52649
rect 57980 52640 58032 52692
rect 33784 52572 33836 52624
rect 34060 52504 34112 52556
rect 34336 52504 34388 52556
rect 36268 52504 36320 52556
rect 26240 52436 26292 52488
rect 25688 52343 25740 52352
rect 25688 52309 25697 52343
rect 25697 52309 25731 52343
rect 25731 52309 25740 52343
rect 25688 52300 25740 52309
rect 29276 52300 29328 52352
rect 36084 52436 36136 52488
rect 57704 52479 57756 52488
rect 57704 52445 57713 52479
rect 57713 52445 57747 52479
rect 57747 52445 57756 52479
rect 57704 52436 57756 52445
rect 33508 52300 33560 52352
rect 35716 52343 35768 52352
rect 35716 52309 35725 52343
rect 35725 52309 35759 52343
rect 35759 52309 35768 52343
rect 35716 52300 35768 52309
rect 36176 52300 36228 52352
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 25964 52139 26016 52148
rect 25964 52105 25973 52139
rect 25973 52105 26007 52139
rect 26007 52105 26016 52139
rect 25964 52096 26016 52105
rect 26332 52096 26384 52148
rect 32036 52096 32088 52148
rect 36268 52139 36320 52148
rect 36268 52105 36277 52139
rect 36277 52105 36311 52139
rect 36311 52105 36320 52139
rect 36268 52096 36320 52105
rect 57704 52096 57756 52148
rect 32128 52071 32180 52080
rect 32128 52037 32137 52071
rect 32137 52037 32171 52071
rect 32171 52037 32180 52071
rect 32128 52028 32180 52037
rect 58164 52071 58216 52080
rect 58164 52037 58173 52071
rect 58173 52037 58207 52071
rect 58207 52037 58216 52071
rect 58164 52028 58216 52037
rect 21364 51960 21416 52012
rect 22836 51960 22888 52012
rect 33600 52003 33652 52012
rect 1400 51935 1452 51944
rect 1400 51901 1409 51935
rect 1409 51901 1443 51935
rect 1443 51901 1452 51935
rect 1400 51892 1452 51901
rect 20904 51892 20956 51944
rect 21456 51935 21508 51944
rect 21456 51901 21465 51935
rect 21465 51901 21499 51935
rect 21499 51901 21508 51935
rect 21456 51892 21508 51901
rect 23296 51935 23348 51944
rect 23296 51901 23305 51935
rect 23305 51901 23339 51935
rect 23339 51901 23348 51935
rect 23296 51892 23348 51901
rect 23664 51892 23716 51944
rect 24032 51892 24084 51944
rect 28172 51935 28224 51944
rect 23756 51824 23808 51876
rect 25044 51824 25096 51876
rect 28172 51901 28181 51935
rect 28181 51901 28215 51935
rect 28215 51901 28224 51935
rect 28172 51892 28224 51901
rect 28632 51892 28684 51944
rect 21088 51799 21140 51808
rect 21088 51765 21097 51799
rect 21097 51765 21131 51799
rect 21131 51765 21140 51799
rect 21088 51756 21140 51765
rect 22928 51799 22980 51808
rect 22928 51765 22937 51799
rect 22937 51765 22971 51799
rect 22971 51765 22980 51799
rect 22928 51756 22980 51765
rect 25596 51756 25648 51808
rect 28816 51824 28868 51876
rect 25872 51756 25924 51808
rect 26148 51799 26200 51808
rect 26148 51765 26157 51799
rect 26157 51765 26191 51799
rect 26191 51765 26200 51799
rect 26148 51756 26200 51765
rect 27804 51799 27856 51808
rect 27804 51765 27813 51799
rect 27813 51765 27847 51799
rect 27847 51765 27856 51799
rect 27804 51756 27856 51765
rect 29644 51892 29696 51944
rect 30012 51935 30064 51944
rect 30012 51901 30021 51935
rect 30021 51901 30055 51935
rect 30055 51901 30064 51935
rect 30012 51892 30064 51901
rect 33600 51969 33609 52003
rect 33609 51969 33643 52003
rect 33643 51969 33652 52003
rect 33600 51960 33652 51969
rect 31760 51892 31812 51944
rect 33416 51935 33468 51944
rect 33416 51901 33425 51935
rect 33425 51901 33459 51935
rect 33459 51901 33468 51935
rect 33416 51892 33468 51901
rect 34336 51935 34388 51944
rect 34336 51901 34345 51935
rect 34345 51901 34379 51935
rect 34379 51901 34388 51935
rect 34336 51892 34388 51901
rect 35716 51892 35768 51944
rect 36176 51935 36228 51944
rect 36176 51901 36185 51935
rect 36185 51901 36219 51935
rect 36219 51901 36228 51935
rect 36176 51892 36228 51901
rect 29184 51867 29236 51876
rect 29184 51833 29193 51867
rect 29193 51833 29227 51867
rect 29227 51833 29236 51867
rect 29184 51824 29236 51833
rect 29276 51867 29328 51876
rect 29276 51833 29285 51867
rect 29285 51833 29319 51867
rect 29319 51833 29328 51867
rect 29276 51824 29328 51833
rect 29552 51756 29604 51808
rect 32588 51824 32640 51876
rect 33508 51799 33560 51808
rect 33508 51765 33517 51799
rect 33517 51765 33551 51799
rect 33551 51765 33560 51799
rect 36084 51824 36136 51876
rect 56508 51892 56560 51944
rect 57520 51892 57572 51944
rect 58348 51824 58400 51876
rect 33508 51756 33560 51765
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 50326 51654 50378 51706
rect 50390 51654 50442 51706
rect 50454 51654 50506 51706
rect 50518 51654 50570 51706
rect 23664 51595 23716 51604
rect 23664 51561 23673 51595
rect 23673 51561 23707 51595
rect 23707 51561 23716 51595
rect 23664 51552 23716 51561
rect 23756 51552 23808 51604
rect 25964 51552 26016 51604
rect 28632 51595 28684 51604
rect 28632 51561 28641 51595
rect 28641 51561 28675 51595
rect 28675 51561 28684 51595
rect 28632 51552 28684 51561
rect 29000 51552 29052 51604
rect 29092 51595 29144 51604
rect 29092 51561 29101 51595
rect 29101 51561 29135 51595
rect 29135 51561 29144 51595
rect 29092 51552 29144 51561
rect 33140 51552 33192 51604
rect 33508 51552 33560 51604
rect 21088 51484 21140 51536
rect 22928 51484 22980 51536
rect 25688 51527 25740 51536
rect 1400 51459 1452 51468
rect 1400 51425 1409 51459
rect 1409 51425 1443 51459
rect 1443 51425 1452 51459
rect 1400 51416 1452 51425
rect 22284 51459 22336 51468
rect 22284 51425 22293 51459
rect 22293 51425 22327 51459
rect 22327 51425 22336 51459
rect 22284 51416 22336 51425
rect 22836 51416 22888 51468
rect 23296 51416 23348 51468
rect 25688 51493 25722 51527
rect 25722 51493 25740 51527
rect 25688 51484 25740 51493
rect 27804 51484 27856 51536
rect 29552 51484 29604 51536
rect 20444 51391 20496 51400
rect 20444 51357 20453 51391
rect 20453 51357 20487 51391
rect 20487 51357 20496 51391
rect 20444 51348 20496 51357
rect 26148 51416 26200 51468
rect 29644 51416 29696 51468
rect 30564 51416 30616 51468
rect 30840 51416 30892 51468
rect 32312 51459 32364 51468
rect 32312 51425 32346 51459
rect 32346 51425 32364 51459
rect 32312 51416 32364 51425
rect 32588 51416 32640 51468
rect 57980 51459 58032 51468
rect 57980 51425 57989 51459
rect 57989 51425 58023 51459
rect 58023 51425 58032 51459
rect 57980 51416 58032 51425
rect 21364 51212 21416 51264
rect 29368 51348 29420 51400
rect 30656 51348 30708 51400
rect 31944 51348 31996 51400
rect 58164 51323 58216 51332
rect 58164 51289 58173 51323
rect 58173 51289 58207 51323
rect 58207 51289 58216 51323
rect 58164 51280 58216 51289
rect 26332 51212 26384 51264
rect 29184 51212 29236 51264
rect 57428 51255 57480 51264
rect 57428 51221 57437 51255
rect 57437 51221 57471 51255
rect 57471 51221 57480 51255
rect 57428 51212 57480 51221
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 20904 51051 20956 51060
rect 20904 51017 20913 51051
rect 20913 51017 20947 51051
rect 20947 51017 20956 51051
rect 20904 51008 20956 51017
rect 21456 51008 21508 51060
rect 25044 51051 25096 51060
rect 25044 51017 25053 51051
rect 25053 51017 25087 51051
rect 25087 51017 25096 51051
rect 25044 51008 25096 51017
rect 26240 51008 26292 51060
rect 28172 51008 28224 51060
rect 25872 50872 25924 50924
rect 21364 50804 21416 50856
rect 21640 50804 21692 50856
rect 24032 50804 24084 50856
rect 25504 50804 25556 50856
rect 25964 50804 26016 50856
rect 26700 50804 26752 50856
rect 28172 50847 28224 50856
rect 28172 50813 28181 50847
rect 28181 50813 28215 50847
rect 28215 50813 28224 50847
rect 28172 50804 28224 50813
rect 28816 51008 28868 51060
rect 29184 51008 29236 51060
rect 30564 51051 30616 51060
rect 29000 50847 29052 50856
rect 29000 50813 29009 50847
rect 29009 50813 29043 50847
rect 29043 50813 29052 50847
rect 29000 50804 29052 50813
rect 30564 51017 30573 51051
rect 30573 51017 30607 51051
rect 30607 51017 30616 51051
rect 30564 51008 30616 51017
rect 36176 51008 36228 51060
rect 57980 51051 58032 51060
rect 57980 51017 57989 51051
rect 57989 51017 58023 51051
rect 58023 51017 58032 51051
rect 57980 51008 58032 51017
rect 31484 50872 31536 50924
rect 30656 50847 30708 50856
rect 30656 50813 30665 50847
rect 30665 50813 30699 50847
rect 30699 50813 30708 50847
rect 30656 50804 30708 50813
rect 31852 50847 31904 50856
rect 31852 50813 31861 50847
rect 31861 50813 31895 50847
rect 31895 50813 31904 50847
rect 34796 50872 34848 50924
rect 31852 50804 31904 50813
rect 33232 50847 33284 50856
rect 33232 50813 33241 50847
rect 33241 50813 33275 50847
rect 33275 50813 33284 50847
rect 33232 50804 33284 50813
rect 32956 50736 33008 50788
rect 34704 50804 34756 50856
rect 57428 50872 57480 50924
rect 57520 50736 57572 50788
rect 22284 50668 22336 50720
rect 22652 50711 22704 50720
rect 22652 50677 22661 50711
rect 22661 50677 22695 50711
rect 22695 50677 22704 50711
rect 22652 50668 22704 50677
rect 25872 50668 25924 50720
rect 31392 50711 31444 50720
rect 31392 50677 31401 50711
rect 31401 50677 31435 50711
rect 31435 50677 31444 50711
rect 31392 50668 31444 50677
rect 34152 50711 34204 50720
rect 34152 50677 34161 50711
rect 34161 50677 34195 50711
rect 34195 50677 34204 50711
rect 34152 50668 34204 50677
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 50326 50566 50378 50618
rect 50390 50566 50442 50618
rect 50454 50566 50506 50618
rect 50518 50566 50570 50618
rect 24032 50464 24084 50516
rect 31852 50507 31904 50516
rect 31852 50473 31861 50507
rect 31861 50473 31895 50507
rect 31895 50473 31904 50507
rect 31852 50464 31904 50473
rect 32312 50507 32364 50516
rect 32312 50473 32321 50507
rect 32321 50473 32355 50507
rect 32355 50473 32364 50507
rect 32312 50464 32364 50473
rect 1400 50371 1452 50380
rect 1400 50337 1409 50371
rect 1409 50337 1443 50371
rect 1443 50337 1452 50371
rect 1400 50328 1452 50337
rect 21272 50328 21324 50380
rect 21456 50371 21508 50380
rect 21456 50337 21490 50371
rect 21490 50337 21508 50371
rect 21456 50328 21508 50337
rect 23480 50328 23532 50380
rect 25504 50328 25556 50380
rect 25872 50328 25924 50380
rect 26700 50328 26752 50380
rect 28172 50396 28224 50448
rect 31392 50396 31444 50448
rect 33232 50464 33284 50516
rect 34796 50507 34848 50516
rect 34796 50473 34805 50507
rect 34805 50473 34839 50507
rect 34839 50473 34848 50507
rect 34796 50464 34848 50473
rect 33508 50396 33560 50448
rect 34152 50396 34204 50448
rect 58164 50439 58216 50448
rect 58164 50405 58173 50439
rect 58173 50405 58207 50439
rect 58207 50405 58216 50439
rect 58164 50396 58216 50405
rect 20812 50260 20864 50312
rect 19432 50192 19484 50244
rect 20444 50192 20496 50244
rect 20168 50167 20220 50176
rect 20168 50133 20177 50167
rect 20177 50133 20211 50167
rect 20211 50133 20220 50167
rect 20168 50124 20220 50133
rect 20536 50167 20588 50176
rect 20536 50133 20545 50167
rect 20545 50133 20579 50167
rect 20579 50133 20588 50167
rect 20536 50124 20588 50133
rect 22652 50192 22704 50244
rect 22560 50167 22612 50176
rect 22560 50133 22569 50167
rect 22569 50133 22603 50167
rect 22603 50133 22612 50167
rect 25780 50167 25832 50176
rect 22560 50124 22612 50133
rect 25780 50133 25789 50167
rect 25789 50133 25823 50167
rect 25823 50133 25832 50167
rect 25780 50124 25832 50133
rect 27896 50167 27948 50176
rect 27896 50133 27905 50167
rect 27905 50133 27939 50167
rect 27939 50133 27948 50167
rect 27896 50124 27948 50133
rect 29000 50371 29052 50380
rect 29000 50337 29009 50371
rect 29009 50337 29043 50371
rect 29043 50337 29052 50371
rect 29000 50328 29052 50337
rect 30012 50328 30064 50380
rect 31944 50328 31996 50380
rect 32496 50371 32548 50380
rect 32496 50337 32505 50371
rect 32505 50337 32539 50371
rect 32539 50337 32548 50371
rect 32496 50328 32548 50337
rect 32956 50371 33008 50380
rect 31484 50260 31536 50312
rect 32956 50337 32965 50371
rect 32965 50337 32999 50371
rect 32999 50337 33008 50371
rect 32956 50328 33008 50337
rect 57244 50371 57296 50380
rect 57244 50337 57253 50371
rect 57253 50337 57287 50371
rect 57287 50337 57296 50371
rect 57244 50328 57296 50337
rect 58256 50328 58308 50380
rect 31944 50192 31996 50244
rect 28356 50124 28408 50176
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 20812 49963 20864 49972
rect 20812 49929 20821 49963
rect 20821 49929 20855 49963
rect 20855 49929 20864 49963
rect 20812 49920 20864 49929
rect 21272 49920 21324 49972
rect 19432 49827 19484 49836
rect 19432 49793 19441 49827
rect 19441 49793 19475 49827
rect 19475 49793 19484 49827
rect 19432 49784 19484 49793
rect 29000 49920 29052 49972
rect 31484 49920 31536 49972
rect 32496 49920 32548 49972
rect 34336 49920 34388 49972
rect 20168 49716 20220 49768
rect 20536 49716 20588 49768
rect 22652 49784 22704 49836
rect 31116 49784 31168 49836
rect 33140 49784 33192 49836
rect 25228 49716 25280 49768
rect 25780 49759 25832 49768
rect 25780 49725 25814 49759
rect 25814 49725 25832 49759
rect 25780 49716 25832 49725
rect 26332 49716 26384 49768
rect 27528 49716 27580 49768
rect 27896 49716 27948 49768
rect 30472 49716 30524 49768
rect 31484 49716 31536 49768
rect 31668 49759 31720 49768
rect 31668 49725 31677 49759
rect 31677 49725 31711 49759
rect 31711 49725 31720 49759
rect 31668 49716 31720 49725
rect 30932 49648 30984 49700
rect 31760 49648 31812 49700
rect 33508 49716 33560 49768
rect 34244 49716 34296 49768
rect 34704 49759 34756 49768
rect 34704 49725 34713 49759
rect 34713 49725 34747 49759
rect 34747 49725 34756 49759
rect 34704 49716 34756 49725
rect 57520 49716 57572 49768
rect 58164 49759 58216 49768
rect 58164 49725 58173 49759
rect 58173 49725 58207 49759
rect 58207 49725 58216 49759
rect 58164 49716 58216 49725
rect 57980 49691 58032 49700
rect 57980 49657 57989 49691
rect 57989 49657 58023 49691
rect 58023 49657 58032 49691
rect 57980 49648 58032 49657
rect 22376 49580 22428 49632
rect 24952 49623 25004 49632
rect 24952 49589 24961 49623
rect 24961 49589 24995 49623
rect 24995 49589 25004 49623
rect 24952 49580 25004 49589
rect 26516 49580 26568 49632
rect 34612 49623 34664 49632
rect 34612 49589 34621 49623
rect 34621 49589 34655 49623
rect 34655 49589 34664 49623
rect 34612 49580 34664 49589
rect 57244 49623 57296 49632
rect 57244 49589 57253 49623
rect 57253 49589 57287 49623
rect 57287 49589 57296 49623
rect 57244 49580 57296 49589
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 50326 49478 50378 49530
rect 50390 49478 50442 49530
rect 50454 49478 50506 49530
rect 50518 49478 50570 49530
rect 21456 49419 21508 49428
rect 21456 49385 21465 49419
rect 21465 49385 21499 49419
rect 21499 49385 21508 49419
rect 21456 49376 21508 49385
rect 25228 49419 25280 49428
rect 25228 49385 25237 49419
rect 25237 49385 25271 49419
rect 25271 49385 25280 49419
rect 25228 49376 25280 49385
rect 26700 49419 26752 49428
rect 26700 49385 26709 49419
rect 26709 49385 26743 49419
rect 26743 49385 26752 49419
rect 26700 49376 26752 49385
rect 28356 49376 28408 49428
rect 1400 49283 1452 49292
rect 1400 49249 1409 49283
rect 1409 49249 1443 49283
rect 1443 49249 1452 49283
rect 1400 49240 1452 49249
rect 21640 49283 21692 49292
rect 21640 49249 21649 49283
rect 21649 49249 21683 49283
rect 21683 49249 21692 49283
rect 21640 49240 21692 49249
rect 22376 49283 22428 49292
rect 22376 49249 22385 49283
rect 22385 49249 22419 49283
rect 22419 49249 22428 49283
rect 22376 49240 22428 49249
rect 22560 49283 22612 49292
rect 22560 49249 22569 49283
rect 22569 49249 22603 49283
rect 22603 49249 22612 49283
rect 22560 49240 22612 49249
rect 24952 49240 25004 49292
rect 25688 49240 25740 49292
rect 25780 49215 25832 49224
rect 25780 49181 25789 49215
rect 25789 49181 25823 49215
rect 25823 49181 25832 49215
rect 29276 49283 29328 49292
rect 29276 49249 29285 49283
rect 29285 49249 29319 49283
rect 29319 49249 29328 49283
rect 29276 49240 29328 49249
rect 34796 49419 34848 49428
rect 34796 49385 34805 49419
rect 34805 49385 34839 49419
rect 34839 49385 34848 49419
rect 34796 49376 34848 49385
rect 57980 49376 58032 49428
rect 34428 49351 34480 49360
rect 31300 49283 31352 49292
rect 31300 49249 31334 49283
rect 31334 49249 31352 49283
rect 31300 49240 31352 49249
rect 27436 49215 27488 49224
rect 25780 49172 25832 49181
rect 27436 49181 27445 49215
rect 27445 49181 27479 49215
rect 27479 49181 27488 49215
rect 27436 49172 27488 49181
rect 30656 49172 30708 49224
rect 34428 49317 34463 49351
rect 34463 49317 34480 49351
rect 34428 49308 34480 49317
rect 35256 49308 35308 49360
rect 55036 49240 55088 49292
rect 57244 49240 57296 49292
rect 33692 49172 33744 49224
rect 26516 49079 26568 49088
rect 26516 49045 26525 49079
rect 26525 49045 26559 49079
rect 26559 49045 26568 49079
rect 26516 49036 26568 49045
rect 28448 49036 28500 49088
rect 31760 49036 31812 49088
rect 33324 49079 33376 49088
rect 33324 49045 33333 49079
rect 33333 49045 33367 49079
rect 33367 49045 33376 49079
rect 33324 49036 33376 49045
rect 57428 49172 57480 49224
rect 57060 49147 57112 49156
rect 57060 49113 57069 49147
rect 57069 49113 57103 49147
rect 57103 49113 57112 49147
rect 57060 49104 57112 49113
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 20444 48875 20496 48884
rect 20444 48841 20453 48875
rect 20453 48841 20487 48875
rect 20487 48841 20496 48875
rect 20444 48832 20496 48841
rect 20536 48832 20588 48884
rect 25504 48875 25556 48884
rect 25504 48841 25513 48875
rect 25513 48841 25547 48875
rect 25547 48841 25556 48875
rect 25504 48832 25556 48841
rect 30472 48875 30524 48884
rect 30472 48841 30481 48875
rect 30481 48841 30515 48875
rect 30515 48841 30524 48875
rect 30472 48832 30524 48841
rect 30932 48832 30984 48884
rect 31668 48832 31720 48884
rect 34428 48875 34480 48884
rect 34428 48841 34437 48875
rect 34437 48841 34471 48875
rect 34471 48841 34480 48875
rect 34428 48832 34480 48841
rect 35256 48832 35308 48884
rect 57428 48875 57480 48884
rect 57428 48841 57437 48875
rect 57437 48841 57471 48875
rect 57471 48841 57480 48875
rect 57428 48832 57480 48841
rect 18144 48671 18196 48680
rect 18144 48637 18153 48671
rect 18153 48637 18187 48671
rect 18187 48637 18196 48671
rect 18144 48628 18196 48637
rect 21088 48671 21140 48680
rect 21088 48637 21097 48671
rect 21097 48637 21131 48671
rect 21131 48637 21140 48671
rect 21088 48628 21140 48637
rect 27528 48696 27580 48748
rect 30656 48764 30708 48816
rect 24860 48671 24912 48680
rect 24860 48637 24869 48671
rect 24869 48637 24903 48671
rect 24903 48637 24912 48671
rect 24860 48628 24912 48637
rect 25688 48671 25740 48680
rect 25688 48637 25697 48671
rect 25697 48637 25731 48671
rect 25731 48637 25740 48671
rect 25688 48628 25740 48637
rect 25780 48671 25832 48680
rect 25780 48637 25789 48671
rect 25789 48637 25823 48671
rect 25823 48637 25832 48671
rect 26700 48671 26752 48680
rect 25780 48628 25832 48637
rect 26700 48637 26709 48671
rect 26709 48637 26743 48671
rect 26743 48637 26752 48671
rect 26700 48628 26752 48637
rect 27804 48671 27856 48680
rect 27804 48637 27813 48671
rect 27813 48637 27847 48671
rect 27847 48637 27856 48671
rect 27804 48628 27856 48637
rect 28448 48671 28500 48680
rect 28448 48637 28457 48671
rect 28457 48637 28491 48671
rect 28491 48637 28500 48671
rect 28448 48628 28500 48637
rect 31116 48671 31168 48680
rect 31116 48637 31125 48671
rect 31125 48637 31159 48671
rect 31159 48637 31168 48671
rect 31116 48628 31168 48637
rect 34336 48696 34388 48748
rect 18420 48603 18472 48612
rect 18420 48569 18454 48603
rect 18454 48569 18472 48603
rect 18420 48560 18472 48569
rect 19340 48492 19392 48544
rect 20352 48560 20404 48612
rect 20536 48560 20588 48612
rect 26516 48560 26568 48612
rect 33324 48671 33376 48680
rect 33324 48637 33358 48671
rect 33358 48637 33376 48671
rect 33324 48628 33376 48637
rect 56508 48628 56560 48680
rect 34612 48560 34664 48612
rect 57980 48603 58032 48612
rect 57980 48569 57989 48603
rect 57989 48569 58023 48603
rect 58023 48569 58032 48603
rect 57980 48560 58032 48569
rect 21180 48535 21232 48544
rect 21180 48501 21189 48535
rect 21189 48501 21223 48535
rect 21223 48501 21232 48535
rect 21180 48492 21232 48501
rect 26608 48492 26660 48544
rect 27712 48492 27764 48544
rect 28540 48535 28592 48544
rect 28540 48501 28549 48535
rect 28549 48501 28583 48535
rect 28583 48501 28592 48535
rect 28540 48492 28592 48501
rect 57888 48492 57940 48544
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 50326 48390 50378 48442
rect 50390 48390 50442 48442
rect 50454 48390 50506 48442
rect 50518 48390 50570 48442
rect 18420 48331 18472 48340
rect 18420 48297 18429 48331
rect 18429 48297 18463 48331
rect 18463 48297 18472 48331
rect 18420 48288 18472 48297
rect 31300 48331 31352 48340
rect 1400 48195 1452 48204
rect 1400 48161 1409 48195
rect 1409 48161 1443 48195
rect 1443 48161 1452 48195
rect 1400 48152 1452 48161
rect 16488 48220 16540 48272
rect 31300 48297 31309 48331
rect 31309 48297 31343 48331
rect 31343 48297 31352 48331
rect 31300 48288 31352 48297
rect 33692 48331 33744 48340
rect 33692 48297 33701 48331
rect 33701 48297 33735 48331
rect 33735 48297 33744 48331
rect 33692 48288 33744 48297
rect 34428 48331 34480 48340
rect 34428 48297 34437 48331
rect 34437 48297 34471 48331
rect 34471 48297 34480 48331
rect 34428 48288 34480 48297
rect 57980 48288 58032 48340
rect 16120 48152 16172 48204
rect 15016 47991 15068 48000
rect 15016 47957 15025 47991
rect 15025 47957 15059 47991
rect 15059 47957 15068 47991
rect 15016 47948 15068 47957
rect 15752 48084 15804 48136
rect 17960 48152 18012 48204
rect 21180 48220 21232 48272
rect 19340 48152 19392 48204
rect 19432 48084 19484 48136
rect 24216 48152 24268 48204
rect 25320 48152 25372 48204
rect 27528 48220 27580 48272
rect 28540 48220 28592 48272
rect 30932 48220 30984 48272
rect 26332 48152 26384 48204
rect 31484 48195 31536 48204
rect 25136 48084 25188 48136
rect 27712 48084 27764 48136
rect 31484 48161 31493 48195
rect 31493 48161 31527 48195
rect 31527 48161 31536 48195
rect 31484 48152 31536 48161
rect 31668 48195 31720 48204
rect 31668 48161 31677 48195
rect 31677 48161 31711 48195
rect 31711 48161 31720 48195
rect 31668 48152 31720 48161
rect 31760 48195 31812 48204
rect 31760 48161 31769 48195
rect 31769 48161 31803 48195
rect 31803 48161 31812 48195
rect 32220 48195 32272 48204
rect 31760 48152 31812 48161
rect 32220 48161 32229 48195
rect 32229 48161 32263 48195
rect 32263 48161 32272 48195
rect 32220 48152 32272 48161
rect 33048 48195 33100 48204
rect 33048 48161 33057 48195
rect 33057 48161 33091 48195
rect 33091 48161 33100 48195
rect 33048 48152 33100 48161
rect 33692 48152 33744 48204
rect 35256 48220 35308 48272
rect 31852 48084 31904 48136
rect 57704 48127 57756 48136
rect 57704 48093 57713 48127
rect 57713 48093 57747 48127
rect 57747 48093 57756 48127
rect 57704 48084 57756 48093
rect 20444 48016 20496 48068
rect 23480 48059 23532 48068
rect 23480 48025 23489 48059
rect 23489 48025 23523 48059
rect 23523 48025 23532 48059
rect 23480 48016 23532 48025
rect 27804 48016 27856 48068
rect 16396 47991 16448 48000
rect 16396 47957 16405 47991
rect 16405 47957 16439 47991
rect 16439 47957 16448 47991
rect 16396 47948 16448 47957
rect 17408 47948 17460 48000
rect 20536 47948 20588 48000
rect 24860 47948 24912 48000
rect 25412 47948 25464 48000
rect 29276 48016 29328 48068
rect 34244 48059 34296 48068
rect 34244 48025 34253 48059
rect 34253 48025 34287 48059
rect 34287 48025 34296 48059
rect 34244 48016 34296 48025
rect 28080 47991 28132 48000
rect 28080 47957 28089 47991
rect 28089 47957 28123 47991
rect 28123 47957 28132 47991
rect 28080 47948 28132 47957
rect 28264 47948 28316 48000
rect 29920 47948 29972 48000
rect 31760 47948 31812 48000
rect 31944 47948 31996 48000
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 16488 47744 16540 47796
rect 21088 47744 21140 47796
rect 25320 47787 25372 47796
rect 25320 47753 25329 47787
rect 25329 47753 25363 47787
rect 25363 47753 25372 47787
rect 25320 47744 25372 47753
rect 26332 47787 26384 47796
rect 26332 47753 26341 47787
rect 26341 47753 26375 47787
rect 26375 47753 26384 47787
rect 26332 47744 26384 47753
rect 26700 47744 26752 47796
rect 28080 47744 28132 47796
rect 29920 47787 29972 47796
rect 18788 47608 18840 47660
rect 27804 47676 27856 47728
rect 29920 47753 29929 47787
rect 29929 47753 29963 47787
rect 29963 47753 29972 47787
rect 29920 47744 29972 47753
rect 1400 47583 1452 47592
rect 1400 47549 1409 47583
rect 1409 47549 1443 47583
rect 1443 47549 1452 47583
rect 1400 47540 1452 47549
rect 13912 47540 13964 47592
rect 15016 47540 15068 47592
rect 17408 47540 17460 47592
rect 19156 47583 19208 47592
rect 19156 47549 19165 47583
rect 19165 47549 19199 47583
rect 19199 47549 19208 47583
rect 19156 47540 19208 47549
rect 19340 47583 19392 47592
rect 19340 47549 19349 47583
rect 19349 47549 19383 47583
rect 19383 47549 19392 47583
rect 19340 47540 19392 47549
rect 20352 47583 20404 47592
rect 20352 47549 20361 47583
rect 20361 47549 20395 47583
rect 20395 47549 20404 47583
rect 20352 47540 20404 47549
rect 20444 47583 20496 47592
rect 20444 47549 20453 47583
rect 20453 47549 20487 47583
rect 20487 47549 20496 47583
rect 20444 47540 20496 47549
rect 18144 47472 18196 47524
rect 19432 47472 19484 47524
rect 20536 47472 20588 47524
rect 23572 47540 23624 47592
rect 32220 47744 32272 47796
rect 57704 47744 57756 47796
rect 26608 47583 26660 47592
rect 26608 47549 26617 47583
rect 26617 47549 26651 47583
rect 26651 47549 26660 47583
rect 26608 47540 26660 47549
rect 27712 47540 27764 47592
rect 25228 47472 25280 47524
rect 15752 47447 15804 47456
rect 15752 47413 15761 47447
rect 15761 47413 15795 47447
rect 15795 47413 15804 47447
rect 15752 47404 15804 47413
rect 27896 47583 27948 47592
rect 27896 47549 27905 47583
rect 27905 47549 27939 47583
rect 27939 47549 27948 47583
rect 27896 47540 27948 47549
rect 29736 47583 29788 47592
rect 27988 47472 28040 47524
rect 29736 47549 29745 47583
rect 29745 47549 29779 47583
rect 29779 47549 29788 47583
rect 29736 47540 29788 47549
rect 30288 47540 30340 47592
rect 30472 47540 30524 47592
rect 30656 47583 30708 47592
rect 30656 47549 30665 47583
rect 30665 47549 30699 47583
rect 30699 47549 30708 47583
rect 30656 47540 30708 47549
rect 33508 47583 33560 47592
rect 31024 47472 31076 47524
rect 33508 47549 33517 47583
rect 33517 47549 33551 47583
rect 33551 47549 33560 47583
rect 33508 47540 33560 47549
rect 34336 47540 34388 47592
rect 57520 47540 57572 47592
rect 57704 47540 57756 47592
rect 33692 47472 33744 47524
rect 34244 47472 34296 47524
rect 55680 47472 55732 47524
rect 58164 47515 58216 47524
rect 58164 47481 58173 47515
rect 58173 47481 58207 47515
rect 58207 47481 58216 47515
rect 58164 47472 58216 47481
rect 28448 47404 28500 47456
rect 29552 47447 29604 47456
rect 29552 47413 29561 47447
rect 29561 47413 29595 47447
rect 29595 47413 29604 47447
rect 29552 47404 29604 47413
rect 32036 47447 32088 47456
rect 32036 47413 32045 47447
rect 32045 47413 32079 47447
rect 32079 47413 32088 47447
rect 32036 47404 32088 47413
rect 33140 47447 33192 47456
rect 33140 47413 33149 47447
rect 33149 47413 33183 47447
rect 33183 47413 33192 47447
rect 33140 47404 33192 47413
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 50326 47302 50378 47354
rect 50390 47302 50442 47354
rect 50454 47302 50506 47354
rect 50518 47302 50570 47354
rect 15752 47200 15804 47252
rect 24216 47243 24268 47252
rect 24216 47209 24225 47243
rect 24225 47209 24259 47243
rect 24259 47209 24268 47243
rect 24216 47200 24268 47209
rect 25228 47243 25280 47252
rect 25228 47209 25237 47243
rect 25237 47209 25271 47243
rect 25271 47209 25280 47243
rect 25228 47200 25280 47209
rect 28356 47200 28408 47252
rect 29736 47200 29788 47252
rect 31024 47243 31076 47252
rect 31024 47209 31033 47243
rect 31033 47209 31067 47243
rect 31067 47209 31076 47243
rect 31024 47200 31076 47209
rect 33508 47200 33560 47252
rect 34244 47243 34296 47252
rect 16488 47132 16540 47184
rect 15384 47064 15436 47116
rect 16396 47107 16448 47116
rect 16396 47073 16405 47107
rect 16405 47073 16439 47107
rect 16439 47073 16448 47107
rect 16396 47064 16448 47073
rect 17040 47107 17092 47116
rect 15292 46996 15344 47048
rect 17040 47073 17049 47107
rect 17049 47073 17083 47107
rect 17083 47073 17092 47107
rect 17040 47064 17092 47073
rect 18788 47107 18840 47116
rect 18788 47073 18797 47107
rect 18797 47073 18831 47107
rect 18831 47073 18840 47107
rect 18788 47064 18840 47073
rect 19156 47064 19208 47116
rect 17960 46996 18012 47048
rect 19340 46996 19392 47048
rect 20168 47064 20220 47116
rect 21456 47064 21508 47116
rect 23480 47064 23532 47116
rect 20628 46996 20680 47048
rect 16120 46971 16172 46980
rect 16120 46937 16129 46971
rect 16129 46937 16163 46971
rect 16163 46937 16172 46971
rect 16120 46928 16172 46937
rect 22744 46971 22796 46980
rect 22744 46937 22753 46971
rect 22753 46937 22787 46971
rect 22787 46937 22796 46971
rect 22744 46928 22796 46937
rect 23480 46971 23532 46980
rect 23480 46937 23489 46971
rect 23489 46937 23523 46971
rect 23523 46937 23532 46971
rect 23480 46928 23532 46937
rect 25320 47132 25372 47184
rect 25412 47107 25464 47116
rect 25412 47073 25421 47107
rect 25421 47073 25455 47107
rect 25455 47073 25464 47107
rect 25412 47064 25464 47073
rect 26700 47064 26752 47116
rect 27620 46996 27672 47048
rect 27896 47064 27948 47116
rect 28264 47107 28316 47116
rect 28264 47073 28273 47107
rect 28273 47073 28307 47107
rect 28307 47073 28316 47107
rect 28264 47064 28316 47073
rect 28448 47107 28500 47116
rect 28448 47073 28457 47107
rect 28457 47073 28491 47107
rect 28491 47073 28500 47107
rect 28448 47064 28500 47073
rect 29920 47132 29972 47184
rect 30472 47132 30524 47184
rect 30288 47064 30340 47116
rect 32036 47064 32088 47116
rect 33140 47132 33192 47184
rect 34244 47209 34253 47243
rect 34253 47209 34287 47243
rect 34287 47209 34296 47243
rect 34244 47200 34296 47209
rect 57704 47243 57756 47252
rect 57704 47209 57713 47243
rect 57713 47209 57747 47243
rect 57747 47209 57756 47243
rect 57704 47200 57756 47209
rect 34336 47107 34388 47116
rect 34336 47073 34345 47107
rect 34345 47073 34379 47107
rect 34379 47073 34388 47107
rect 34336 47064 34388 47073
rect 56876 47107 56928 47116
rect 56876 47073 56885 47107
rect 56885 47073 56919 47107
rect 56919 47073 56928 47107
rect 56876 47064 56928 47073
rect 57612 47064 57664 47116
rect 31852 46996 31904 47048
rect 32312 47039 32364 47048
rect 32312 47005 32321 47039
rect 32321 47005 32355 47039
rect 32355 47005 32364 47039
rect 32312 46996 32364 47005
rect 24768 46928 24820 46980
rect 27804 46928 27856 46980
rect 27988 46928 28040 46980
rect 31944 46928 31996 46980
rect 14740 46903 14792 46912
rect 14740 46869 14749 46903
rect 14749 46869 14783 46903
rect 14783 46869 14792 46903
rect 14740 46860 14792 46869
rect 15108 46903 15160 46912
rect 15108 46869 15117 46903
rect 15117 46869 15151 46903
rect 15151 46869 15160 46903
rect 15108 46860 15160 46869
rect 17776 46860 17828 46912
rect 18604 46903 18656 46912
rect 18604 46869 18613 46903
rect 18613 46869 18647 46903
rect 18647 46869 18656 46903
rect 18604 46860 18656 46869
rect 20076 46903 20128 46912
rect 20076 46869 20085 46903
rect 20085 46869 20119 46903
rect 20119 46869 20128 46903
rect 20076 46860 20128 46869
rect 22560 46860 22612 46912
rect 26608 46903 26660 46912
rect 26608 46869 26617 46903
rect 26617 46869 26651 46903
rect 26651 46869 26660 46903
rect 26608 46860 26660 46869
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 15108 46656 15160 46708
rect 15384 46699 15436 46708
rect 15384 46665 15393 46699
rect 15393 46665 15427 46699
rect 15427 46665 15436 46699
rect 15384 46656 15436 46665
rect 16396 46656 16448 46708
rect 19156 46656 19208 46708
rect 20168 46656 20220 46708
rect 22468 46656 22520 46708
rect 27804 46699 27856 46708
rect 27804 46665 27813 46699
rect 27813 46665 27847 46699
rect 27847 46665 27856 46699
rect 27804 46656 27856 46665
rect 30288 46699 30340 46708
rect 30288 46665 30297 46699
rect 30297 46665 30331 46699
rect 30331 46665 30340 46699
rect 30288 46656 30340 46665
rect 31852 46656 31904 46708
rect 32404 46588 32456 46640
rect 19432 46563 19484 46572
rect 1400 46495 1452 46504
rect 1400 46461 1409 46495
rect 1409 46461 1443 46495
rect 1443 46461 1452 46495
rect 1400 46452 1452 46461
rect 14740 46452 14792 46504
rect 15108 46452 15160 46504
rect 15384 46452 15436 46504
rect 19432 46529 19441 46563
rect 19441 46529 19475 46563
rect 19475 46529 19484 46563
rect 19432 46520 19484 46529
rect 24676 46520 24728 46572
rect 16764 46452 16816 46504
rect 18604 46452 18656 46504
rect 20076 46452 20128 46504
rect 20904 46452 20956 46504
rect 23388 46495 23440 46504
rect 23388 46461 23397 46495
rect 23397 46461 23431 46495
rect 23431 46461 23440 46495
rect 23388 46452 23440 46461
rect 24768 46495 24820 46504
rect 13912 46384 13964 46436
rect 22560 46427 22612 46436
rect 22560 46393 22569 46427
rect 22569 46393 22603 46427
rect 22603 46393 22612 46427
rect 22560 46384 22612 46393
rect 22100 46316 22152 46368
rect 22836 46384 22888 46436
rect 24768 46461 24777 46495
rect 24777 46461 24811 46495
rect 24811 46461 24820 46495
rect 24768 46452 24820 46461
rect 24952 46495 25004 46504
rect 24952 46461 24961 46495
rect 24961 46461 24995 46495
rect 24995 46461 25004 46495
rect 24952 46452 25004 46461
rect 25044 46495 25096 46504
rect 25044 46461 25053 46495
rect 25053 46461 25087 46495
rect 25087 46461 25096 46495
rect 25044 46452 25096 46461
rect 26608 46452 26660 46504
rect 27988 46495 28040 46504
rect 27988 46461 27997 46495
rect 27997 46461 28031 46495
rect 28031 46461 28040 46495
rect 27988 46452 28040 46461
rect 31760 46520 31812 46572
rect 32312 46520 32364 46572
rect 58164 46563 58216 46572
rect 58164 46529 58173 46563
rect 58173 46529 58207 46563
rect 58207 46529 58216 46563
rect 58164 46520 58216 46529
rect 31484 46495 31536 46504
rect 31484 46461 31493 46495
rect 31493 46461 31527 46495
rect 31527 46461 31536 46495
rect 31484 46452 31536 46461
rect 31944 46495 31996 46504
rect 31944 46461 31953 46495
rect 31953 46461 31987 46495
rect 31987 46461 31996 46495
rect 31944 46452 31996 46461
rect 32036 46452 32088 46504
rect 28448 46384 28500 46436
rect 29552 46384 29604 46436
rect 31208 46427 31260 46436
rect 31208 46393 31217 46427
rect 31217 46393 31251 46427
rect 31251 46393 31260 46427
rect 31208 46384 31260 46393
rect 33508 46384 33560 46436
rect 57980 46427 58032 46436
rect 57980 46393 57989 46427
rect 57989 46393 58023 46427
rect 58023 46393 58032 46427
rect 57980 46384 58032 46393
rect 22928 46359 22980 46368
rect 22928 46325 22937 46359
rect 22937 46325 22971 46359
rect 22971 46325 22980 46359
rect 22928 46316 22980 46325
rect 23020 46316 23072 46368
rect 24584 46359 24636 46368
rect 24584 46325 24593 46359
rect 24593 46325 24627 46359
rect 24627 46325 24636 46359
rect 24584 46316 24636 46325
rect 27620 46316 27672 46368
rect 31392 46359 31444 46368
rect 31392 46325 31401 46359
rect 31401 46325 31435 46359
rect 31435 46325 31444 46359
rect 31392 46316 31444 46325
rect 33416 46316 33468 46368
rect 34336 46316 34388 46368
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 50326 46214 50378 46266
rect 50390 46214 50442 46266
rect 50454 46214 50506 46266
rect 50518 46214 50570 46266
rect 17040 46112 17092 46164
rect 19432 46112 19484 46164
rect 20628 46155 20680 46164
rect 20628 46121 20637 46155
rect 20637 46121 20671 46155
rect 20671 46121 20680 46155
rect 20628 46112 20680 46121
rect 21456 46155 21508 46164
rect 21456 46121 21465 46155
rect 21465 46121 21499 46155
rect 21499 46121 21508 46155
rect 21456 46112 21508 46121
rect 22100 46112 22152 46164
rect 25044 46112 25096 46164
rect 15384 45976 15436 46028
rect 17776 46019 17828 46028
rect 17776 45985 17785 46019
rect 17785 45985 17819 46019
rect 17819 45985 17828 46019
rect 17776 45976 17828 45985
rect 19892 45976 19944 46028
rect 20168 46019 20220 46028
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 22744 46044 22796 46096
rect 23020 46087 23072 46096
rect 23020 46053 23054 46087
rect 23054 46053 23072 46087
rect 23020 46044 23072 46053
rect 24584 46044 24636 46096
rect 22560 45976 22612 46028
rect 13912 45908 13964 45960
rect 17040 45908 17092 45960
rect 23480 45976 23532 46028
rect 24952 45976 25004 46028
rect 27436 45976 27488 46028
rect 29276 46044 29328 46096
rect 31208 46112 31260 46164
rect 33508 46155 33560 46164
rect 33508 46121 33517 46155
rect 33517 46121 33551 46155
rect 33551 46121 33560 46155
rect 33508 46112 33560 46121
rect 57980 46112 58032 46164
rect 33048 46044 33100 46096
rect 27804 45976 27856 46028
rect 30472 45976 30524 46028
rect 30656 46019 30708 46028
rect 30656 45985 30665 46019
rect 30665 45985 30699 46019
rect 30699 45985 30708 46019
rect 30656 45976 30708 45985
rect 32956 45976 33008 46028
rect 33416 46019 33468 46028
rect 33416 45985 33425 46019
rect 33425 45985 33459 46019
rect 33459 45985 33468 46019
rect 33416 45976 33468 45985
rect 17960 45883 18012 45892
rect 17960 45849 17969 45883
rect 17969 45849 18003 45883
rect 18003 45849 18012 45883
rect 17960 45840 18012 45849
rect 22100 45840 22152 45892
rect 22560 45840 22612 45892
rect 24676 45908 24728 45960
rect 57704 45951 57756 45960
rect 57704 45917 57713 45951
rect 57713 45917 57747 45951
rect 57747 45917 57756 45951
rect 57704 45908 57756 45917
rect 14832 45815 14884 45824
rect 14832 45781 14841 45815
rect 14841 45781 14875 45815
rect 14875 45781 14884 45815
rect 14832 45772 14884 45781
rect 18604 45815 18656 45824
rect 18604 45781 18613 45815
rect 18613 45781 18647 45815
rect 18647 45781 18656 45815
rect 18604 45772 18656 45781
rect 20076 45815 20128 45824
rect 20076 45781 20085 45815
rect 20085 45781 20119 45815
rect 20119 45781 20128 45815
rect 20076 45772 20128 45781
rect 22468 45772 22520 45824
rect 24768 45772 24820 45824
rect 29092 45815 29144 45824
rect 29092 45781 29101 45815
rect 29101 45781 29135 45815
rect 29135 45781 29144 45815
rect 29092 45772 29144 45781
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 15384 45611 15436 45620
rect 15384 45577 15393 45611
rect 15393 45577 15427 45611
rect 15427 45577 15436 45611
rect 15384 45568 15436 45577
rect 23388 45568 23440 45620
rect 24952 45568 25004 45620
rect 27804 45611 27856 45620
rect 27804 45577 27813 45611
rect 27813 45577 27847 45611
rect 27847 45577 27856 45611
rect 27804 45568 27856 45577
rect 31208 45568 31260 45620
rect 57704 45568 57756 45620
rect 17960 45500 18012 45552
rect 18604 45500 18656 45552
rect 31944 45500 31996 45552
rect 58164 45543 58216 45552
rect 14004 45475 14056 45484
rect 14004 45441 14013 45475
rect 14013 45441 14047 45475
rect 14047 45441 14056 45475
rect 14004 45432 14056 45441
rect 24308 45432 24360 45484
rect 29276 45475 29328 45484
rect 1400 45407 1452 45416
rect 1400 45373 1409 45407
rect 1409 45373 1443 45407
rect 1443 45373 1452 45407
rect 1400 45364 1452 45373
rect 14832 45364 14884 45416
rect 17592 45407 17644 45416
rect 17592 45373 17601 45407
rect 17601 45373 17635 45407
rect 17635 45373 17644 45407
rect 17592 45364 17644 45373
rect 18144 45364 18196 45416
rect 19432 45364 19484 45416
rect 20904 45407 20956 45416
rect 20904 45373 20913 45407
rect 20913 45373 20947 45407
rect 20947 45373 20956 45407
rect 20904 45364 20956 45373
rect 20996 45364 21048 45416
rect 21640 45364 21692 45416
rect 22468 45364 22520 45416
rect 22836 45407 22888 45416
rect 22836 45373 22845 45407
rect 22845 45373 22879 45407
rect 22879 45373 22888 45407
rect 22836 45364 22888 45373
rect 22928 45364 22980 45416
rect 23940 45364 23992 45416
rect 24216 45364 24268 45416
rect 26240 45407 26292 45416
rect 18696 45296 18748 45348
rect 22652 45296 22704 45348
rect 26240 45373 26249 45407
rect 26249 45373 26283 45407
rect 26283 45373 26292 45407
rect 26240 45364 26292 45373
rect 27712 45364 27764 45416
rect 29276 45441 29285 45475
rect 29285 45441 29319 45475
rect 29319 45441 29328 45475
rect 29276 45432 29328 45441
rect 32956 45432 33008 45484
rect 28448 45364 28500 45416
rect 29092 45364 29144 45416
rect 32404 45364 32456 45416
rect 58164 45509 58173 45543
rect 58173 45509 58207 45543
rect 58207 45509 58216 45543
rect 58164 45500 58216 45509
rect 56508 45364 56560 45416
rect 57336 45364 57388 45416
rect 26424 45339 26476 45348
rect 26424 45305 26433 45339
rect 26433 45305 26467 45339
rect 26467 45305 26476 45339
rect 26424 45296 26476 45305
rect 27988 45339 28040 45348
rect 27988 45305 27997 45339
rect 27997 45305 28031 45339
rect 28031 45305 28040 45339
rect 27988 45296 28040 45305
rect 30472 45296 30524 45348
rect 17408 45271 17460 45280
rect 17408 45237 17417 45271
rect 17417 45237 17451 45271
rect 17451 45237 17460 45271
rect 17408 45228 17460 45237
rect 19984 45271 20036 45280
rect 19984 45237 19993 45271
rect 19993 45237 20027 45271
rect 20027 45237 20036 45271
rect 19984 45228 20036 45237
rect 20168 45228 20220 45280
rect 20720 45271 20772 45280
rect 20720 45237 20729 45271
rect 20729 45237 20763 45271
rect 20763 45237 20772 45271
rect 20720 45228 20772 45237
rect 23388 45271 23440 45280
rect 23388 45237 23397 45271
rect 23397 45237 23431 45271
rect 23431 45237 23440 45271
rect 23388 45228 23440 45237
rect 24492 45271 24544 45280
rect 24492 45237 24501 45271
rect 24501 45237 24535 45271
rect 24535 45237 24544 45271
rect 24492 45228 24544 45237
rect 31392 45296 31444 45348
rect 31484 45339 31536 45348
rect 31484 45305 31514 45339
rect 31514 45305 31536 45339
rect 31484 45296 31536 45305
rect 58808 45296 58860 45348
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 50326 45126 50378 45178
rect 50390 45126 50442 45178
rect 50454 45126 50506 45178
rect 50518 45126 50570 45178
rect 18144 45067 18196 45076
rect 18144 45033 18153 45067
rect 18153 45033 18187 45067
rect 18187 45033 18196 45067
rect 18144 45024 18196 45033
rect 18696 45024 18748 45076
rect 21640 45067 21692 45076
rect 21640 45033 21649 45067
rect 21649 45033 21683 45067
rect 21683 45033 21692 45067
rect 21640 45024 21692 45033
rect 25136 45024 25188 45076
rect 27896 45067 27948 45076
rect 17408 44956 17460 45008
rect 1400 44931 1452 44940
rect 1400 44897 1409 44931
rect 1409 44897 1443 44931
rect 1443 44897 1452 44931
rect 1400 44888 1452 44897
rect 16764 44931 16816 44940
rect 16764 44897 16773 44931
rect 16773 44897 16807 44931
rect 16807 44897 16816 44931
rect 16764 44888 16816 44897
rect 20076 44956 20128 45008
rect 20352 44956 20404 45008
rect 20720 44956 20772 45008
rect 26424 44956 26476 45008
rect 27896 45033 27905 45067
rect 27905 45033 27939 45067
rect 27939 45033 27948 45067
rect 27896 45024 27948 45033
rect 30472 45067 30524 45076
rect 30472 45033 30481 45067
rect 30481 45033 30515 45067
rect 30515 45033 30524 45067
rect 30472 45024 30524 45033
rect 31484 45024 31536 45076
rect 19984 44888 20036 44940
rect 23388 44888 23440 44940
rect 24492 44888 24544 44940
rect 24676 44888 24728 44940
rect 19432 44820 19484 44872
rect 22928 44863 22980 44872
rect 22928 44829 22937 44863
rect 22937 44829 22971 44863
rect 22971 44829 22980 44863
rect 22928 44820 22980 44829
rect 23940 44820 23992 44872
rect 24308 44863 24360 44872
rect 24308 44829 24317 44863
rect 24317 44829 24351 44863
rect 24351 44829 24360 44863
rect 24308 44820 24360 44829
rect 19340 44752 19392 44804
rect 19892 44752 19944 44804
rect 27620 44888 27672 44940
rect 31944 44956 31996 45008
rect 33968 44956 34020 45008
rect 28908 44888 28960 44940
rect 29000 44820 29052 44872
rect 31392 44888 31444 44940
rect 32220 44931 32272 44940
rect 32220 44897 32229 44931
rect 32229 44897 32263 44931
rect 32263 44897 32272 44931
rect 32220 44888 32272 44897
rect 32312 44931 32364 44940
rect 32312 44897 32321 44931
rect 32321 44897 32355 44931
rect 32355 44897 32364 44931
rect 32312 44888 32364 44897
rect 56968 44888 57020 44940
rect 57612 44888 57664 44940
rect 57980 44931 58032 44940
rect 57980 44897 57989 44931
rect 57989 44897 58023 44931
rect 58023 44897 58032 44931
rect 57980 44888 58032 44897
rect 58164 44931 58216 44940
rect 58164 44897 58173 44931
rect 58173 44897 58207 44931
rect 58207 44897 58216 44931
rect 58164 44888 58216 44897
rect 30656 44752 30708 44804
rect 31484 44752 31536 44804
rect 32128 44752 32180 44804
rect 22652 44684 22704 44736
rect 23848 44727 23900 44736
rect 23848 44693 23857 44727
rect 23857 44693 23891 44727
rect 23891 44693 23900 44727
rect 23848 44684 23900 44693
rect 24216 44727 24268 44736
rect 24216 44693 24225 44727
rect 24225 44693 24259 44727
rect 24259 44693 24268 44727
rect 24216 44684 24268 44693
rect 27252 44727 27304 44736
rect 27252 44693 27261 44727
rect 27261 44693 27295 44727
rect 27295 44693 27304 44727
rect 27252 44684 27304 44693
rect 29092 44727 29144 44736
rect 29092 44693 29101 44727
rect 29101 44693 29135 44727
rect 29135 44693 29144 44727
rect 29092 44684 29144 44693
rect 32036 44727 32088 44736
rect 32036 44693 32045 44727
rect 32045 44693 32079 44727
rect 32079 44693 32088 44727
rect 32036 44684 32088 44693
rect 57336 44684 57388 44736
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 17592 44480 17644 44532
rect 19340 44480 19392 44532
rect 20904 44480 20956 44532
rect 23940 44523 23992 44532
rect 23940 44489 23949 44523
rect 23949 44489 23983 44523
rect 23983 44489 23992 44523
rect 23940 44480 23992 44489
rect 24308 44480 24360 44532
rect 28448 44523 28500 44532
rect 28448 44489 28457 44523
rect 28457 44489 28491 44523
rect 28491 44489 28500 44523
rect 28448 44480 28500 44489
rect 31944 44523 31996 44532
rect 31944 44489 31953 44523
rect 31953 44489 31987 44523
rect 31987 44489 31996 44523
rect 31944 44480 31996 44489
rect 32128 44523 32180 44532
rect 32128 44489 32137 44523
rect 32137 44489 32171 44523
rect 32171 44489 32180 44523
rect 32128 44480 32180 44489
rect 57980 44523 58032 44532
rect 57980 44489 57989 44523
rect 57989 44489 58023 44523
rect 58023 44489 58032 44523
rect 57980 44480 58032 44489
rect 28264 44455 28316 44464
rect 28264 44421 28273 44455
rect 28273 44421 28307 44455
rect 28307 44421 28316 44455
rect 28264 44412 28316 44421
rect 18144 44276 18196 44328
rect 23848 44344 23900 44396
rect 20352 44319 20404 44328
rect 20352 44285 20361 44319
rect 20361 44285 20395 44319
rect 20395 44285 20404 44319
rect 20352 44276 20404 44285
rect 20996 44319 21048 44328
rect 20996 44285 21005 44319
rect 21005 44285 21039 44319
rect 21039 44285 21048 44319
rect 20996 44276 21048 44285
rect 21640 44276 21692 44328
rect 22560 44319 22612 44328
rect 22560 44285 22569 44319
rect 22569 44285 22603 44319
rect 22603 44285 22612 44319
rect 22560 44276 22612 44285
rect 22652 44276 22704 44328
rect 29000 44344 29052 44396
rect 33048 44455 33100 44464
rect 33048 44421 33057 44455
rect 33057 44421 33091 44455
rect 33091 44421 33100 44455
rect 33048 44412 33100 44421
rect 17960 44208 18012 44260
rect 26332 44276 26384 44328
rect 27252 44276 27304 44328
rect 30564 44276 30616 44328
rect 32036 44276 32088 44328
rect 57336 44276 57388 44328
rect 25228 44208 25280 44260
rect 26700 44251 26752 44260
rect 26700 44217 26709 44251
rect 26709 44217 26743 44251
rect 26743 44217 26752 44251
rect 26700 44208 26752 44217
rect 28080 44208 28132 44260
rect 29368 44208 29420 44260
rect 32220 44208 32272 44260
rect 30472 44140 30524 44192
rect 31944 44183 31996 44192
rect 31944 44149 31974 44183
rect 31974 44149 31996 44183
rect 31944 44140 31996 44149
rect 32312 44140 32364 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 24216 43936 24268 43988
rect 25136 43936 25188 43988
rect 26240 43936 26292 43988
rect 21088 43911 21140 43920
rect 21088 43877 21097 43911
rect 21097 43877 21131 43911
rect 21131 43877 21140 43911
rect 21088 43868 21140 43877
rect 21180 43868 21232 43920
rect 1400 43843 1452 43852
rect 1400 43809 1409 43843
rect 1409 43809 1443 43843
rect 1443 43809 1452 43843
rect 1400 43800 1452 43809
rect 20904 43732 20956 43784
rect 23388 43800 23440 43852
rect 25320 43800 25372 43852
rect 26332 43843 26384 43852
rect 26332 43809 26341 43843
rect 26341 43809 26375 43843
rect 26375 43809 26384 43843
rect 26332 43800 26384 43809
rect 27896 43800 27948 43852
rect 28080 43843 28132 43852
rect 28080 43809 28089 43843
rect 28089 43809 28123 43843
rect 28123 43809 28132 43843
rect 28080 43800 28132 43809
rect 28264 43800 28316 43852
rect 29000 43868 29052 43920
rect 31944 43936 31996 43988
rect 33968 43979 34020 43988
rect 33968 43945 33977 43979
rect 33977 43945 34011 43979
rect 34011 43945 34020 43979
rect 33968 43936 34020 43945
rect 29092 43800 29144 43852
rect 30472 43843 30524 43852
rect 26700 43732 26752 43784
rect 27528 43732 27580 43784
rect 30472 43809 30481 43843
rect 30481 43809 30515 43843
rect 30515 43809 30524 43843
rect 30472 43800 30524 43809
rect 32220 43868 32272 43920
rect 33048 43868 33100 43920
rect 58164 43911 58216 43920
rect 58164 43877 58173 43911
rect 58173 43877 58207 43911
rect 58207 43877 58216 43911
rect 58164 43868 58216 43877
rect 22744 43664 22796 43716
rect 26332 43664 26384 43716
rect 28080 43664 28132 43716
rect 28908 43664 28960 43716
rect 30564 43732 30616 43784
rect 31668 43732 31720 43784
rect 54944 43800 54996 43852
rect 32220 43732 32272 43784
rect 29368 43664 29420 43716
rect 20444 43639 20496 43648
rect 20444 43605 20453 43639
rect 20453 43605 20487 43639
rect 20487 43605 20496 43639
rect 20444 43596 20496 43605
rect 21364 43596 21416 43648
rect 31392 43639 31444 43648
rect 31392 43605 31401 43639
rect 31401 43605 31435 43639
rect 31435 43605 31444 43639
rect 31392 43596 31444 43605
rect 31944 43639 31996 43648
rect 31944 43605 31953 43639
rect 31953 43605 31987 43639
rect 31987 43605 31996 43639
rect 31944 43596 31996 43605
rect 32864 43596 32916 43648
rect 57428 43639 57480 43648
rect 57428 43605 57437 43639
rect 57437 43605 57471 43639
rect 57471 43605 57480 43639
rect 57428 43596 57480 43605
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 26332 43435 26384 43444
rect 26332 43401 26341 43435
rect 26341 43401 26375 43435
rect 26375 43401 26384 43435
rect 26332 43392 26384 43401
rect 32220 43392 32272 43444
rect 22744 43324 22796 43376
rect 23664 43324 23716 43376
rect 30564 43324 30616 43376
rect 58164 43367 58216 43376
rect 58164 43333 58173 43367
rect 58173 43333 58207 43367
rect 58207 43333 58216 43367
rect 58164 43324 58216 43333
rect 20168 43231 20220 43240
rect 20168 43197 20177 43231
rect 20177 43197 20211 43231
rect 20211 43197 20220 43231
rect 20168 43188 20220 43197
rect 20444 43231 20496 43240
rect 20444 43197 20478 43231
rect 20478 43197 20496 43231
rect 20444 43188 20496 43197
rect 23388 43188 23440 43240
rect 22652 43120 22704 43172
rect 24308 43120 24360 43172
rect 26240 43188 26292 43240
rect 26700 43188 26752 43240
rect 27160 43188 27212 43240
rect 27804 43231 27856 43240
rect 27804 43197 27813 43231
rect 27813 43197 27847 43231
rect 27847 43197 27856 43231
rect 27804 43188 27856 43197
rect 28908 43188 28960 43240
rect 30564 43188 30616 43240
rect 31392 43188 31444 43240
rect 56508 43188 56560 43240
rect 57336 43188 57388 43240
rect 26608 43120 26660 43172
rect 27988 43120 28040 43172
rect 29736 43120 29788 43172
rect 57980 43163 58032 43172
rect 57980 43129 57989 43163
rect 57989 43129 58023 43163
rect 58023 43129 58032 43163
rect 57980 43120 58032 43129
rect 21364 43052 21416 43104
rect 22560 43095 22612 43104
rect 22560 43061 22569 43095
rect 22569 43061 22603 43095
rect 22603 43061 22612 43095
rect 22560 43052 22612 43061
rect 22744 43095 22796 43104
rect 22744 43061 22753 43095
rect 22753 43061 22787 43095
rect 22787 43061 22796 43095
rect 22744 43052 22796 43061
rect 25136 43095 25188 43104
rect 25136 43061 25145 43095
rect 25145 43061 25179 43095
rect 25179 43061 25188 43095
rect 25136 43052 25188 43061
rect 25872 43095 25924 43104
rect 25872 43061 25881 43095
rect 25881 43061 25915 43095
rect 25915 43061 25924 43095
rect 25872 43052 25924 43061
rect 27896 43052 27948 43104
rect 57704 43052 57756 43104
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 21180 42848 21232 42900
rect 22560 42780 22612 42832
rect 23664 42848 23716 42900
rect 23848 42848 23900 42900
rect 26608 42891 26660 42900
rect 26608 42857 26617 42891
rect 26617 42857 26651 42891
rect 26651 42857 26660 42891
rect 26608 42848 26660 42857
rect 27160 42891 27212 42900
rect 27160 42857 27169 42891
rect 27169 42857 27203 42891
rect 27203 42857 27212 42891
rect 27160 42848 27212 42857
rect 27988 42891 28040 42900
rect 27988 42857 27997 42891
rect 27997 42857 28031 42891
rect 28031 42857 28040 42891
rect 27988 42848 28040 42857
rect 57980 42848 58032 42900
rect 23388 42780 23440 42832
rect 25872 42780 25924 42832
rect 1400 42755 1452 42764
rect 1400 42721 1409 42755
rect 1409 42721 1443 42755
rect 1443 42721 1452 42755
rect 1400 42712 1452 42721
rect 21088 42712 21140 42764
rect 22652 42712 22704 42764
rect 25228 42755 25280 42764
rect 25228 42721 25237 42755
rect 25237 42721 25271 42755
rect 25271 42721 25280 42755
rect 25228 42712 25280 42721
rect 27528 42712 27580 42764
rect 29092 42712 29144 42764
rect 21180 42644 21232 42696
rect 27896 42644 27948 42696
rect 29552 42712 29604 42764
rect 30472 42755 30524 42764
rect 30472 42721 30481 42755
rect 30481 42721 30515 42755
rect 30515 42721 30524 42755
rect 30472 42712 30524 42721
rect 30656 42712 30708 42764
rect 20260 42551 20312 42560
rect 20260 42517 20269 42551
rect 20269 42517 20303 42551
rect 20303 42517 20312 42551
rect 20260 42508 20312 42517
rect 23572 42508 23624 42560
rect 25136 42576 25188 42628
rect 24492 42508 24544 42560
rect 28448 42508 28500 42560
rect 32864 42712 32916 42764
rect 56876 42755 56928 42764
rect 56876 42721 56885 42755
rect 56885 42721 56919 42755
rect 56919 42721 56928 42755
rect 56876 42712 56928 42721
rect 57060 42755 57112 42764
rect 57060 42721 57069 42755
rect 57069 42721 57103 42755
rect 57103 42721 57112 42755
rect 57060 42712 57112 42721
rect 57428 42712 57480 42764
rect 57704 42755 57756 42764
rect 57704 42721 57713 42755
rect 57713 42721 57747 42755
rect 57747 42721 57756 42755
rect 57704 42712 57756 42721
rect 33232 42644 33284 42696
rect 30840 42508 30892 42560
rect 31116 42551 31168 42560
rect 31116 42517 31125 42551
rect 31125 42517 31159 42551
rect 31159 42517 31168 42551
rect 31116 42508 31168 42517
rect 31668 42508 31720 42560
rect 33140 42508 33192 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 20904 42304 20956 42356
rect 24308 42347 24360 42356
rect 24308 42313 24317 42347
rect 24317 42313 24351 42347
rect 24351 42313 24360 42347
rect 24308 42304 24360 42313
rect 24952 42304 25004 42356
rect 25228 42304 25280 42356
rect 26148 42304 26200 42356
rect 26240 42304 26292 42356
rect 28448 42304 28500 42356
rect 30472 42347 30524 42356
rect 30472 42313 30481 42347
rect 30481 42313 30515 42347
rect 30515 42313 30524 42347
rect 30472 42304 30524 42313
rect 21180 42168 21232 42220
rect 27804 42236 27856 42288
rect 28172 42279 28224 42288
rect 28172 42245 28181 42279
rect 28181 42245 28215 42279
rect 28215 42245 28224 42279
rect 28172 42236 28224 42245
rect 30932 42236 30984 42288
rect 31668 42236 31720 42288
rect 1400 42143 1452 42152
rect 1400 42109 1409 42143
rect 1409 42109 1443 42143
rect 1443 42109 1452 42143
rect 1400 42100 1452 42109
rect 20260 42100 20312 42152
rect 21364 42143 21416 42152
rect 21364 42109 21373 42143
rect 21373 42109 21407 42143
rect 21407 42109 21416 42143
rect 21364 42100 21416 42109
rect 23388 42100 23440 42152
rect 23848 42143 23900 42152
rect 23848 42109 23857 42143
rect 23857 42109 23891 42143
rect 23891 42109 23900 42143
rect 28448 42168 28500 42220
rect 23848 42100 23900 42109
rect 24492 42143 24544 42152
rect 24492 42109 24501 42143
rect 24501 42109 24535 42143
rect 24535 42109 24544 42143
rect 24492 42100 24544 42109
rect 24584 42100 24636 42152
rect 20168 42032 20220 42084
rect 20720 42032 20772 42084
rect 23572 42075 23624 42084
rect 23572 42041 23581 42075
rect 23581 42041 23615 42075
rect 23615 42041 23624 42075
rect 23572 42032 23624 42041
rect 21088 41964 21140 42016
rect 25688 41964 25740 42016
rect 26332 42100 26384 42152
rect 28080 42100 28132 42152
rect 28816 42100 28868 42152
rect 29736 42100 29788 42152
rect 27896 42075 27948 42084
rect 27896 42041 27905 42075
rect 27905 42041 27939 42075
rect 27939 42041 27948 42075
rect 27896 42032 27948 42041
rect 31116 42032 31168 42084
rect 31484 42007 31536 42016
rect 31484 41973 31493 42007
rect 31493 41973 31527 42007
rect 31527 41973 31536 42007
rect 31484 41964 31536 41973
rect 32680 42168 32732 42220
rect 32128 42143 32180 42152
rect 32128 42109 32137 42143
rect 32137 42109 32171 42143
rect 32171 42109 32180 42143
rect 32128 42100 32180 42109
rect 33140 42100 33192 42152
rect 56508 42100 56560 42152
rect 57520 42100 57572 42152
rect 57980 42075 58032 42084
rect 57980 42041 57989 42075
rect 57989 42041 58023 42075
rect 58023 42041 58032 42075
rect 57980 42032 58032 42041
rect 58164 42075 58216 42084
rect 58164 42041 58173 42075
rect 58173 42041 58207 42075
rect 58207 42041 58216 42075
rect 58164 42032 58216 42041
rect 33324 41964 33376 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 21180 41760 21232 41812
rect 20812 41667 20864 41676
rect 20812 41633 20821 41667
rect 20821 41633 20855 41667
rect 20855 41633 20864 41667
rect 20812 41624 20864 41633
rect 21180 41624 21232 41676
rect 24216 41692 24268 41744
rect 24584 41692 24636 41744
rect 27804 41760 27856 41812
rect 28816 41760 28868 41812
rect 24032 41667 24084 41676
rect 24032 41633 24041 41667
rect 24041 41633 24075 41667
rect 24075 41633 24084 41667
rect 24032 41624 24084 41633
rect 24492 41624 24544 41676
rect 25504 41667 25556 41676
rect 25504 41633 25513 41667
rect 25513 41633 25547 41667
rect 25547 41633 25556 41667
rect 25504 41624 25556 41633
rect 25688 41667 25740 41676
rect 25688 41633 25697 41667
rect 25697 41633 25731 41667
rect 25731 41633 25740 41667
rect 25688 41624 25740 41633
rect 26148 41624 26200 41676
rect 27804 41624 27856 41676
rect 27896 41624 27948 41676
rect 28080 41624 28132 41676
rect 28448 41667 28500 41676
rect 28448 41633 28457 41667
rect 28457 41633 28491 41667
rect 28491 41633 28500 41667
rect 28448 41624 28500 41633
rect 20720 41556 20772 41608
rect 24124 41599 24176 41608
rect 24124 41565 24133 41599
rect 24133 41565 24167 41599
rect 24167 41565 24176 41599
rect 24124 41556 24176 41565
rect 25872 41556 25924 41608
rect 28908 41599 28960 41608
rect 28908 41565 28917 41599
rect 28917 41565 28951 41599
rect 28951 41565 28960 41599
rect 28908 41556 28960 41565
rect 32128 41760 32180 41812
rect 31484 41692 31536 41744
rect 57980 41760 58032 41812
rect 32680 41735 32732 41744
rect 32680 41701 32710 41735
rect 32710 41701 32732 41735
rect 33324 41735 33376 41744
rect 32680 41692 32732 41701
rect 33324 41701 33333 41735
rect 33333 41701 33367 41735
rect 33367 41701 33376 41735
rect 33324 41692 33376 41701
rect 28172 41488 28224 41540
rect 22376 41420 22428 41472
rect 23664 41463 23716 41472
rect 23664 41429 23673 41463
rect 23673 41429 23707 41463
rect 23707 41429 23716 41463
rect 23664 41420 23716 41429
rect 25228 41420 25280 41472
rect 57060 41667 57112 41676
rect 33048 41556 33100 41608
rect 57060 41633 57069 41667
rect 57069 41633 57103 41667
rect 57103 41633 57112 41667
rect 57060 41624 57112 41633
rect 57336 41624 57388 41676
rect 57520 41667 57572 41676
rect 57520 41633 57529 41667
rect 57529 41633 57563 41667
rect 57563 41633 57572 41667
rect 57520 41624 57572 41633
rect 32864 41531 32916 41540
rect 32864 41497 32873 41531
rect 32873 41497 32907 41531
rect 32907 41497 32916 41531
rect 32864 41488 32916 41497
rect 33232 41488 33284 41540
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 21180 41259 21232 41268
rect 21180 41225 21189 41259
rect 21189 41225 21223 41259
rect 21223 41225 21232 41259
rect 21180 41216 21232 41225
rect 24124 41216 24176 41268
rect 25872 41216 25924 41268
rect 27804 41259 27856 41268
rect 27804 41225 27813 41259
rect 27813 41225 27847 41259
rect 27847 41225 27856 41259
rect 27804 41216 27856 41225
rect 30564 41216 30616 41268
rect 57336 41259 57388 41268
rect 57336 41225 57345 41259
rect 57345 41225 57379 41259
rect 57379 41225 57388 41259
rect 57336 41216 57388 41225
rect 22652 41080 22704 41132
rect 28816 41123 28868 41132
rect 28816 41089 28825 41123
rect 28825 41089 28859 41123
rect 28859 41089 28868 41123
rect 28816 41080 28868 41089
rect 29828 41080 29880 41132
rect 1400 41055 1452 41064
rect 1400 41021 1409 41055
rect 1409 41021 1443 41055
rect 1443 41021 1452 41055
rect 1400 41012 1452 41021
rect 20812 41012 20864 41064
rect 21548 41055 21600 41064
rect 21548 41021 21557 41055
rect 21557 41021 21591 41055
rect 21591 41021 21600 41055
rect 21548 41012 21600 41021
rect 22376 41012 22428 41064
rect 23664 41012 23716 41064
rect 24952 41055 25004 41064
rect 24952 41021 24961 41055
rect 24961 41021 24995 41055
rect 24995 41021 25004 41055
rect 24952 41012 25004 41021
rect 25228 41055 25280 41064
rect 25228 41021 25262 41055
rect 25262 41021 25280 41055
rect 25228 41012 25280 41021
rect 27620 41012 27672 41064
rect 28080 41055 28132 41064
rect 28080 41021 28089 41055
rect 28089 41021 28123 41055
rect 28123 41021 28132 41055
rect 28080 41012 28132 41021
rect 28908 41012 28960 41064
rect 30840 41055 30892 41064
rect 30840 41021 30849 41055
rect 30849 41021 30883 41055
rect 30883 41021 30892 41055
rect 30840 41012 30892 41021
rect 21732 40944 21784 40996
rect 25412 40944 25464 40996
rect 27804 40987 27856 40996
rect 27804 40953 27813 40987
rect 27813 40953 27847 40987
rect 27847 40953 27856 40987
rect 27804 40944 27856 40953
rect 27988 40987 28040 40996
rect 27988 40953 27997 40987
rect 27997 40953 28031 40987
rect 28031 40953 28040 40987
rect 27988 40944 28040 40953
rect 28448 40944 28500 40996
rect 29000 40944 29052 40996
rect 29552 40944 29604 40996
rect 31760 41012 31812 41064
rect 32588 41012 32640 41064
rect 33140 41012 33192 41064
rect 56508 41055 56560 41064
rect 56508 41021 56517 41055
rect 56517 41021 56551 41055
rect 56551 41021 56560 41055
rect 56508 41012 56560 41021
rect 57520 40944 57572 40996
rect 57980 40987 58032 40996
rect 57980 40953 57989 40987
rect 57989 40953 58023 40987
rect 58023 40953 58032 40987
rect 57980 40944 58032 40953
rect 58164 40987 58216 40996
rect 58164 40953 58173 40987
rect 58173 40953 58207 40987
rect 58207 40953 58216 40987
rect 58164 40944 58216 40953
rect 30196 40919 30248 40928
rect 30196 40885 30205 40919
rect 30205 40885 30239 40919
rect 30239 40885 30248 40919
rect 30196 40876 30248 40885
rect 31852 40876 31904 40928
rect 33140 40919 33192 40928
rect 33140 40885 33149 40919
rect 33149 40885 33183 40919
rect 33183 40885 33192 40919
rect 33140 40876 33192 40885
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 21548 40672 21600 40724
rect 20076 40647 20128 40656
rect 15200 40536 15252 40588
rect 15292 40579 15344 40588
rect 15292 40545 15301 40579
rect 15301 40545 15335 40579
rect 15335 40545 15344 40579
rect 20076 40613 20085 40647
rect 20085 40613 20119 40647
rect 20119 40613 20128 40647
rect 20076 40604 20128 40613
rect 15292 40536 15344 40545
rect 19984 40579 20036 40588
rect 19984 40545 19993 40579
rect 19993 40545 20027 40579
rect 20027 40545 20036 40579
rect 19984 40536 20036 40545
rect 19708 40468 19760 40520
rect 20904 40536 20956 40588
rect 21732 40672 21784 40724
rect 24216 40715 24268 40724
rect 24216 40681 24225 40715
rect 24225 40681 24259 40715
rect 24259 40681 24268 40715
rect 24216 40672 24268 40681
rect 29000 40715 29052 40724
rect 29000 40681 29009 40715
rect 29009 40681 29043 40715
rect 29043 40681 29052 40715
rect 29000 40672 29052 40681
rect 32588 40715 32640 40724
rect 32588 40681 32597 40715
rect 32597 40681 32631 40715
rect 32631 40681 32640 40715
rect 32588 40672 32640 40681
rect 57980 40672 58032 40724
rect 22376 40579 22428 40588
rect 22376 40545 22385 40579
rect 22385 40545 22419 40579
rect 22419 40545 22428 40579
rect 22376 40536 22428 40545
rect 24032 40579 24084 40588
rect 24032 40545 24041 40579
rect 24041 40545 24075 40579
rect 24075 40545 24084 40579
rect 24032 40536 24084 40545
rect 24124 40536 24176 40588
rect 25688 40579 25740 40588
rect 25688 40545 25697 40579
rect 25697 40545 25731 40579
rect 25731 40545 25740 40579
rect 25688 40536 25740 40545
rect 25872 40579 25924 40588
rect 25872 40545 25881 40579
rect 25881 40545 25915 40579
rect 25915 40545 25924 40579
rect 25872 40536 25924 40545
rect 27988 40604 28040 40656
rect 21088 40511 21140 40520
rect 21088 40477 21097 40511
rect 21097 40477 21131 40511
rect 21131 40477 21140 40511
rect 21088 40468 21140 40477
rect 28908 40536 28960 40588
rect 30196 40604 30248 40656
rect 29276 40579 29328 40588
rect 29276 40545 29285 40579
rect 29285 40545 29319 40579
rect 29319 40545 29328 40579
rect 29552 40579 29604 40588
rect 29276 40536 29328 40545
rect 29552 40545 29561 40579
rect 29561 40545 29595 40579
rect 29595 40545 29604 40579
rect 29552 40536 29604 40545
rect 25504 40400 25556 40452
rect 27620 40468 27672 40520
rect 27988 40511 28040 40520
rect 27988 40477 27997 40511
rect 27997 40477 28031 40511
rect 28031 40477 28040 40511
rect 27988 40468 28040 40477
rect 31576 40579 31628 40588
rect 31576 40545 31585 40579
rect 31585 40545 31619 40579
rect 31619 40545 31628 40579
rect 31852 40579 31904 40588
rect 31576 40536 31628 40545
rect 31852 40545 31861 40579
rect 31861 40545 31895 40579
rect 31895 40545 31904 40579
rect 31852 40536 31904 40545
rect 34060 40604 34112 40656
rect 57060 40579 57112 40588
rect 31760 40468 31812 40520
rect 57060 40545 57069 40579
rect 57069 40545 57103 40579
rect 57103 40545 57112 40579
rect 57060 40536 57112 40545
rect 57428 40468 57480 40520
rect 27804 40400 27856 40452
rect 29828 40400 29880 40452
rect 15384 40332 15436 40384
rect 18604 40375 18656 40384
rect 18604 40341 18613 40375
rect 18613 40341 18647 40375
rect 18647 40341 18656 40375
rect 18604 40332 18656 40341
rect 20444 40332 20496 40384
rect 20812 40332 20864 40384
rect 27712 40332 27764 40384
rect 31300 40375 31352 40384
rect 31300 40341 31309 40375
rect 31309 40341 31343 40375
rect 31343 40341 31352 40375
rect 31300 40332 31352 40341
rect 31852 40332 31904 40384
rect 33876 40375 33928 40384
rect 33876 40341 33885 40375
rect 33885 40341 33919 40375
rect 33919 40341 33928 40375
rect 33876 40332 33928 40341
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 19708 40171 19760 40180
rect 19708 40137 19717 40171
rect 19717 40137 19751 40171
rect 19751 40137 19760 40171
rect 19708 40128 19760 40137
rect 21088 40128 21140 40180
rect 29276 40128 29328 40180
rect 31760 40128 31812 40180
rect 57428 40171 57480 40180
rect 57428 40137 57437 40171
rect 57437 40137 57471 40171
rect 57471 40137 57480 40171
rect 57428 40128 57480 40137
rect 1400 39967 1452 39976
rect 1400 39933 1409 39967
rect 1409 39933 1443 39967
rect 1443 39933 1452 39967
rect 1400 39924 1452 39933
rect 12624 39967 12676 39976
rect 12624 39933 12633 39967
rect 12633 39933 12667 39967
rect 12667 39933 12676 39967
rect 12624 39924 12676 39933
rect 13268 39924 13320 39976
rect 15752 40060 15804 40112
rect 34060 39992 34112 40044
rect 13452 39856 13504 39908
rect 12256 39831 12308 39840
rect 12256 39797 12265 39831
rect 12265 39797 12299 39831
rect 12299 39797 12308 39831
rect 12256 39788 12308 39797
rect 13728 39788 13780 39840
rect 14004 39788 14056 39840
rect 16764 39924 16816 39976
rect 17684 39924 17736 39976
rect 18604 39967 18656 39976
rect 18604 39933 18638 39967
rect 18638 39933 18656 39967
rect 18604 39924 18656 39933
rect 20444 39967 20496 39976
rect 20444 39933 20478 39967
rect 20478 39933 20496 39967
rect 20444 39924 20496 39933
rect 25964 39967 26016 39976
rect 25964 39933 25973 39967
rect 25973 39933 26007 39967
rect 26007 39933 26016 39967
rect 25964 39924 26016 39933
rect 20720 39856 20772 39908
rect 27712 39856 27764 39908
rect 29828 39924 29880 39976
rect 31300 39924 31352 39976
rect 30932 39856 30984 39908
rect 33140 39924 33192 39976
rect 33416 39856 33468 39908
rect 15476 39788 15528 39840
rect 26056 39831 26108 39840
rect 26056 39797 26065 39831
rect 26065 39797 26099 39831
rect 26099 39797 26108 39831
rect 26056 39788 26108 39797
rect 27896 39788 27948 39840
rect 58624 39924 58676 39976
rect 58164 39899 58216 39908
rect 58164 39865 58173 39899
rect 58173 39865 58207 39899
rect 58207 39865 58216 39899
rect 58164 39856 58216 39865
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 12624 39584 12676 39636
rect 13452 39627 13504 39636
rect 12256 39516 12308 39568
rect 13452 39593 13461 39627
rect 13461 39593 13495 39627
rect 13495 39593 13504 39627
rect 13452 39584 13504 39593
rect 16764 39584 16816 39636
rect 20904 39627 20956 39636
rect 20904 39593 20913 39627
rect 20913 39593 20947 39627
rect 20947 39593 20956 39627
rect 20904 39584 20956 39593
rect 25964 39584 26016 39636
rect 28172 39627 28224 39636
rect 28172 39593 28181 39627
rect 28181 39593 28215 39627
rect 28215 39593 28224 39627
rect 28172 39584 28224 39593
rect 31576 39584 31628 39636
rect 33048 39627 33100 39636
rect 33048 39593 33057 39627
rect 33057 39593 33091 39627
rect 33091 39593 33100 39627
rect 33048 39584 33100 39593
rect 15384 39516 15436 39568
rect 26056 39516 26108 39568
rect 13268 39380 13320 39432
rect 18052 39448 18104 39500
rect 20076 39448 20128 39500
rect 20812 39491 20864 39500
rect 20812 39457 20821 39491
rect 20821 39457 20855 39491
rect 20855 39457 20864 39491
rect 20812 39448 20864 39457
rect 21088 39448 21140 39500
rect 27344 39491 27396 39500
rect 27344 39457 27353 39491
rect 27353 39457 27387 39491
rect 27387 39457 27396 39491
rect 27344 39448 27396 39457
rect 27988 39448 28040 39500
rect 31760 39448 31812 39500
rect 32128 39448 32180 39500
rect 13728 39380 13780 39432
rect 25504 39423 25556 39432
rect 25504 39389 25513 39423
rect 25513 39389 25547 39423
rect 25547 39389 25556 39423
rect 25504 39380 25556 39389
rect 32864 39380 32916 39432
rect 15568 39244 15620 39296
rect 28540 39244 28592 39296
rect 33876 39516 33928 39568
rect 57980 39491 58032 39500
rect 57980 39457 57989 39491
rect 57989 39457 58023 39491
rect 58023 39457 58032 39491
rect 57980 39448 58032 39457
rect 33048 39312 33100 39364
rect 33232 39244 33284 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 1400 38879 1452 38888
rect 1400 38845 1409 38879
rect 1409 38845 1443 38879
rect 1443 38845 1452 38879
rect 1400 38836 1452 38845
rect 13268 38836 13320 38888
rect 13452 38836 13504 38888
rect 12532 38743 12584 38752
rect 12532 38709 12541 38743
rect 12541 38709 12575 38743
rect 12575 38709 12584 38743
rect 12532 38700 12584 38709
rect 15200 39040 15252 39092
rect 19984 39040 20036 39092
rect 15292 38972 15344 39024
rect 25872 39015 25924 39024
rect 25872 38981 25881 39015
rect 25881 38981 25915 39015
rect 25915 38981 25924 39015
rect 25872 38972 25924 38981
rect 33692 38972 33744 39024
rect 17684 38947 17736 38956
rect 17684 38913 17693 38947
rect 17693 38913 17727 38947
rect 17727 38913 17736 38947
rect 17684 38904 17736 38913
rect 25964 38904 26016 38956
rect 32128 38947 32180 38956
rect 32128 38913 32137 38947
rect 32137 38913 32171 38947
rect 32171 38913 32180 38947
rect 32128 38904 32180 38913
rect 15568 38879 15620 38888
rect 15568 38845 15577 38879
rect 15577 38845 15611 38879
rect 15611 38845 15620 38879
rect 15568 38836 15620 38845
rect 15752 38879 15804 38888
rect 15752 38845 15761 38879
rect 15761 38845 15795 38879
rect 15795 38845 15804 38879
rect 15752 38836 15804 38845
rect 19892 38879 19944 38888
rect 15476 38700 15528 38752
rect 18972 38768 19024 38820
rect 19892 38845 19901 38879
rect 19901 38845 19935 38879
rect 19935 38845 19944 38879
rect 19892 38836 19944 38845
rect 19984 38879 20036 38888
rect 19984 38845 19993 38879
rect 19993 38845 20027 38879
rect 20027 38845 20036 38879
rect 20444 38879 20496 38888
rect 19984 38836 20036 38845
rect 20444 38845 20453 38879
rect 20453 38845 20487 38879
rect 20487 38845 20496 38879
rect 20444 38836 20496 38845
rect 20720 38836 20772 38888
rect 26516 38879 26568 38888
rect 26516 38845 26525 38879
rect 26525 38845 26559 38879
rect 26559 38845 26568 38879
rect 26516 38836 26568 38845
rect 27344 38836 27396 38888
rect 30932 38836 30984 38888
rect 31760 38836 31812 38888
rect 32404 38836 32456 38888
rect 33048 38879 33100 38888
rect 33048 38845 33057 38879
rect 33057 38845 33091 38879
rect 33091 38845 33100 38879
rect 33048 38836 33100 38845
rect 33232 38879 33284 38888
rect 33232 38845 33241 38879
rect 33241 38845 33275 38879
rect 33275 38845 33284 38879
rect 33232 38836 33284 38845
rect 33416 38836 33468 38888
rect 28816 38768 28868 38820
rect 33968 38811 34020 38820
rect 33968 38777 34002 38811
rect 34002 38777 34020 38811
rect 57980 38811 58032 38820
rect 33968 38768 34020 38777
rect 57980 38777 57989 38811
rect 57989 38777 58023 38811
rect 58023 38777 58032 38811
rect 57980 38768 58032 38777
rect 58164 38811 58216 38820
rect 58164 38777 58173 38811
rect 58173 38777 58207 38811
rect 58207 38777 58216 38811
rect 58164 38768 58216 38777
rect 18236 38700 18288 38752
rect 20168 38700 20220 38752
rect 29184 38700 29236 38752
rect 31668 38743 31720 38752
rect 31668 38709 31677 38743
rect 31677 38709 31711 38743
rect 31711 38709 31720 38743
rect 31668 38700 31720 38709
rect 35256 38700 35308 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 13268 38539 13320 38548
rect 13268 38505 13277 38539
rect 13277 38505 13311 38539
rect 13311 38505 13320 38539
rect 13268 38496 13320 38505
rect 18972 38539 19024 38548
rect 12532 38428 12584 38480
rect 1400 38403 1452 38412
rect 1400 38369 1409 38403
rect 1409 38369 1443 38403
rect 1443 38369 1452 38403
rect 1400 38360 1452 38369
rect 13728 38360 13780 38412
rect 15660 38360 15712 38412
rect 16764 38428 16816 38480
rect 17960 38428 18012 38480
rect 18972 38505 18981 38539
rect 18981 38505 19015 38539
rect 19015 38505 19024 38539
rect 18972 38496 19024 38505
rect 19984 38496 20036 38548
rect 26516 38496 26568 38548
rect 18696 38428 18748 38480
rect 20168 38428 20220 38480
rect 32128 38496 32180 38548
rect 32404 38496 32456 38548
rect 57980 38496 58032 38548
rect 28448 38428 28500 38480
rect 29184 38471 29236 38480
rect 29184 38437 29193 38471
rect 29193 38437 29227 38471
rect 29227 38437 29236 38471
rect 29184 38428 29236 38437
rect 31668 38428 31720 38480
rect 33692 38428 33744 38480
rect 17316 38360 17368 38412
rect 18880 38403 18932 38412
rect 18880 38369 18889 38403
rect 18889 38369 18923 38403
rect 18923 38369 18932 38403
rect 18880 38360 18932 38369
rect 15108 38292 15160 38344
rect 19892 38360 19944 38412
rect 20720 38360 20772 38412
rect 25872 38403 25924 38412
rect 25872 38369 25881 38403
rect 25881 38369 25915 38403
rect 25915 38369 25924 38403
rect 25872 38360 25924 38369
rect 25964 38360 26016 38412
rect 27804 38360 27856 38412
rect 30932 38403 30984 38412
rect 30932 38369 30941 38403
rect 30941 38369 30975 38403
rect 30975 38369 30984 38403
rect 30932 38360 30984 38369
rect 25504 38292 25556 38344
rect 28540 38292 28592 38344
rect 32864 38403 32916 38412
rect 32864 38369 32873 38403
rect 32873 38369 32907 38403
rect 32907 38369 32916 38403
rect 32864 38360 32916 38369
rect 33232 38360 33284 38412
rect 34152 38403 34204 38412
rect 34152 38369 34161 38403
rect 34161 38369 34195 38403
rect 34195 38369 34204 38403
rect 34152 38360 34204 38369
rect 57704 38335 57756 38344
rect 57704 38301 57713 38335
rect 57713 38301 57747 38335
rect 57747 38301 57756 38335
rect 57704 38292 57756 38301
rect 33048 38224 33100 38276
rect 33968 38267 34020 38276
rect 33968 38233 33977 38267
rect 33977 38233 34011 38267
rect 34011 38233 34020 38267
rect 33968 38224 34020 38233
rect 14740 38199 14792 38208
rect 14740 38165 14749 38199
rect 14749 38165 14783 38199
rect 14783 38165 14792 38199
rect 14740 38156 14792 38165
rect 15292 38156 15344 38208
rect 18236 38199 18288 38208
rect 18236 38165 18245 38199
rect 18245 38165 18279 38199
rect 18279 38165 18288 38199
rect 18236 38156 18288 38165
rect 28540 38199 28592 38208
rect 28540 38165 28549 38199
rect 28549 38165 28583 38199
rect 28583 38165 28592 38199
rect 28540 38156 28592 38165
rect 28724 38199 28776 38208
rect 28724 38165 28733 38199
rect 28733 38165 28767 38199
rect 28767 38165 28776 38199
rect 28724 38156 28776 38165
rect 28908 38156 28960 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 15108 37995 15160 38004
rect 15108 37961 15117 37995
rect 15117 37961 15151 37995
rect 15151 37961 15160 37995
rect 15108 37952 15160 37961
rect 15660 37995 15712 38004
rect 15660 37961 15669 37995
rect 15669 37961 15703 37995
rect 15703 37961 15712 37995
rect 15660 37952 15712 37961
rect 17316 37995 17368 38004
rect 17316 37961 17325 37995
rect 17325 37961 17359 37995
rect 17359 37961 17368 37995
rect 17316 37952 17368 37961
rect 18880 37952 18932 38004
rect 27804 37995 27856 38004
rect 27804 37961 27813 37995
rect 27813 37961 27847 37995
rect 27847 37961 27856 37995
rect 27804 37952 27856 37961
rect 28540 37952 28592 38004
rect 28816 37952 28868 38004
rect 34152 37952 34204 38004
rect 57704 37952 57756 38004
rect 58164 37927 58216 37936
rect 17960 37859 18012 37868
rect 13728 37791 13780 37800
rect 13728 37757 13737 37791
rect 13737 37757 13771 37791
rect 13771 37757 13780 37791
rect 13728 37748 13780 37757
rect 14740 37748 14792 37800
rect 15292 37748 15344 37800
rect 16396 37791 16448 37800
rect 16396 37757 16405 37791
rect 16405 37757 16439 37791
rect 16439 37757 16448 37791
rect 16396 37748 16448 37757
rect 17960 37825 17969 37859
rect 17969 37825 18003 37859
rect 18003 37825 18012 37859
rect 17960 37816 18012 37825
rect 18236 37748 18288 37800
rect 58164 37893 58173 37927
rect 58173 37893 58207 37927
rect 58207 37893 58216 37927
rect 58164 37884 58216 37893
rect 20996 37816 21048 37868
rect 25320 37816 25372 37868
rect 28448 37859 28500 37868
rect 18696 37791 18748 37800
rect 18696 37757 18705 37791
rect 18705 37757 18739 37791
rect 18739 37757 18748 37791
rect 18696 37748 18748 37757
rect 28448 37825 28457 37859
rect 28457 37825 28491 37859
rect 28491 37825 28500 37859
rect 28448 37816 28500 37825
rect 28724 37816 28776 37868
rect 28908 37791 28960 37800
rect 28908 37757 28917 37791
rect 28917 37757 28951 37791
rect 28951 37757 28960 37791
rect 28908 37748 28960 37757
rect 33324 37791 33376 37800
rect 33324 37757 33333 37791
rect 33333 37757 33367 37791
rect 33367 37757 33376 37791
rect 33324 37748 33376 37757
rect 34796 37748 34848 37800
rect 35256 37748 35308 37800
rect 56508 37748 56560 37800
rect 57428 37791 57480 37800
rect 57428 37757 57437 37791
rect 57437 37757 57471 37791
rect 57471 37757 57480 37791
rect 57428 37748 57480 37757
rect 1308 37680 1360 37732
rect 33048 37680 33100 37732
rect 33508 37723 33560 37732
rect 33508 37689 33517 37723
rect 33517 37689 33551 37723
rect 33551 37689 33560 37723
rect 33508 37680 33560 37689
rect 58716 37680 58768 37732
rect 16212 37655 16264 37664
rect 16212 37621 16221 37655
rect 16221 37621 16255 37655
rect 16255 37621 16264 37655
rect 16212 37612 16264 37621
rect 18696 37612 18748 37664
rect 20996 37655 21048 37664
rect 20996 37621 21005 37655
rect 21005 37621 21039 37655
rect 21039 37621 21048 37655
rect 20996 37612 21048 37621
rect 28540 37612 28592 37664
rect 34520 37655 34572 37664
rect 34520 37621 34529 37655
rect 34529 37621 34563 37655
rect 34563 37621 34572 37655
rect 34520 37612 34572 37621
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 16396 37408 16448 37460
rect 17960 37408 18012 37460
rect 18696 37408 18748 37460
rect 20444 37408 20496 37460
rect 20720 37408 20772 37460
rect 34796 37451 34848 37460
rect 34796 37417 34805 37451
rect 34805 37417 34839 37451
rect 34839 37417 34848 37451
rect 34796 37408 34848 37417
rect 57888 37408 57940 37460
rect 15752 37383 15804 37392
rect 1400 37315 1452 37324
rect 1400 37281 1409 37315
rect 1409 37281 1443 37315
rect 1443 37281 1452 37315
rect 1400 37272 1452 37281
rect 15752 37349 15761 37383
rect 15761 37349 15795 37383
rect 15795 37349 15804 37383
rect 15752 37340 15804 37349
rect 18604 37340 18656 37392
rect 15660 37315 15712 37324
rect 15660 37281 15669 37315
rect 15669 37281 15703 37315
rect 15703 37281 15712 37315
rect 15660 37272 15712 37281
rect 15200 37247 15252 37256
rect 15200 37213 15209 37247
rect 15209 37213 15243 37247
rect 15243 37213 15252 37247
rect 15200 37204 15252 37213
rect 16948 37315 17000 37324
rect 16948 37281 16957 37315
rect 16957 37281 16991 37315
rect 16991 37281 17000 37315
rect 16948 37272 17000 37281
rect 17132 37315 17184 37324
rect 17132 37281 17141 37315
rect 17141 37281 17175 37315
rect 17175 37281 17184 37315
rect 17132 37272 17184 37281
rect 18052 37315 18104 37324
rect 18052 37281 18061 37315
rect 18061 37281 18095 37315
rect 18095 37281 18104 37315
rect 18052 37272 18104 37281
rect 18236 37315 18288 37324
rect 18236 37281 18245 37315
rect 18245 37281 18279 37315
rect 18279 37281 18288 37315
rect 18236 37272 18288 37281
rect 28080 37340 28132 37392
rect 19892 37272 19944 37324
rect 20076 37272 20128 37324
rect 20720 37272 20772 37324
rect 28264 37204 28316 37256
rect 28632 37272 28684 37324
rect 30472 37315 30524 37324
rect 30472 37281 30481 37315
rect 30481 37281 30515 37315
rect 30515 37281 30524 37315
rect 30472 37272 30524 37281
rect 30656 37315 30708 37324
rect 30656 37281 30665 37315
rect 30665 37281 30699 37315
rect 30699 37281 30708 37315
rect 30656 37272 30708 37281
rect 30932 37272 30984 37324
rect 33508 37340 33560 37392
rect 32220 37272 32272 37324
rect 33140 37272 33192 37324
rect 33416 37315 33468 37324
rect 33416 37281 33425 37315
rect 33425 37281 33459 37315
rect 33459 37281 33468 37315
rect 33416 37272 33468 37281
rect 56784 37272 56836 37324
rect 56968 37272 57020 37324
rect 57980 37315 58032 37324
rect 57980 37281 57989 37315
rect 57989 37281 58023 37315
rect 58023 37281 58032 37315
rect 57980 37272 58032 37281
rect 28724 37204 28776 37256
rect 15844 37136 15896 37188
rect 14740 37111 14792 37120
rect 14740 37077 14749 37111
rect 14749 37077 14783 37111
rect 14783 37077 14792 37111
rect 14740 37068 14792 37077
rect 17684 37068 17736 37120
rect 30564 37111 30616 37120
rect 30564 37077 30573 37111
rect 30573 37077 30607 37111
rect 30607 37077 30616 37111
rect 30564 37068 30616 37077
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 57428 37111 57480 37120
rect 57428 37077 57437 37111
rect 57437 37077 57471 37111
rect 57471 37077 57480 37111
rect 57428 37068 57480 37077
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 15200 36864 15252 36916
rect 15844 36907 15896 36916
rect 15844 36873 15853 36907
rect 15853 36873 15887 36907
rect 15887 36873 15896 36907
rect 15844 36864 15896 36873
rect 18236 36864 18288 36916
rect 18880 36864 18932 36916
rect 28264 36907 28316 36916
rect 28264 36873 28273 36907
rect 28273 36873 28307 36907
rect 28307 36873 28316 36907
rect 28264 36864 28316 36873
rect 30472 36864 30524 36916
rect 57980 36907 58032 36916
rect 57980 36873 57989 36907
rect 57989 36873 58023 36907
rect 58023 36873 58032 36907
rect 57980 36864 58032 36873
rect 30656 36796 30708 36848
rect 17592 36771 17644 36780
rect 13728 36660 13780 36712
rect 14740 36660 14792 36712
rect 15752 36703 15804 36712
rect 15752 36669 15761 36703
rect 15761 36669 15795 36703
rect 15795 36669 15804 36703
rect 15752 36660 15804 36669
rect 17592 36737 17601 36771
rect 17601 36737 17635 36771
rect 17635 36737 17644 36771
rect 17592 36728 17644 36737
rect 28080 36703 28132 36712
rect 28080 36669 28089 36703
rect 28089 36669 28123 36703
rect 28123 36669 28132 36703
rect 28080 36660 28132 36669
rect 28632 36660 28684 36712
rect 30932 36728 30984 36780
rect 34520 36796 34572 36848
rect 30564 36660 30616 36712
rect 32496 36660 32548 36712
rect 33784 36728 33836 36780
rect 57704 36703 57756 36712
rect 16212 36592 16264 36644
rect 18420 36592 18472 36644
rect 57704 36669 57713 36703
rect 57713 36669 57747 36703
rect 57747 36669 57756 36703
rect 57704 36660 57756 36669
rect 57060 36635 57112 36644
rect 27896 36567 27948 36576
rect 27896 36533 27905 36567
rect 27905 36533 27939 36567
rect 27939 36533 27948 36567
rect 27896 36524 27948 36533
rect 32772 36524 32824 36576
rect 33048 36524 33100 36576
rect 57060 36601 57069 36635
rect 57069 36601 57103 36635
rect 57103 36601 57112 36635
rect 57060 36592 57112 36601
rect 56968 36524 57020 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 17132 36320 17184 36372
rect 18420 36363 18472 36372
rect 18420 36329 18429 36363
rect 18429 36329 18463 36363
rect 18463 36329 18472 36363
rect 18420 36320 18472 36329
rect 28632 36363 28684 36372
rect 28632 36329 28641 36363
rect 28641 36329 28675 36363
rect 28675 36329 28684 36363
rect 28632 36320 28684 36329
rect 32220 36363 32272 36372
rect 32220 36329 32229 36363
rect 32229 36329 32263 36363
rect 32263 36329 32272 36363
rect 32220 36320 32272 36329
rect 33324 36320 33376 36372
rect 57704 36320 57756 36372
rect 1400 36227 1452 36236
rect 1400 36193 1409 36227
rect 1409 36193 1443 36227
rect 1443 36193 1452 36227
rect 1400 36184 1452 36193
rect 16212 36252 16264 36304
rect 17684 36227 17736 36236
rect 17684 36193 17693 36227
rect 17693 36193 17727 36227
rect 17727 36193 17736 36227
rect 17684 36184 17736 36193
rect 27896 36252 27948 36304
rect 18604 36227 18656 36236
rect 18604 36193 18613 36227
rect 18613 36193 18647 36227
rect 18647 36193 18656 36227
rect 18604 36184 18656 36193
rect 18880 36227 18932 36236
rect 18880 36193 18889 36227
rect 18889 36193 18923 36227
rect 18923 36193 18932 36227
rect 18880 36184 18932 36193
rect 30564 36184 30616 36236
rect 32404 36227 32456 36236
rect 32404 36193 32413 36227
rect 32413 36193 32447 36227
rect 32447 36193 32456 36227
rect 32404 36184 32456 36193
rect 32772 36227 32824 36236
rect 16948 36116 17000 36168
rect 27252 36159 27304 36168
rect 27252 36125 27261 36159
rect 27261 36125 27295 36159
rect 27295 36125 27304 36159
rect 27252 36116 27304 36125
rect 32772 36193 32781 36227
rect 32781 36193 32815 36227
rect 32815 36193 32824 36227
rect 32772 36184 32824 36193
rect 34520 36252 34572 36304
rect 33784 36184 33836 36236
rect 57428 36227 57480 36236
rect 57428 36193 57437 36227
rect 57437 36193 57471 36227
rect 57471 36193 57480 36227
rect 57428 36184 57480 36193
rect 57980 36227 58032 36236
rect 57980 36193 57989 36227
rect 57989 36193 58023 36227
rect 58023 36193 58032 36227
rect 57980 36184 58032 36193
rect 34244 36091 34296 36100
rect 34244 36057 34253 36091
rect 34253 36057 34287 36091
rect 34287 36057 34296 36091
rect 34244 36048 34296 36057
rect 18788 36023 18840 36032
rect 18788 35989 18797 36023
rect 18797 35989 18831 36023
rect 18831 35989 18840 36023
rect 18788 35980 18840 35989
rect 31116 35980 31168 36032
rect 33692 35980 33744 36032
rect 57888 35980 57940 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 18052 35776 18104 35828
rect 18788 35776 18840 35828
rect 31116 35819 31168 35828
rect 31116 35785 31125 35819
rect 31125 35785 31159 35819
rect 31159 35785 31168 35819
rect 31116 35776 31168 35785
rect 57980 35819 58032 35828
rect 57980 35785 57989 35819
rect 57989 35785 58023 35819
rect 58023 35785 58032 35819
rect 57980 35776 58032 35785
rect 17960 35708 18012 35760
rect 33140 35683 33192 35692
rect 1400 35615 1452 35624
rect 1400 35581 1409 35615
rect 1409 35581 1443 35615
rect 1443 35581 1452 35615
rect 1400 35572 1452 35581
rect 17684 35572 17736 35624
rect 18328 35615 18380 35624
rect 18328 35581 18337 35615
rect 18337 35581 18371 35615
rect 18371 35581 18380 35615
rect 18328 35572 18380 35581
rect 33140 35649 33149 35683
rect 33149 35649 33183 35683
rect 33183 35649 33192 35683
rect 33140 35640 33192 35649
rect 34244 35640 34296 35692
rect 31852 35615 31904 35624
rect 30748 35479 30800 35488
rect 30748 35445 30757 35479
rect 30757 35445 30791 35479
rect 30791 35445 30800 35479
rect 30748 35436 30800 35445
rect 31852 35581 31861 35615
rect 31861 35581 31895 35615
rect 31895 35581 31904 35615
rect 31852 35572 31904 35581
rect 34980 35615 35032 35624
rect 34980 35581 34989 35615
rect 34989 35581 35023 35615
rect 35023 35581 35032 35615
rect 34980 35572 35032 35581
rect 56232 35615 56284 35624
rect 56232 35581 56241 35615
rect 56241 35581 56275 35615
rect 56275 35581 56284 35615
rect 56232 35572 56284 35581
rect 57704 35615 57756 35624
rect 57704 35581 57713 35615
rect 57713 35581 57747 35615
rect 57747 35581 57756 35615
rect 57704 35572 57756 35581
rect 31760 35479 31812 35488
rect 31760 35445 31769 35479
rect 31769 35445 31803 35479
rect 31803 35445 31812 35479
rect 31760 35436 31812 35445
rect 34428 35436 34480 35488
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 31852 35275 31904 35284
rect 31852 35241 31861 35275
rect 31861 35241 31895 35275
rect 31895 35241 31904 35275
rect 31852 35232 31904 35241
rect 34980 35232 35032 35284
rect 57704 35232 57756 35284
rect 30748 35207 30800 35216
rect 30748 35173 30782 35207
rect 30782 35173 30800 35207
rect 30748 35164 30800 35173
rect 18328 35096 18380 35148
rect 33232 35139 33284 35148
rect 27252 35028 27304 35080
rect 30472 35071 30524 35080
rect 30472 35037 30481 35071
rect 30481 35037 30515 35071
rect 30515 35037 30524 35071
rect 30472 35028 30524 35037
rect 33232 35105 33241 35139
rect 33241 35105 33275 35139
rect 33275 35105 33284 35139
rect 33232 35096 33284 35105
rect 33784 35096 33836 35148
rect 34428 35139 34480 35148
rect 34428 35105 34437 35139
rect 34437 35105 34471 35139
rect 34471 35105 34480 35139
rect 34428 35096 34480 35105
rect 57428 35139 57480 35148
rect 57428 35105 57437 35139
rect 57437 35105 57471 35139
rect 57471 35105 57480 35139
rect 57428 35096 57480 35105
rect 57520 35096 57572 35148
rect 57704 35096 57756 35148
rect 58072 35096 58124 35148
rect 33692 35071 33744 35080
rect 33692 35037 33701 35071
rect 33701 35037 33735 35071
rect 33735 35037 33744 35071
rect 33692 35028 33744 35037
rect 58164 35003 58216 35012
rect 58164 34969 58173 35003
rect 58173 34969 58207 35003
rect 58207 34969 58216 35003
rect 58164 34960 58216 34969
rect 20720 34892 20772 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 18328 34688 18380 34740
rect 27252 34688 27304 34740
rect 33232 34688 33284 34740
rect 34152 34688 34204 34740
rect 33784 34620 33836 34672
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 17868 34527 17920 34536
rect 17868 34493 17877 34527
rect 17877 34493 17911 34527
rect 17911 34493 17920 34527
rect 17868 34484 17920 34493
rect 20720 34484 20772 34536
rect 31024 34527 31076 34536
rect 31024 34493 31033 34527
rect 31033 34493 31067 34527
rect 31067 34493 31076 34527
rect 31024 34484 31076 34493
rect 31208 34527 31260 34536
rect 31208 34493 31217 34527
rect 31217 34493 31251 34527
rect 31251 34493 31260 34527
rect 31208 34484 31260 34493
rect 31300 34527 31352 34536
rect 31300 34493 31309 34527
rect 31309 34493 31343 34527
rect 31343 34493 31352 34527
rect 31300 34484 31352 34493
rect 31760 34527 31812 34536
rect 31760 34493 31769 34527
rect 31769 34493 31803 34527
rect 31803 34493 31812 34527
rect 31760 34484 31812 34493
rect 30840 34391 30892 34400
rect 30840 34357 30849 34391
rect 30849 34357 30883 34391
rect 30883 34357 30892 34391
rect 30840 34348 30892 34357
rect 33048 34391 33100 34400
rect 33048 34357 33057 34391
rect 33057 34357 33091 34391
rect 33091 34357 33100 34391
rect 33048 34348 33100 34357
rect 33324 34527 33376 34536
rect 33324 34493 33333 34527
rect 33333 34493 33367 34527
rect 33367 34493 33376 34527
rect 33324 34484 33376 34493
rect 33876 34552 33928 34604
rect 34060 34527 34112 34536
rect 34060 34493 34069 34527
rect 34069 34493 34103 34527
rect 34103 34493 34112 34527
rect 34060 34484 34112 34493
rect 57520 34552 57572 34604
rect 55312 34527 55364 34536
rect 55312 34493 55321 34527
rect 55321 34493 55355 34527
rect 55355 34493 55364 34527
rect 55312 34484 55364 34493
rect 57336 34484 57388 34536
rect 57428 34527 57480 34536
rect 57428 34493 57437 34527
rect 57437 34493 57471 34527
rect 57471 34493 57480 34527
rect 57428 34484 57480 34493
rect 57888 34484 57940 34536
rect 57060 34416 57112 34468
rect 57980 34459 58032 34468
rect 57980 34425 57989 34459
rect 57989 34425 58023 34459
rect 58023 34425 58032 34459
rect 57980 34416 58032 34425
rect 33876 34348 33928 34400
rect 34244 34348 34296 34400
rect 57244 34391 57296 34400
rect 57244 34357 57253 34391
rect 57253 34357 57287 34391
rect 57287 34357 57296 34391
rect 57244 34348 57296 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 20628 34008 20680 34060
rect 31300 34144 31352 34196
rect 33876 34144 33928 34196
rect 57980 34144 58032 34196
rect 30840 34076 30892 34128
rect 33048 34076 33100 34128
rect 33324 34076 33376 34128
rect 22652 34008 22704 34060
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 25688 34008 25740 34060
rect 19892 33940 19944 33992
rect 23112 33983 23164 33992
rect 23112 33949 23121 33983
rect 23121 33949 23155 33983
rect 23155 33949 23164 33983
rect 23112 33940 23164 33949
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 22928 33872 22980 33924
rect 23664 33804 23716 33856
rect 34152 34051 34204 34060
rect 34152 34017 34161 34051
rect 34161 34017 34195 34051
rect 34195 34017 34204 34051
rect 34152 34008 34204 34017
rect 35348 34008 35400 34060
rect 54116 34008 54168 34060
rect 55220 34008 55272 34060
rect 55864 34008 55916 34060
rect 57060 34051 57112 34060
rect 57060 34017 57069 34051
rect 57069 34017 57103 34051
rect 57103 34017 57112 34051
rect 57060 34008 57112 34017
rect 57520 34051 57572 34060
rect 57520 34017 57529 34051
rect 57529 34017 57563 34051
rect 57563 34017 57572 34051
rect 57520 34008 57572 34017
rect 35900 33804 35952 33856
rect 55772 33804 55824 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 20628 33643 20680 33652
rect 20628 33609 20637 33643
rect 20637 33609 20671 33643
rect 20671 33609 20680 33643
rect 20628 33600 20680 33609
rect 22192 33600 22244 33652
rect 54116 33643 54168 33652
rect 1400 33439 1452 33448
rect 1400 33405 1409 33439
rect 1409 33405 1443 33439
rect 1443 33405 1452 33439
rect 1400 33396 1452 33405
rect 20628 33439 20680 33448
rect 20628 33405 20637 33439
rect 20637 33405 20671 33439
rect 20671 33405 20680 33439
rect 20628 33396 20680 33405
rect 22100 33396 22152 33448
rect 22652 33439 22704 33448
rect 22652 33405 22661 33439
rect 22661 33405 22695 33439
rect 22695 33405 22704 33439
rect 22652 33396 22704 33405
rect 24952 33396 25004 33448
rect 31024 33532 31076 33584
rect 31852 33532 31904 33584
rect 32956 33532 33008 33584
rect 35348 33575 35400 33584
rect 35348 33541 35357 33575
rect 35357 33541 35391 33575
rect 35391 33541 35400 33575
rect 35348 33532 35400 33541
rect 31208 33439 31260 33448
rect 31208 33405 31217 33439
rect 31217 33405 31251 33439
rect 31251 33405 31260 33439
rect 31208 33396 31260 33405
rect 31300 33396 31352 33448
rect 32864 33396 32916 33448
rect 33232 33439 33284 33448
rect 33232 33405 33241 33439
rect 33241 33405 33275 33439
rect 33275 33405 33284 33439
rect 33232 33396 33284 33405
rect 33876 33396 33928 33448
rect 34244 33439 34296 33448
rect 34244 33405 34278 33439
rect 34278 33405 34296 33439
rect 34244 33396 34296 33405
rect 35900 33396 35952 33448
rect 36176 33396 36228 33448
rect 23940 33328 23992 33380
rect 34060 33328 34112 33380
rect 35716 33328 35768 33380
rect 21364 33303 21416 33312
rect 21364 33269 21373 33303
rect 21373 33269 21407 33303
rect 21407 33269 21416 33303
rect 21364 33260 21416 33269
rect 23664 33260 23716 33312
rect 24860 33303 24912 33312
rect 24860 33269 24869 33303
rect 24869 33269 24903 33303
rect 24903 33269 24912 33303
rect 24860 33260 24912 33269
rect 26148 33260 26200 33312
rect 34520 33260 34572 33312
rect 54116 33609 54125 33643
rect 54125 33609 54159 33643
rect 54159 33609 54168 33643
rect 54116 33600 54168 33609
rect 56968 33600 57020 33652
rect 57704 33600 57756 33652
rect 56784 33532 56836 33584
rect 57612 33532 57664 33584
rect 55036 33507 55088 33516
rect 55036 33473 55045 33507
rect 55045 33473 55079 33507
rect 55079 33473 55088 33507
rect 55036 33464 55088 33473
rect 57060 33507 57112 33516
rect 57060 33473 57069 33507
rect 57069 33473 57103 33507
rect 57103 33473 57112 33507
rect 57060 33464 57112 33473
rect 57244 33464 57296 33516
rect 54484 33371 54536 33380
rect 54484 33337 54493 33371
rect 54493 33337 54527 33371
rect 54527 33337 54536 33371
rect 54484 33328 54536 33337
rect 55772 33371 55824 33380
rect 55772 33337 55781 33371
rect 55781 33337 55815 33371
rect 55815 33337 55824 33371
rect 55772 33328 55824 33337
rect 56784 33328 56836 33380
rect 57336 33396 57388 33448
rect 58808 33328 58860 33380
rect 58164 33303 58216 33312
rect 58164 33269 58173 33303
rect 58173 33269 58207 33303
rect 58207 33269 58216 33303
rect 58164 33260 58216 33269
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 50326 33158 50378 33210
rect 50390 33158 50442 33210
rect 50454 33158 50506 33210
rect 50518 33158 50570 33210
rect 22100 33056 22152 33108
rect 23388 33099 23440 33108
rect 13728 32988 13780 33040
rect 23388 33065 23397 33099
rect 23397 33065 23431 33099
rect 23431 33065 23440 33099
rect 23388 33056 23440 33065
rect 23940 33099 23992 33108
rect 23940 33065 23949 33099
rect 23949 33065 23983 33099
rect 23983 33065 23992 33099
rect 23940 33056 23992 33065
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 21088 32920 21140 32972
rect 21364 32920 21416 32972
rect 22192 32920 22244 32972
rect 19892 32852 19944 32904
rect 22836 32963 22888 32972
rect 22836 32929 22845 32963
rect 22845 32929 22879 32963
rect 22879 32929 22888 32963
rect 22836 32920 22888 32929
rect 23572 32988 23624 33040
rect 32956 33056 33008 33108
rect 35716 33099 35768 33108
rect 35716 33065 35725 33099
rect 35725 33065 35759 33099
rect 35759 33065 35768 33099
rect 35716 33056 35768 33065
rect 34704 32988 34756 33040
rect 55864 33056 55916 33108
rect 23112 32963 23164 32972
rect 23112 32929 23121 32963
rect 23121 32929 23155 32963
rect 23155 32929 23164 32963
rect 23112 32920 23164 32929
rect 23848 32963 23900 32972
rect 22652 32852 22704 32904
rect 23848 32929 23857 32963
rect 23857 32929 23891 32963
rect 23891 32929 23900 32963
rect 23848 32920 23900 32929
rect 24032 32963 24084 32972
rect 24032 32929 24041 32963
rect 24041 32929 24075 32963
rect 24075 32929 24084 32963
rect 24032 32920 24084 32929
rect 24952 32920 25004 32972
rect 25780 32963 25832 32972
rect 25780 32929 25789 32963
rect 25789 32929 25823 32963
rect 25823 32929 25832 32963
rect 25780 32920 25832 32929
rect 31760 32963 31812 32972
rect 31760 32929 31769 32963
rect 31769 32929 31803 32963
rect 31803 32929 31812 32963
rect 31760 32920 31812 32929
rect 31852 32963 31904 32972
rect 31852 32929 31861 32963
rect 31861 32929 31895 32963
rect 31895 32929 31904 32963
rect 32864 32963 32916 32972
rect 31852 32920 31904 32929
rect 32864 32929 32873 32963
rect 32873 32929 32907 32963
rect 32907 32929 32916 32963
rect 32864 32920 32916 32929
rect 34520 32920 34572 32972
rect 35900 32963 35952 32972
rect 35900 32929 35909 32963
rect 35909 32929 35943 32963
rect 35943 32929 35952 32963
rect 35900 32920 35952 32929
rect 54576 32988 54628 33040
rect 58256 32988 58308 33040
rect 53840 32963 53892 32972
rect 53840 32929 53849 32963
rect 53849 32929 53883 32963
rect 53883 32929 53892 32963
rect 53840 32920 53892 32929
rect 56232 32920 56284 32972
rect 31668 32852 31720 32904
rect 33232 32852 33284 32904
rect 36176 32895 36228 32904
rect 36176 32861 36185 32895
rect 36185 32861 36219 32895
rect 36219 32861 36228 32895
rect 36176 32852 36228 32861
rect 49976 32852 50028 32904
rect 30932 32784 30984 32836
rect 34060 32784 34112 32836
rect 50344 32784 50396 32836
rect 54944 32827 54996 32836
rect 54944 32793 54953 32827
rect 54953 32793 54987 32827
rect 54987 32793 54996 32827
rect 54944 32784 54996 32793
rect 21640 32716 21692 32768
rect 22652 32716 22704 32768
rect 22836 32716 22888 32768
rect 23296 32716 23348 32768
rect 24860 32716 24912 32768
rect 31576 32759 31628 32768
rect 31576 32725 31585 32759
rect 31585 32725 31619 32759
rect 31619 32725 31628 32759
rect 31576 32716 31628 32725
rect 34152 32716 34204 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 20720 32512 20772 32564
rect 50344 32512 50396 32564
rect 54484 32512 54536 32564
rect 17040 32444 17092 32496
rect 20996 32444 21048 32496
rect 23296 32444 23348 32496
rect 13728 32419 13780 32428
rect 13728 32385 13737 32419
rect 13737 32385 13771 32419
rect 13771 32385 13780 32419
rect 13728 32376 13780 32385
rect 13360 32351 13412 32360
rect 13360 32317 13369 32351
rect 13369 32317 13403 32351
rect 13403 32317 13412 32351
rect 13360 32308 13412 32317
rect 13820 32308 13872 32360
rect 14924 32376 14976 32428
rect 15384 32308 15436 32360
rect 13176 32283 13228 32292
rect 13176 32249 13185 32283
rect 13185 32249 13219 32283
rect 13219 32249 13228 32283
rect 13176 32240 13228 32249
rect 13912 32240 13964 32292
rect 15568 32308 15620 32360
rect 18880 32308 18932 32360
rect 19432 32351 19484 32360
rect 19432 32317 19441 32351
rect 19441 32317 19475 32351
rect 19475 32317 19484 32351
rect 19432 32308 19484 32317
rect 20628 32308 20680 32360
rect 20996 32351 21048 32360
rect 20996 32317 21005 32351
rect 21005 32317 21039 32351
rect 21039 32317 21048 32351
rect 20996 32308 21048 32317
rect 21456 32351 21508 32360
rect 21456 32317 21465 32351
rect 21465 32317 21499 32351
rect 21499 32317 21508 32351
rect 21456 32308 21508 32317
rect 22836 32308 22888 32360
rect 31760 32444 31812 32496
rect 33232 32444 33284 32496
rect 55496 32444 55548 32496
rect 25688 32419 25740 32428
rect 25688 32385 25697 32419
rect 25697 32385 25731 32419
rect 25731 32385 25740 32419
rect 25688 32376 25740 32385
rect 30472 32376 30524 32428
rect 31668 32376 31720 32428
rect 22560 32240 22612 32292
rect 14740 32215 14792 32224
rect 14740 32181 14749 32215
rect 14749 32181 14783 32215
rect 14783 32181 14792 32215
rect 14740 32172 14792 32181
rect 16028 32172 16080 32224
rect 17960 32172 18012 32224
rect 19340 32172 19392 32224
rect 20444 32172 20496 32224
rect 20904 32215 20956 32224
rect 20904 32181 20913 32215
rect 20913 32181 20947 32215
rect 20947 32181 20956 32215
rect 20904 32172 20956 32181
rect 21180 32172 21232 32224
rect 23480 32308 23532 32360
rect 23940 32351 23992 32360
rect 23940 32317 23949 32351
rect 23949 32317 23983 32351
rect 23983 32317 23992 32351
rect 23940 32308 23992 32317
rect 24952 32351 25004 32360
rect 24952 32317 24961 32351
rect 24961 32317 24995 32351
rect 24995 32317 25004 32351
rect 24952 32308 25004 32317
rect 25412 32351 25464 32360
rect 25412 32317 25421 32351
rect 25421 32317 25455 32351
rect 25455 32317 25464 32351
rect 25412 32308 25464 32317
rect 26148 32351 26200 32360
rect 26148 32317 26157 32351
rect 26157 32317 26191 32351
rect 26191 32317 26200 32351
rect 26148 32308 26200 32317
rect 31576 32308 31628 32360
rect 23112 32283 23164 32292
rect 23112 32249 23121 32283
rect 23121 32249 23155 32283
rect 23155 32249 23164 32283
rect 23112 32240 23164 32249
rect 23572 32240 23624 32292
rect 24032 32283 24084 32292
rect 24032 32249 24041 32283
rect 24041 32249 24075 32283
rect 24075 32249 24084 32283
rect 24032 32240 24084 32249
rect 25780 32172 25832 32224
rect 33876 32351 33928 32360
rect 33876 32317 33885 32351
rect 33885 32317 33919 32351
rect 33919 32317 33928 32351
rect 33876 32308 33928 32317
rect 53840 32376 53892 32428
rect 55864 32376 55916 32428
rect 58532 32444 58584 32496
rect 57152 32419 57204 32428
rect 57152 32385 57161 32419
rect 57161 32385 57195 32419
rect 57195 32385 57204 32419
rect 57152 32376 57204 32385
rect 34244 32240 34296 32292
rect 54668 32308 54720 32360
rect 55036 32308 55088 32360
rect 58164 32308 58216 32360
rect 49976 32240 50028 32292
rect 34428 32172 34480 32224
rect 35716 32172 35768 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 50326 32070 50378 32122
rect 50390 32070 50442 32122
rect 50454 32070 50506 32122
rect 50518 32070 50570 32122
rect 16856 32011 16908 32020
rect 16856 31977 16865 32011
rect 16865 31977 16899 32011
rect 16899 31977 16908 32011
rect 16856 31968 16908 31977
rect 17868 31968 17920 32020
rect 19432 31968 19484 32020
rect 21088 31968 21140 32020
rect 12440 31943 12492 31952
rect 12440 31909 12449 31943
rect 12449 31909 12483 31943
rect 12483 31909 12492 31943
rect 12440 31900 12492 31909
rect 1400 31875 1452 31884
rect 1400 31841 1409 31875
rect 1409 31841 1443 31875
rect 1443 31841 1452 31875
rect 1400 31832 1452 31841
rect 12072 31832 12124 31884
rect 13268 31832 13320 31884
rect 12900 31764 12952 31816
rect 14556 31900 14608 31952
rect 14924 31875 14976 31884
rect 14924 31841 14933 31875
rect 14933 31841 14967 31875
rect 14967 31841 14976 31875
rect 14924 31832 14976 31841
rect 15476 31900 15528 31952
rect 15568 31875 15620 31884
rect 15568 31841 15577 31875
rect 15577 31841 15611 31875
rect 15611 31841 15620 31875
rect 15568 31832 15620 31841
rect 17684 31900 17736 31952
rect 17960 31943 18012 31952
rect 17960 31909 17994 31943
rect 17994 31909 18012 31943
rect 20720 31943 20772 31952
rect 17960 31900 18012 31909
rect 20720 31909 20729 31943
rect 20729 31909 20763 31943
rect 20763 31909 20772 31943
rect 20720 31900 20772 31909
rect 24952 31968 25004 32020
rect 33876 31968 33928 32020
rect 34244 32011 34296 32020
rect 34244 31977 34253 32011
rect 34253 31977 34287 32011
rect 34287 31977 34296 32011
rect 34244 31968 34296 31977
rect 17040 31875 17092 31884
rect 15016 31764 15068 31816
rect 16304 31807 16356 31816
rect 16304 31773 16313 31807
rect 16313 31773 16347 31807
rect 16347 31773 16356 31807
rect 16304 31764 16356 31773
rect 14004 31696 14056 31748
rect 17040 31841 17049 31875
rect 17049 31841 17083 31875
rect 17083 31841 17092 31875
rect 17040 31832 17092 31841
rect 19984 31875 20036 31884
rect 19984 31841 19993 31875
rect 19993 31841 20027 31875
rect 20027 31841 20036 31875
rect 19984 31832 20036 31841
rect 20444 31875 20496 31884
rect 20444 31841 20453 31875
rect 20453 31841 20487 31875
rect 20487 31841 20496 31875
rect 20444 31832 20496 31841
rect 19892 31764 19944 31816
rect 20536 31764 20588 31816
rect 21088 31832 21140 31884
rect 22100 31900 22152 31952
rect 22744 31900 22796 31952
rect 21824 31875 21876 31884
rect 12624 31628 12676 31680
rect 13452 31628 13504 31680
rect 14924 31671 14976 31680
rect 14924 31637 14933 31671
rect 14933 31637 14967 31671
rect 14967 31637 14976 31671
rect 14924 31628 14976 31637
rect 15108 31628 15160 31680
rect 19984 31696 20036 31748
rect 18052 31628 18104 31680
rect 20812 31628 20864 31680
rect 21824 31841 21833 31875
rect 21833 31841 21867 31875
rect 21867 31841 21876 31875
rect 21824 31832 21876 31841
rect 22468 31875 22520 31884
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 22560 31832 22612 31884
rect 22652 31807 22704 31816
rect 22652 31773 22661 31807
rect 22661 31773 22695 31807
rect 22695 31773 22704 31807
rect 22652 31764 22704 31773
rect 23388 31832 23440 31884
rect 25780 31900 25832 31952
rect 55680 31968 55732 32020
rect 56416 31968 56468 32020
rect 23848 31764 23900 31816
rect 24768 31764 24820 31816
rect 26332 31832 26384 31884
rect 55220 31943 55272 31952
rect 55220 31909 55229 31943
rect 55229 31909 55263 31943
rect 55263 31909 55272 31943
rect 55220 31900 55272 31909
rect 58348 31900 58400 31952
rect 27804 31832 27856 31884
rect 30472 31832 30524 31884
rect 32956 31832 33008 31884
rect 34428 31875 34480 31884
rect 34428 31841 34437 31875
rect 34437 31841 34471 31875
rect 34471 31841 34480 31875
rect 34428 31832 34480 31841
rect 34520 31875 34572 31884
rect 34520 31841 34529 31875
rect 34529 31841 34563 31875
rect 34563 31841 34572 31875
rect 34520 31832 34572 31841
rect 35716 31875 35768 31884
rect 27068 31807 27120 31816
rect 27068 31773 27077 31807
rect 27077 31773 27111 31807
rect 27111 31773 27120 31807
rect 27068 31764 27120 31773
rect 34704 31807 34756 31816
rect 34704 31773 34713 31807
rect 34713 31773 34747 31807
rect 34747 31773 34756 31807
rect 34704 31764 34756 31773
rect 35716 31841 35725 31875
rect 35725 31841 35759 31875
rect 35759 31841 35768 31875
rect 35716 31832 35768 31841
rect 53840 31832 53892 31884
rect 54668 31832 54720 31884
rect 56692 31832 56744 31884
rect 56968 31875 57020 31884
rect 56968 31841 56977 31875
rect 56977 31841 57011 31875
rect 57011 31841 57020 31875
rect 56968 31832 57020 31841
rect 36176 31764 36228 31816
rect 22744 31696 22796 31748
rect 23480 31696 23532 31748
rect 55220 31764 55272 31816
rect 57888 31764 57940 31816
rect 54576 31696 54628 31748
rect 23020 31628 23072 31680
rect 28448 31671 28500 31680
rect 28448 31637 28457 31671
rect 28457 31637 28491 31671
rect 28491 31637 28500 31671
rect 28448 31628 28500 31637
rect 33508 31671 33560 31680
rect 33508 31637 33517 31671
rect 33517 31637 33551 31671
rect 33551 31637 33560 31671
rect 33508 31628 33560 31637
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 12072 31424 12124 31476
rect 12256 31424 12308 31476
rect 19340 31424 19392 31476
rect 21824 31424 21876 31476
rect 23664 31424 23716 31476
rect 12624 31399 12676 31408
rect 12624 31365 12648 31399
rect 12648 31365 12676 31399
rect 12624 31356 12676 31365
rect 13268 31288 13320 31340
rect 19984 31356 20036 31408
rect 22836 31356 22888 31408
rect 12348 31220 12400 31272
rect 13636 31263 13688 31272
rect 13636 31229 13645 31263
rect 13645 31229 13679 31263
rect 13679 31229 13688 31263
rect 13636 31220 13688 31229
rect 15200 31220 15252 31272
rect 15660 31220 15712 31272
rect 18512 31288 18564 31340
rect 18880 31288 18932 31340
rect 13176 31195 13228 31204
rect 13176 31161 13185 31195
rect 13185 31161 13219 31195
rect 13219 31161 13228 31195
rect 13176 31152 13228 31161
rect 17500 31152 17552 31204
rect 18052 31263 18104 31272
rect 18052 31229 18061 31263
rect 18061 31229 18095 31263
rect 18095 31229 18104 31263
rect 18052 31220 18104 31229
rect 18420 31220 18472 31272
rect 19432 31220 19484 31272
rect 20076 31263 20128 31272
rect 20076 31229 20085 31263
rect 20085 31229 20119 31263
rect 20119 31229 20128 31263
rect 20076 31220 20128 31229
rect 21180 31263 21232 31272
rect 21180 31229 21187 31263
rect 21187 31229 21232 31263
rect 14556 31127 14608 31136
rect 14556 31093 14565 31127
rect 14565 31093 14599 31127
rect 14599 31093 14608 31127
rect 14556 31084 14608 31093
rect 17592 31127 17644 31136
rect 17592 31093 17601 31127
rect 17601 31093 17635 31127
rect 17635 31093 17644 31127
rect 17592 31084 17644 31093
rect 19156 31084 19208 31136
rect 19432 31084 19484 31136
rect 20628 31084 20680 31136
rect 21180 31220 21232 31229
rect 21640 31288 21692 31340
rect 22100 31288 22152 31340
rect 23480 31288 23532 31340
rect 27068 31424 27120 31476
rect 27252 31424 27304 31476
rect 27804 31467 27856 31476
rect 27804 31433 27813 31467
rect 27813 31433 27847 31467
rect 27847 31433 27856 31467
rect 27804 31424 27856 31433
rect 32956 31424 33008 31476
rect 33140 31424 33192 31476
rect 34060 31467 34112 31476
rect 34060 31433 34069 31467
rect 34069 31433 34103 31467
rect 34103 31433 34112 31467
rect 34060 31424 34112 31433
rect 34520 31424 34572 31476
rect 33508 31331 33560 31340
rect 33508 31297 33517 31331
rect 33517 31297 33551 31331
rect 33551 31297 33560 31331
rect 33508 31288 33560 31297
rect 21456 31263 21508 31272
rect 21456 31229 21470 31263
rect 21470 31229 21504 31263
rect 21504 31229 21508 31263
rect 21456 31220 21508 31229
rect 22744 31263 22796 31272
rect 22744 31229 22753 31263
rect 22753 31229 22787 31263
rect 22787 31229 22796 31263
rect 22744 31220 22796 31229
rect 23112 31263 23164 31272
rect 22468 31152 22520 31204
rect 23112 31229 23121 31263
rect 23121 31229 23155 31263
rect 23155 31229 23164 31263
rect 23112 31220 23164 31229
rect 23480 31152 23532 31204
rect 23848 31220 23900 31272
rect 24676 31220 24728 31272
rect 28172 31220 28224 31272
rect 25964 31152 26016 31204
rect 34704 31220 34756 31272
rect 56508 31356 56560 31408
rect 36544 31152 36596 31204
rect 54576 31195 54628 31204
rect 54576 31161 54585 31195
rect 54585 31161 54619 31195
rect 54619 31161 54628 31195
rect 54576 31152 54628 31161
rect 56876 31288 56928 31340
rect 58440 31288 58492 31340
rect 56232 31263 56284 31272
rect 56232 31229 56241 31263
rect 56241 31229 56275 31263
rect 56275 31229 56284 31263
rect 56232 31220 56284 31229
rect 23296 31084 23348 31136
rect 26516 31127 26568 31136
rect 26516 31093 26525 31127
rect 26525 31093 26559 31127
rect 26559 31093 26568 31127
rect 26516 31084 26568 31093
rect 55036 31084 55088 31136
rect 55772 31127 55824 31136
rect 55772 31093 55781 31127
rect 55781 31093 55815 31127
rect 55815 31093 55824 31127
rect 55772 31084 55824 31093
rect 56876 31127 56928 31136
rect 56876 31093 56885 31127
rect 56885 31093 56919 31127
rect 56919 31093 56928 31127
rect 57244 31195 57296 31204
rect 57244 31161 57253 31195
rect 57253 31161 57287 31195
rect 57287 31161 57296 31195
rect 57244 31152 57296 31161
rect 56876 31084 56928 31093
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 50326 30982 50378 31034
rect 50390 30982 50442 31034
rect 50454 30982 50506 31034
rect 50518 30982 50570 31034
rect 11428 30880 11480 30932
rect 13912 30880 13964 30932
rect 15384 30923 15436 30932
rect 15384 30889 15393 30923
rect 15393 30889 15427 30923
rect 15427 30889 15436 30923
rect 15384 30880 15436 30889
rect 16396 30880 16448 30932
rect 18420 30923 18472 30932
rect 18420 30889 18429 30923
rect 18429 30889 18463 30923
rect 18463 30889 18472 30923
rect 18420 30880 18472 30889
rect 20076 30880 20128 30932
rect 22468 30880 22520 30932
rect 25964 30923 26016 30932
rect 25964 30889 25973 30923
rect 25973 30889 26007 30923
rect 26007 30889 26016 30923
rect 25964 30880 26016 30889
rect 1400 30787 1452 30796
rect 1400 30753 1409 30787
rect 1409 30753 1443 30787
rect 1443 30753 1452 30787
rect 1400 30744 1452 30753
rect 10508 30787 10560 30796
rect 10508 30753 10517 30787
rect 10517 30753 10551 30787
rect 10551 30753 10560 30787
rect 10508 30744 10560 30753
rect 12440 30855 12492 30864
rect 12440 30821 12449 30855
rect 12449 30821 12483 30855
rect 12483 30821 12492 30855
rect 12440 30812 12492 30821
rect 11520 30676 11572 30728
rect 12992 30744 13044 30796
rect 17592 30812 17644 30864
rect 18604 30812 18656 30864
rect 20536 30812 20588 30864
rect 16764 30744 16816 30796
rect 17960 30787 18012 30796
rect 17960 30753 17967 30787
rect 17967 30753 18012 30787
rect 12532 30676 12584 30728
rect 12900 30676 12952 30728
rect 14372 30676 14424 30728
rect 15108 30676 15160 30728
rect 12256 30608 12308 30660
rect 17960 30744 18012 30753
rect 18144 30787 18196 30796
rect 18144 30753 18153 30787
rect 18153 30753 18187 30787
rect 18187 30753 18196 30787
rect 18144 30744 18196 30753
rect 18328 30744 18380 30796
rect 20076 30744 20128 30796
rect 20260 30787 20312 30796
rect 20260 30753 20294 30787
rect 20294 30753 20312 30787
rect 20260 30744 20312 30753
rect 21640 30744 21692 30796
rect 22376 30744 22428 30796
rect 19432 30608 19484 30660
rect 22468 30608 22520 30660
rect 23296 30787 23348 30796
rect 23296 30753 23305 30787
rect 23305 30753 23339 30787
rect 23339 30753 23348 30787
rect 23296 30744 23348 30753
rect 23664 30744 23716 30796
rect 23940 30676 23992 30728
rect 24492 30676 24544 30728
rect 26516 30744 26568 30796
rect 26976 30787 27028 30796
rect 26976 30753 26985 30787
rect 26985 30753 27019 30787
rect 27019 30753 27028 30787
rect 26976 30744 27028 30753
rect 54576 30880 54628 30932
rect 56416 30880 56468 30932
rect 55772 30812 55824 30864
rect 57796 30855 57848 30864
rect 57796 30821 57805 30855
rect 57805 30821 57839 30855
rect 57839 30821 57848 30855
rect 57796 30812 57848 30821
rect 27252 30676 27304 30728
rect 53840 30744 53892 30796
rect 55036 30744 55088 30796
rect 29828 30676 29880 30728
rect 56968 30676 57020 30728
rect 25504 30608 25556 30660
rect 8760 30540 8812 30592
rect 10416 30540 10468 30592
rect 12808 30540 12860 30592
rect 13728 30540 13780 30592
rect 16672 30540 16724 30592
rect 17500 30540 17552 30592
rect 17960 30540 18012 30592
rect 20720 30540 20772 30592
rect 23756 30583 23808 30592
rect 23756 30549 23765 30583
rect 23765 30549 23799 30583
rect 23799 30549 23808 30583
rect 23756 30540 23808 30549
rect 26700 30540 26752 30592
rect 26792 30540 26844 30592
rect 30104 30540 30156 30592
rect 57244 30608 57296 30660
rect 55680 30540 55732 30592
rect 56968 30540 57020 30592
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 1400 30175 1452 30184
rect 1400 30141 1409 30175
rect 1409 30141 1443 30175
rect 1443 30141 1452 30175
rect 1400 30132 1452 30141
rect 10508 30336 10560 30388
rect 12808 30336 12860 30388
rect 13636 30336 13688 30388
rect 13820 30379 13872 30388
rect 13820 30345 13829 30379
rect 13829 30345 13863 30379
rect 13863 30345 13872 30379
rect 13820 30336 13872 30345
rect 18328 30379 18380 30388
rect 18328 30345 18337 30379
rect 18337 30345 18371 30379
rect 18371 30345 18380 30379
rect 18328 30336 18380 30345
rect 12532 30268 12584 30320
rect 11428 30200 11480 30252
rect 12256 30200 12308 30252
rect 12900 30268 12952 30320
rect 15844 30268 15896 30320
rect 10968 30175 11020 30184
rect 10968 30141 10977 30175
rect 10977 30141 11011 30175
rect 11011 30141 11020 30175
rect 10968 30132 11020 30141
rect 12440 30175 12492 30184
rect 12440 30141 12449 30175
rect 12449 30141 12483 30175
rect 12483 30141 12492 30175
rect 12440 30132 12492 30141
rect 13176 30132 13228 30184
rect 15108 30175 15160 30184
rect 15108 30141 15117 30175
rect 15117 30141 15151 30175
rect 15151 30141 15160 30175
rect 15108 30132 15160 30141
rect 17132 30200 17184 30252
rect 18144 30268 18196 30320
rect 20260 30336 20312 30388
rect 19524 30268 19576 30320
rect 17868 30243 17920 30252
rect 16396 30175 16448 30184
rect 9588 29996 9640 30048
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 13084 30039 13136 30048
rect 13084 30005 13093 30039
rect 13093 30005 13127 30039
rect 13127 30005 13136 30039
rect 13084 29996 13136 30005
rect 13360 29996 13412 30048
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 16396 30141 16405 30175
rect 16405 30141 16439 30175
rect 16439 30141 16448 30175
rect 16396 30132 16448 30141
rect 16580 30132 16632 30184
rect 17500 30175 17552 30184
rect 17500 30141 17509 30175
rect 17509 30141 17543 30175
rect 17543 30141 17552 30175
rect 17500 30132 17552 30141
rect 17868 30209 17877 30243
rect 17877 30209 17911 30243
rect 17911 30209 17920 30243
rect 17868 30200 17920 30209
rect 18512 30175 18564 30184
rect 18512 30141 18521 30175
rect 18521 30141 18555 30175
rect 18555 30141 18564 30175
rect 18512 30132 18564 30141
rect 18696 30132 18748 30184
rect 17868 30064 17920 30116
rect 18972 30200 19024 30252
rect 19892 30200 19944 30252
rect 23664 30336 23716 30388
rect 25504 30379 25556 30388
rect 25504 30345 25513 30379
rect 25513 30345 25547 30379
rect 25547 30345 25556 30379
rect 25504 30336 25556 30345
rect 31116 30379 31168 30388
rect 20720 30311 20772 30320
rect 20720 30277 20729 30311
rect 20729 30277 20763 30311
rect 20763 30277 20772 30311
rect 20720 30268 20772 30277
rect 20996 30268 21048 30320
rect 22008 30268 22060 30320
rect 24492 30268 24544 30320
rect 26332 30268 26384 30320
rect 26608 30268 26660 30320
rect 26976 30268 27028 30320
rect 28724 30268 28776 30320
rect 29828 30311 29880 30320
rect 29828 30277 29837 30311
rect 29837 30277 29871 30311
rect 29871 30277 29880 30311
rect 29828 30268 29880 30277
rect 31116 30345 31125 30379
rect 31125 30345 31159 30379
rect 31159 30345 31168 30379
rect 31116 30336 31168 30345
rect 18880 30175 18932 30184
rect 18880 30141 18889 30175
rect 18889 30141 18923 30175
rect 18923 30141 18932 30175
rect 18880 30132 18932 30141
rect 19340 30064 19392 30116
rect 18880 29996 18932 30048
rect 19616 30175 19668 30184
rect 19616 30141 19625 30175
rect 19625 30141 19659 30175
rect 19659 30141 19668 30175
rect 27988 30200 28040 30252
rect 19616 30132 19668 30141
rect 19524 30064 19576 30116
rect 20996 30132 21048 30184
rect 22284 30132 22336 30184
rect 23204 30132 23256 30184
rect 23572 30132 23624 30184
rect 23756 30175 23808 30184
rect 23756 30141 23790 30175
rect 23790 30141 23808 30175
rect 23756 30132 23808 30141
rect 22652 30064 22704 30116
rect 24492 30064 24544 30116
rect 25780 30175 25832 30184
rect 25780 30141 25789 30175
rect 25789 30141 25823 30175
rect 25823 30141 25832 30175
rect 26056 30175 26108 30184
rect 25780 30132 25832 30141
rect 26056 30141 26065 30175
rect 26065 30141 26099 30175
rect 26099 30141 26108 30175
rect 26056 30132 26108 30141
rect 26516 30132 26568 30184
rect 26700 30132 26752 30184
rect 27436 30064 27488 30116
rect 28448 30132 28500 30184
rect 28632 30132 28684 30184
rect 29828 30175 29880 30184
rect 29828 30141 29837 30175
rect 29837 30141 29871 30175
rect 29871 30141 29880 30175
rect 29828 30132 29880 30141
rect 30012 30175 30064 30184
rect 30012 30141 30021 30175
rect 30021 30141 30055 30175
rect 30055 30141 30064 30175
rect 30472 30175 30524 30184
rect 30012 30132 30064 30141
rect 30472 30141 30481 30175
rect 30481 30141 30515 30175
rect 30515 30141 30524 30175
rect 30472 30132 30524 30141
rect 30656 30175 30708 30184
rect 30656 30141 30665 30175
rect 30665 30141 30699 30175
rect 30699 30141 30708 30175
rect 30656 30132 30708 30141
rect 28356 30064 28408 30116
rect 31484 30132 31536 30184
rect 35440 30175 35492 30184
rect 35440 30141 35449 30175
rect 35449 30141 35483 30175
rect 35483 30141 35492 30175
rect 35440 30132 35492 30141
rect 50068 30268 50120 30320
rect 55496 30268 55548 30320
rect 36544 30243 36596 30252
rect 36544 30209 36553 30243
rect 36553 30209 36587 30243
rect 36587 30209 36596 30243
rect 36544 30200 36596 30209
rect 50160 30200 50212 30252
rect 56876 30268 56928 30320
rect 57060 30311 57112 30320
rect 57060 30277 57069 30311
rect 57069 30277 57103 30311
rect 57103 30277 57112 30311
rect 57060 30268 57112 30277
rect 55680 30200 55732 30252
rect 54944 30132 54996 30184
rect 56140 30132 56192 30184
rect 22376 29996 22428 30048
rect 22744 29996 22796 30048
rect 25412 29996 25464 30048
rect 27988 29996 28040 30048
rect 28264 29996 28316 30048
rect 28724 29996 28776 30048
rect 30012 29996 30064 30048
rect 30104 29996 30156 30048
rect 55404 30107 55456 30116
rect 55404 30073 55413 30107
rect 55413 30073 55447 30107
rect 55447 30073 55456 30107
rect 55404 30064 55456 30073
rect 56048 29996 56100 30048
rect 57520 29996 57572 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 50326 29894 50378 29946
rect 50390 29894 50442 29946
rect 50454 29894 50506 29946
rect 50518 29894 50570 29946
rect 11060 29792 11112 29844
rect 15936 29792 15988 29844
rect 12348 29767 12400 29776
rect 1860 29699 1912 29708
rect 1860 29665 1869 29699
rect 1869 29665 1903 29699
rect 1903 29665 1912 29699
rect 1860 29656 1912 29665
rect 6460 29699 6512 29708
rect 6460 29665 6469 29699
rect 6469 29665 6503 29699
rect 6503 29665 6512 29699
rect 6460 29656 6512 29665
rect 7196 29656 7248 29708
rect 7288 29699 7340 29708
rect 7288 29665 7297 29699
rect 7297 29665 7331 29699
rect 7331 29665 7340 29699
rect 7288 29656 7340 29665
rect 8208 29656 8260 29708
rect 9404 29656 9456 29708
rect 12348 29733 12357 29767
rect 12357 29733 12391 29767
rect 12391 29733 12400 29767
rect 12348 29724 12400 29733
rect 11060 29656 11112 29708
rect 12532 29699 12584 29708
rect 12532 29665 12538 29699
rect 12538 29665 12584 29699
rect 12532 29656 12584 29665
rect 9588 29588 9640 29640
rect 12808 29656 12860 29708
rect 14740 29724 14792 29776
rect 15108 29724 15160 29776
rect 17868 29792 17920 29844
rect 16856 29724 16908 29776
rect 31576 29792 31628 29844
rect 20904 29724 20956 29776
rect 12900 29588 12952 29640
rect 15568 29656 15620 29708
rect 16396 29656 16448 29708
rect 16580 29699 16632 29708
rect 16580 29665 16589 29699
rect 16589 29665 16623 29699
rect 16623 29665 16632 29699
rect 16580 29656 16632 29665
rect 16672 29656 16724 29708
rect 17224 29699 17276 29708
rect 17224 29665 17233 29699
rect 17233 29665 17267 29699
rect 17267 29665 17276 29699
rect 17224 29656 17276 29665
rect 17684 29699 17736 29708
rect 17684 29665 17693 29699
rect 17693 29665 17727 29699
rect 17727 29665 17736 29699
rect 17684 29656 17736 29665
rect 18604 29699 18656 29708
rect 18604 29665 18613 29699
rect 18613 29665 18647 29699
rect 18647 29665 18656 29699
rect 18604 29656 18656 29665
rect 18696 29699 18748 29708
rect 18696 29665 18705 29699
rect 18705 29665 18739 29699
rect 18739 29665 18748 29699
rect 18696 29656 18748 29665
rect 14004 29588 14056 29640
rect 14372 29588 14424 29640
rect 15752 29588 15804 29640
rect 19156 29656 19208 29708
rect 20536 29656 20588 29708
rect 22652 29656 22704 29708
rect 23480 29656 23532 29708
rect 25044 29656 25096 29708
rect 20076 29588 20128 29640
rect 22928 29588 22980 29640
rect 23940 29588 23992 29640
rect 24952 29588 25004 29640
rect 12624 29563 12676 29572
rect 12624 29529 12633 29563
rect 12633 29529 12667 29563
rect 12667 29529 12676 29563
rect 12624 29520 12676 29529
rect 18512 29520 18564 29572
rect 19432 29520 19484 29572
rect 22284 29563 22336 29572
rect 22284 29529 22293 29563
rect 22293 29529 22327 29563
rect 22327 29529 22336 29563
rect 22284 29520 22336 29529
rect 22652 29520 22704 29572
rect 26240 29656 26292 29708
rect 26424 29699 26476 29708
rect 26424 29665 26433 29699
rect 26433 29665 26467 29699
rect 26467 29665 26476 29699
rect 26608 29699 26660 29708
rect 26424 29656 26476 29665
rect 26608 29665 26617 29699
rect 26617 29665 26651 29699
rect 26651 29665 26660 29699
rect 26608 29656 26660 29665
rect 26700 29699 26752 29708
rect 26700 29665 26709 29699
rect 26709 29665 26743 29699
rect 26743 29665 26752 29699
rect 26700 29656 26752 29665
rect 27804 29656 27856 29708
rect 28172 29699 28224 29708
rect 28172 29665 28181 29699
rect 28181 29665 28215 29699
rect 28215 29665 28224 29699
rect 28172 29656 28224 29665
rect 28264 29699 28316 29708
rect 28264 29665 28273 29699
rect 28273 29665 28307 29699
rect 28307 29665 28316 29699
rect 28264 29656 28316 29665
rect 28816 29656 28868 29708
rect 31116 29724 31168 29776
rect 50160 29792 50212 29844
rect 55404 29792 55456 29844
rect 31760 29724 31812 29776
rect 50068 29724 50120 29776
rect 54852 29724 54904 29776
rect 58624 29792 58676 29844
rect 56048 29724 56100 29776
rect 57704 29724 57756 29776
rect 28448 29631 28500 29640
rect 28448 29597 28457 29631
rect 28457 29597 28491 29631
rect 28491 29597 28500 29631
rect 28448 29588 28500 29597
rect 30380 29588 30432 29640
rect 28264 29520 28316 29572
rect 31576 29520 31628 29572
rect 54484 29656 54536 29708
rect 54944 29656 54996 29708
rect 57980 29699 58032 29708
rect 57980 29665 57989 29699
rect 57989 29665 58023 29699
rect 58023 29665 58032 29699
rect 57980 29656 58032 29665
rect 50252 29588 50304 29640
rect 50344 29520 50396 29572
rect 58164 29563 58216 29572
rect 58164 29529 58173 29563
rect 58173 29529 58207 29563
rect 58207 29529 58216 29563
rect 58164 29520 58216 29529
rect 1952 29495 2004 29504
rect 1952 29461 1961 29495
rect 1961 29461 1995 29495
rect 1995 29461 2004 29495
rect 1952 29452 2004 29461
rect 6552 29495 6604 29504
rect 6552 29461 6561 29495
rect 6561 29461 6595 29495
rect 6595 29461 6604 29495
rect 6552 29452 6604 29461
rect 7104 29495 7156 29504
rect 7104 29461 7113 29495
rect 7113 29461 7147 29495
rect 7147 29461 7156 29495
rect 7104 29452 7156 29461
rect 8116 29452 8168 29504
rect 9496 29495 9548 29504
rect 9496 29461 9505 29495
rect 9505 29461 9539 29495
rect 9539 29461 9548 29495
rect 9496 29452 9548 29461
rect 12072 29452 12124 29504
rect 13544 29452 13596 29504
rect 14740 29452 14792 29504
rect 17316 29452 17368 29504
rect 18604 29452 18656 29504
rect 21088 29452 21140 29504
rect 22836 29452 22888 29504
rect 24032 29452 24084 29504
rect 24860 29452 24912 29504
rect 25320 29495 25372 29504
rect 25320 29461 25329 29495
rect 25329 29461 25363 29495
rect 25363 29461 25372 29495
rect 25320 29452 25372 29461
rect 25872 29452 25924 29504
rect 27344 29452 27396 29504
rect 28080 29452 28132 29504
rect 30656 29452 30708 29504
rect 31760 29452 31812 29504
rect 35624 29452 35676 29504
rect 54484 29452 54536 29504
rect 56508 29452 56560 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 8208 29291 8260 29300
rect 8208 29257 8217 29291
rect 8217 29257 8251 29291
rect 8251 29257 8260 29291
rect 8208 29248 8260 29257
rect 11520 29248 11572 29300
rect 12256 29248 12308 29300
rect 15936 29248 15988 29300
rect 18512 29248 18564 29300
rect 18972 29248 19024 29300
rect 20444 29291 20496 29300
rect 20444 29257 20453 29291
rect 20453 29257 20487 29291
rect 20487 29257 20496 29291
rect 20444 29248 20496 29257
rect 8760 29155 8812 29164
rect 2964 29044 3016 29096
rect 6828 29087 6880 29096
rect 2044 29019 2096 29028
rect 2044 28985 2053 29019
rect 2053 28985 2087 29019
rect 2087 28985 2096 29019
rect 2044 28976 2096 28985
rect 6828 29053 6837 29087
rect 6837 29053 6871 29087
rect 6871 29053 6880 29087
rect 6828 29044 6880 29053
rect 8760 29121 8769 29155
rect 8769 29121 8803 29155
rect 8803 29121 8812 29155
rect 8760 29112 8812 29121
rect 6920 28976 6972 29028
rect 7104 29087 7156 29096
rect 7104 29053 7138 29087
rect 7138 29053 7156 29087
rect 7104 29044 7156 29053
rect 9496 29044 9548 29096
rect 12992 29180 13044 29232
rect 11152 29112 11204 29164
rect 15292 29180 15344 29232
rect 18696 29180 18748 29232
rect 12072 29087 12124 29096
rect 12072 29053 12081 29087
rect 12081 29053 12115 29087
rect 12115 29053 12124 29087
rect 12072 29044 12124 29053
rect 13084 29087 13136 29096
rect 13084 29053 13093 29087
rect 13093 29053 13127 29087
rect 13127 29053 13136 29087
rect 13084 29044 13136 29053
rect 15108 29044 15160 29096
rect 20536 29112 20588 29164
rect 7288 28976 7340 29028
rect 13820 28976 13872 29028
rect 14464 29019 14516 29028
rect 14464 28985 14473 29019
rect 14473 28985 14507 29019
rect 14507 28985 14516 29019
rect 14464 28976 14516 28985
rect 17224 29044 17276 29096
rect 17132 28976 17184 29028
rect 18052 29019 18104 29028
rect 18052 28985 18061 29019
rect 18061 28985 18095 29019
rect 18095 28985 18104 29019
rect 18052 28976 18104 28985
rect 19156 29087 19208 29096
rect 19156 29053 19165 29087
rect 19165 29053 19199 29087
rect 19199 29053 19208 29087
rect 19432 29087 19484 29096
rect 19156 29044 19208 29053
rect 19432 29053 19441 29087
rect 19441 29053 19475 29087
rect 19475 29053 19484 29087
rect 19432 29044 19484 29053
rect 21088 29248 21140 29300
rect 21824 29248 21876 29300
rect 22560 29248 22612 29300
rect 20904 29180 20956 29232
rect 24584 29248 24636 29300
rect 27896 29248 27948 29300
rect 28632 29248 28684 29300
rect 28816 29248 28868 29300
rect 22652 29112 22704 29164
rect 23112 29155 23164 29164
rect 23112 29121 23121 29155
rect 23121 29121 23155 29155
rect 23155 29121 23164 29155
rect 23112 29112 23164 29121
rect 23204 29155 23256 29164
rect 23204 29121 23213 29155
rect 23213 29121 23247 29155
rect 23247 29121 23256 29155
rect 23204 29112 23256 29121
rect 20904 29087 20956 29096
rect 20904 29053 20913 29087
rect 20913 29053 20947 29087
rect 20947 29053 20956 29087
rect 21088 29087 21140 29096
rect 20904 29044 20956 29053
rect 21088 29053 21097 29087
rect 21097 29053 21131 29087
rect 21131 29053 21140 29087
rect 21088 29044 21140 29053
rect 23296 29087 23348 29096
rect 23296 29053 23305 29087
rect 23305 29053 23339 29087
rect 23339 29053 23348 29087
rect 23296 29044 23348 29053
rect 24952 29180 25004 29232
rect 25780 29180 25832 29232
rect 26332 29180 26384 29232
rect 27528 29180 27580 29232
rect 24860 29112 24912 29164
rect 33324 29180 33376 29232
rect 50344 29248 50396 29300
rect 54852 29291 54904 29300
rect 54852 29257 54861 29291
rect 54861 29257 54895 29291
rect 54895 29257 54904 29291
rect 54852 29248 54904 29257
rect 56140 29291 56192 29300
rect 56140 29257 56149 29291
rect 56149 29257 56183 29291
rect 56183 29257 56192 29291
rect 56140 29248 56192 29257
rect 57980 29291 58032 29300
rect 57980 29257 57989 29291
rect 57989 29257 58023 29291
rect 58023 29257 58032 29291
rect 57980 29248 58032 29257
rect 55220 29180 55272 29232
rect 57152 29180 57204 29232
rect 24492 29087 24544 29096
rect 24492 29053 24501 29087
rect 24501 29053 24535 29087
rect 24535 29053 24544 29087
rect 24492 29044 24544 29053
rect 20536 28976 20588 29028
rect 21272 28976 21324 29028
rect 22652 28976 22704 29028
rect 22928 29019 22980 29028
rect 22928 28985 22937 29019
rect 22937 28985 22971 29019
rect 22971 28985 22980 29019
rect 22928 28976 22980 28985
rect 23480 28976 23532 29028
rect 23756 28976 23808 29028
rect 24584 28976 24636 29028
rect 5816 28951 5868 28960
rect 5816 28917 5825 28951
rect 5825 28917 5859 28951
rect 5859 28917 5868 28951
rect 5816 28908 5868 28917
rect 9772 28908 9824 28960
rect 10140 28908 10192 28960
rect 16488 28908 16540 28960
rect 20812 28908 20864 28960
rect 20996 28908 21048 28960
rect 22560 28908 22612 28960
rect 23296 28908 23348 28960
rect 23848 28951 23900 28960
rect 23848 28917 23857 28951
rect 23857 28917 23891 28951
rect 23891 28917 23900 28951
rect 23848 28908 23900 28917
rect 25044 29087 25096 29096
rect 25044 29053 25053 29087
rect 25053 29053 25087 29087
rect 25087 29053 25096 29087
rect 25044 29044 25096 29053
rect 25872 29087 25924 29096
rect 25872 29053 25881 29087
rect 25881 29053 25915 29087
rect 25915 29053 25924 29087
rect 25872 29044 25924 29053
rect 26148 29087 26200 29096
rect 26148 29053 26157 29087
rect 26157 29053 26191 29087
rect 26191 29053 26200 29087
rect 26148 29044 26200 29053
rect 26332 29044 26384 29096
rect 26424 29087 26476 29096
rect 26424 29053 26433 29087
rect 26433 29053 26467 29087
rect 26467 29053 26476 29087
rect 26424 29044 26476 29053
rect 26700 29044 26752 29096
rect 27988 29087 28040 29096
rect 27712 28976 27764 29028
rect 27988 29053 27997 29087
rect 27997 29053 28031 29087
rect 28031 29053 28040 29087
rect 27988 29044 28040 29053
rect 31208 29112 31260 29164
rect 28724 29044 28776 29096
rect 30380 29044 30432 29096
rect 29000 28976 29052 29028
rect 31576 29087 31628 29096
rect 31576 29053 31585 29087
rect 31585 29053 31619 29087
rect 31619 29053 31628 29087
rect 31576 29044 31628 29053
rect 50252 29112 50304 29164
rect 31116 28976 31168 29028
rect 27620 28908 27672 28960
rect 28356 28908 28408 28960
rect 31484 28908 31536 28960
rect 32036 28951 32088 28960
rect 32036 28917 32045 28951
rect 32045 28917 32079 28951
rect 32079 28917 32088 28951
rect 32036 28908 32088 28917
rect 33416 29087 33468 29096
rect 33416 29053 33425 29087
rect 33425 29053 33459 29087
rect 33459 29053 33468 29087
rect 33416 29044 33468 29053
rect 33692 29087 33744 29096
rect 33140 28976 33192 29028
rect 33692 29053 33701 29087
rect 33701 29053 33735 29087
rect 33735 29053 33744 29087
rect 33692 29044 33744 29053
rect 35440 29087 35492 29096
rect 35440 29053 35449 29087
rect 35449 29053 35483 29087
rect 35483 29053 35492 29087
rect 35440 29044 35492 29053
rect 35624 29087 35676 29096
rect 35624 29053 35633 29087
rect 35633 29053 35667 29087
rect 35667 29053 35676 29087
rect 35624 29044 35676 29053
rect 36452 29087 36504 29096
rect 36452 29053 36461 29087
rect 36461 29053 36495 29087
rect 36495 29053 36504 29087
rect 36452 29044 36504 29053
rect 55220 29044 55272 29096
rect 55680 29044 55732 29096
rect 56232 29044 56284 29096
rect 57428 29044 57480 29096
rect 57704 29087 57756 29096
rect 57704 29053 57713 29087
rect 57713 29053 57747 29087
rect 57747 29053 57756 29087
rect 57704 29044 57756 29053
rect 33508 28954 33560 29006
rect 57336 28976 57388 29028
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 50326 28806 50378 28858
rect 50390 28806 50442 28858
rect 50454 28806 50506 28858
rect 50518 28806 50570 28858
rect 6460 28704 6512 28756
rect 7196 28704 7248 28756
rect 9680 28704 9732 28756
rect 5816 28636 5868 28688
rect 12256 28704 12308 28756
rect 4712 28611 4764 28620
rect 1676 28543 1728 28552
rect 1676 28509 1685 28543
rect 1685 28509 1719 28543
rect 1719 28509 1728 28543
rect 1676 28500 1728 28509
rect 4712 28577 4721 28611
rect 4721 28577 4755 28611
rect 4755 28577 4764 28611
rect 4712 28568 4764 28577
rect 6828 28568 6880 28620
rect 7012 28611 7064 28620
rect 7012 28577 7021 28611
rect 7021 28577 7055 28611
rect 7055 28577 7064 28611
rect 7012 28568 7064 28577
rect 7288 28568 7340 28620
rect 8208 28611 8260 28620
rect 1860 28475 1912 28484
rect 1860 28441 1869 28475
rect 1869 28441 1903 28475
rect 1903 28441 1912 28475
rect 1860 28432 1912 28441
rect 2596 28364 2648 28416
rect 7564 28500 7616 28552
rect 8208 28577 8217 28611
rect 8217 28577 8251 28611
rect 8251 28577 8260 28611
rect 8208 28568 8260 28577
rect 9956 28568 10008 28620
rect 10140 28568 10192 28620
rect 11060 28636 11112 28688
rect 11336 28568 11388 28620
rect 11520 28611 11572 28620
rect 11520 28577 11529 28611
rect 11529 28577 11563 28611
rect 11563 28577 11572 28611
rect 11520 28568 11572 28577
rect 12900 28636 12952 28688
rect 13452 28636 13504 28688
rect 14924 28636 14976 28688
rect 12716 28611 12768 28620
rect 12716 28577 12725 28611
rect 12725 28577 12759 28611
rect 12759 28577 12768 28611
rect 12716 28568 12768 28577
rect 16488 28568 16540 28620
rect 17224 28611 17276 28620
rect 17224 28577 17233 28611
rect 17233 28577 17267 28611
rect 17267 28577 17276 28611
rect 17224 28568 17276 28577
rect 17776 28611 17828 28620
rect 17776 28577 17785 28611
rect 17785 28577 17819 28611
rect 17819 28577 17828 28611
rect 17776 28568 17828 28577
rect 18328 28568 18380 28620
rect 18604 28568 18656 28620
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 11428 28543 11480 28552
rect 9772 28432 9824 28484
rect 11428 28509 11437 28543
rect 11437 28509 11471 28543
rect 11471 28509 11480 28543
rect 11428 28500 11480 28509
rect 12624 28543 12676 28552
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 12624 28500 12676 28509
rect 14372 28500 14424 28552
rect 17868 28543 17920 28552
rect 17868 28509 17877 28543
rect 17877 28509 17911 28543
rect 17911 28509 17920 28543
rect 17868 28500 17920 28509
rect 17960 28500 18012 28552
rect 18880 28611 18932 28620
rect 18880 28577 18889 28611
rect 18889 28577 18923 28611
rect 18923 28577 18932 28611
rect 19064 28611 19116 28620
rect 18880 28568 18932 28577
rect 19064 28577 19073 28611
rect 19073 28577 19107 28611
rect 19107 28577 19116 28611
rect 19064 28568 19116 28577
rect 19156 28568 19208 28620
rect 20444 28636 20496 28688
rect 20996 28704 21048 28756
rect 21824 28747 21876 28756
rect 21824 28713 21833 28747
rect 21833 28713 21867 28747
rect 21867 28713 21876 28747
rect 21824 28704 21876 28713
rect 22928 28747 22980 28756
rect 22928 28713 22937 28747
rect 22937 28713 22971 28747
rect 22971 28713 22980 28747
rect 22928 28704 22980 28713
rect 24860 28704 24912 28756
rect 22836 28636 22888 28688
rect 21180 28568 21232 28620
rect 22008 28611 22060 28620
rect 22008 28577 22017 28611
rect 22017 28577 22051 28611
rect 22051 28577 22060 28611
rect 22008 28568 22060 28577
rect 19340 28500 19392 28552
rect 22560 28568 22612 28620
rect 23756 28636 23808 28688
rect 24032 28636 24084 28688
rect 23480 28611 23532 28620
rect 22284 28543 22336 28552
rect 15752 28432 15804 28484
rect 22284 28509 22293 28543
rect 22293 28509 22327 28543
rect 22327 28509 22336 28543
rect 22284 28500 22336 28509
rect 23480 28577 23489 28611
rect 23489 28577 23523 28611
rect 23523 28577 23532 28611
rect 23480 28568 23532 28577
rect 23940 28611 23992 28620
rect 23940 28577 23949 28611
rect 23949 28577 23983 28611
rect 23983 28577 23992 28611
rect 23940 28568 23992 28577
rect 25688 28568 25740 28620
rect 27804 28679 27856 28688
rect 7104 28364 7156 28416
rect 8116 28407 8168 28416
rect 8116 28373 8125 28407
rect 8125 28373 8159 28407
rect 8159 28373 8168 28407
rect 8116 28364 8168 28373
rect 9404 28364 9456 28416
rect 9956 28407 10008 28416
rect 9956 28373 9965 28407
rect 9965 28373 9999 28407
rect 9999 28373 10008 28407
rect 9956 28364 10008 28373
rect 13268 28364 13320 28416
rect 15108 28364 15160 28416
rect 16580 28364 16632 28416
rect 18236 28364 18288 28416
rect 22744 28432 22796 28484
rect 23940 28432 23992 28484
rect 26056 28500 26108 28552
rect 26884 28611 26936 28620
rect 26884 28577 26893 28611
rect 26893 28577 26927 28611
rect 26927 28577 26936 28611
rect 26884 28568 26936 28577
rect 27804 28645 27813 28679
rect 27813 28645 27847 28679
rect 27847 28645 27856 28679
rect 27804 28636 27856 28645
rect 29000 28704 29052 28756
rect 30380 28704 30432 28756
rect 27620 28568 27672 28620
rect 27344 28500 27396 28552
rect 27896 28611 27948 28620
rect 27896 28577 27910 28611
rect 27910 28577 27944 28611
rect 27944 28577 27948 28611
rect 27896 28568 27948 28577
rect 27804 28432 27856 28484
rect 28540 28500 28592 28552
rect 29000 28611 29052 28620
rect 29000 28577 29009 28611
rect 29009 28577 29043 28611
rect 29043 28577 29052 28611
rect 31024 28636 31076 28688
rect 31208 28679 31260 28688
rect 31208 28645 31217 28679
rect 31217 28645 31251 28679
rect 31251 28645 31260 28679
rect 31208 28636 31260 28645
rect 33692 28704 33744 28756
rect 32864 28636 32916 28688
rect 33232 28636 33284 28688
rect 33416 28636 33468 28688
rect 55312 28636 55364 28688
rect 58072 28704 58124 28756
rect 56232 28636 56284 28688
rect 58164 28679 58216 28688
rect 58164 28645 58173 28679
rect 58173 28645 58207 28679
rect 58207 28645 58216 28679
rect 58164 28636 58216 28645
rect 29000 28568 29052 28577
rect 31116 28611 31168 28620
rect 31116 28577 31125 28611
rect 31125 28577 31159 28611
rect 31159 28577 31168 28611
rect 31116 28568 31168 28577
rect 31760 28611 31812 28620
rect 31760 28577 31770 28611
rect 31770 28577 31804 28611
rect 31804 28577 31812 28611
rect 31944 28611 31996 28620
rect 31760 28568 31812 28577
rect 31944 28577 31953 28611
rect 31953 28577 31987 28611
rect 31987 28577 31996 28611
rect 31944 28568 31996 28577
rect 32036 28611 32088 28620
rect 32036 28577 32045 28611
rect 32045 28577 32079 28611
rect 32079 28577 32088 28611
rect 32036 28568 32088 28577
rect 33784 28568 33836 28620
rect 35716 28611 35768 28620
rect 35716 28577 35725 28611
rect 35725 28577 35759 28611
rect 35759 28577 35768 28611
rect 35716 28568 35768 28577
rect 31300 28432 31352 28484
rect 23204 28364 23256 28416
rect 25596 28364 25648 28416
rect 25872 28364 25924 28416
rect 32588 28500 32640 28552
rect 32864 28500 32916 28552
rect 58072 28568 58124 28620
rect 55128 28543 55180 28552
rect 55128 28509 55137 28543
rect 55137 28509 55171 28543
rect 55171 28509 55180 28543
rect 55128 28500 55180 28509
rect 56784 28543 56836 28552
rect 56784 28509 56793 28543
rect 56793 28509 56827 28543
rect 56827 28509 56836 28543
rect 56784 28500 56836 28509
rect 58716 28500 58768 28552
rect 55588 28432 55640 28484
rect 35440 28364 35492 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 2964 28203 3016 28212
rect 2964 28169 2973 28203
rect 2973 28169 3007 28203
rect 3007 28169 3016 28203
rect 2964 28160 3016 28169
rect 6920 28160 6972 28212
rect 2596 28067 2648 28076
rect 2596 28033 2605 28067
rect 2605 28033 2639 28067
rect 2639 28033 2648 28067
rect 2596 28024 2648 28033
rect 2780 27999 2832 28008
rect 2780 27965 2789 27999
rect 2789 27965 2823 27999
rect 2823 27965 2832 27999
rect 2780 27956 2832 27965
rect 4712 27956 4764 28008
rect 5080 27999 5132 28008
rect 5080 27965 5089 27999
rect 5089 27965 5123 27999
rect 5123 27965 5132 27999
rect 5080 27956 5132 27965
rect 1860 27931 1912 27940
rect 1860 27897 1869 27931
rect 1869 27897 1903 27931
rect 1903 27897 1912 27931
rect 1860 27888 1912 27897
rect 15752 28160 15804 28212
rect 17684 28160 17736 28212
rect 11244 28092 11296 28144
rect 11428 28092 11480 28144
rect 8116 28024 8168 28076
rect 9588 28024 9640 28076
rect 12992 28067 13044 28076
rect 7472 27956 7524 28008
rect 6552 27888 6604 27940
rect 8668 27956 8720 28008
rect 11152 27956 11204 28008
rect 11796 27956 11848 28008
rect 12072 27999 12124 28008
rect 12072 27965 12081 27999
rect 12081 27965 12115 27999
rect 12115 27965 12124 27999
rect 12072 27956 12124 27965
rect 12992 28033 13001 28067
rect 13001 28033 13035 28067
rect 13035 28033 13044 28067
rect 12992 28024 13044 28033
rect 15660 28092 15712 28144
rect 15936 28092 15988 28144
rect 17960 28092 18012 28144
rect 19064 28160 19116 28212
rect 21088 28160 21140 28212
rect 23112 28160 23164 28212
rect 15844 28024 15896 28076
rect 13176 27956 13228 28008
rect 13728 27999 13780 28008
rect 13728 27965 13737 27999
rect 13737 27965 13771 27999
rect 13771 27965 13780 27999
rect 13728 27956 13780 27965
rect 14464 27999 14516 28008
rect 14464 27965 14473 27999
rect 14473 27965 14507 27999
rect 14507 27965 14516 27999
rect 14464 27956 14516 27965
rect 15108 27999 15160 28008
rect 15108 27965 15117 27999
rect 15117 27965 15151 27999
rect 15151 27965 15160 27999
rect 15108 27956 15160 27965
rect 15200 27956 15252 28008
rect 15936 27999 15988 28008
rect 15936 27965 15945 27999
rect 15945 27965 15979 27999
rect 15979 27965 15988 27999
rect 15936 27956 15988 27965
rect 8484 27888 8536 27940
rect 10048 27888 10100 27940
rect 13912 27931 13964 27940
rect 13912 27897 13921 27931
rect 13921 27897 13955 27931
rect 13955 27897 13964 27931
rect 13912 27888 13964 27897
rect 15476 27888 15528 27940
rect 1952 27863 2004 27872
rect 1952 27829 1961 27863
rect 1961 27829 1995 27863
rect 1995 27829 2004 27863
rect 1952 27820 2004 27829
rect 4896 27820 4948 27872
rect 5080 27820 5132 27872
rect 10600 27820 10652 27872
rect 14004 27820 14056 27872
rect 15568 27820 15620 27872
rect 16212 27863 16264 27872
rect 16212 27829 16221 27863
rect 16221 27829 16255 27863
rect 16255 27829 16264 27863
rect 16212 27820 16264 27829
rect 19340 28135 19392 28144
rect 19340 28101 19349 28135
rect 19349 28101 19383 28135
rect 19383 28101 19392 28135
rect 19340 28092 19392 28101
rect 20536 28092 20588 28144
rect 17316 27999 17368 28008
rect 17316 27965 17325 27999
rect 17325 27965 17359 27999
rect 17359 27965 17368 27999
rect 17316 27956 17368 27965
rect 17592 27956 17644 28008
rect 17960 27999 18012 28008
rect 17960 27965 17969 27999
rect 17969 27965 18003 27999
rect 18003 27965 18012 27999
rect 17960 27956 18012 27965
rect 18052 27956 18104 28008
rect 18236 27999 18288 28008
rect 18236 27965 18270 27999
rect 18270 27965 18288 27999
rect 18236 27956 18288 27965
rect 18604 27956 18656 28008
rect 16488 27888 16540 27940
rect 20628 27999 20680 28008
rect 20628 27965 20637 27999
rect 20637 27965 20671 27999
rect 20671 27965 20680 27999
rect 20628 27956 20680 27965
rect 20720 27999 20772 28008
rect 20720 27965 20730 27999
rect 20730 27965 20764 27999
rect 20764 27965 20772 27999
rect 23388 28024 23440 28076
rect 25872 28160 25924 28212
rect 26148 28160 26200 28212
rect 27528 28160 27580 28212
rect 55312 28203 55364 28212
rect 26240 28092 26292 28144
rect 26332 28092 26384 28144
rect 26608 28092 26660 28144
rect 28080 28092 28132 28144
rect 20720 27956 20772 27965
rect 22284 27956 22336 28008
rect 23204 27999 23256 28008
rect 23204 27965 23213 27999
rect 23213 27965 23247 27999
rect 23247 27965 23256 27999
rect 23204 27956 23256 27965
rect 23848 27999 23900 28008
rect 23848 27965 23857 27999
rect 23857 27965 23891 27999
rect 23891 27965 23900 27999
rect 23848 27956 23900 27965
rect 25228 28024 25280 28076
rect 21364 27888 21416 27940
rect 21824 27888 21876 27940
rect 22560 27888 22612 27940
rect 23480 27888 23532 27940
rect 25688 27956 25740 28008
rect 26056 28024 26108 28076
rect 26148 27999 26200 28008
rect 26148 27965 26157 27999
rect 26157 27965 26191 27999
rect 26191 27965 26200 27999
rect 26148 27956 26200 27965
rect 26332 27956 26384 28008
rect 27344 27956 27396 28008
rect 28080 27999 28132 28008
rect 26056 27888 26108 27940
rect 28080 27965 28089 27999
rect 28089 27965 28123 27999
rect 28123 27965 28132 27999
rect 28080 27956 28132 27965
rect 27988 27931 28040 27940
rect 27988 27897 27997 27931
rect 27997 27897 28031 27931
rect 28031 27897 28040 27931
rect 27988 27888 28040 27897
rect 25320 27820 25372 27872
rect 26148 27820 26200 27872
rect 30380 27956 30432 28008
rect 30840 27956 30892 28008
rect 31208 28092 31260 28144
rect 31668 28024 31720 28076
rect 31760 28024 31812 28076
rect 33784 28067 33836 28076
rect 31208 27999 31260 28008
rect 31208 27965 31217 27999
rect 31217 27965 31251 27999
rect 31251 27965 31260 27999
rect 31208 27956 31260 27965
rect 31484 27956 31536 28008
rect 32036 27956 32088 28008
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 34336 27999 34388 28008
rect 34336 27965 34345 27999
rect 34345 27965 34379 27999
rect 34379 27965 34388 27999
rect 34336 27956 34388 27965
rect 55312 28169 55321 28203
rect 55321 28169 55355 28203
rect 55355 28169 55364 28203
rect 55312 28160 55364 28169
rect 56232 28203 56284 28212
rect 56232 28169 56241 28203
rect 56241 28169 56275 28203
rect 56275 28169 56284 28203
rect 56232 28160 56284 28169
rect 57704 28160 57756 28212
rect 56784 28024 56836 28076
rect 35440 27999 35492 28008
rect 35440 27965 35449 27999
rect 35449 27965 35483 27999
rect 35483 27965 35492 27999
rect 35440 27956 35492 27965
rect 35532 27999 35584 28008
rect 35532 27965 35541 27999
rect 35541 27965 35575 27999
rect 35575 27965 35584 27999
rect 36268 27999 36320 28008
rect 35532 27956 35584 27965
rect 36268 27965 36277 27999
rect 36277 27965 36311 27999
rect 36311 27965 36320 27999
rect 36268 27956 36320 27965
rect 34612 27888 34664 27940
rect 55220 27956 55272 28008
rect 57428 27999 57480 28008
rect 57428 27965 57437 27999
rect 57437 27965 57471 27999
rect 57471 27965 57480 27999
rect 57428 27956 57480 27965
rect 55128 27888 55180 27940
rect 57980 27931 58032 27940
rect 57980 27897 57989 27931
rect 57989 27897 58023 27931
rect 58023 27897 58032 27931
rect 57980 27888 58032 27897
rect 58164 27931 58216 27940
rect 58164 27897 58173 27931
rect 58173 27897 58207 27931
rect 58207 27897 58216 27931
rect 58164 27888 58216 27897
rect 29092 27820 29144 27872
rect 30288 27820 30340 27872
rect 30380 27820 30432 27872
rect 30932 27863 30984 27872
rect 30932 27829 30941 27863
rect 30941 27829 30975 27863
rect 30975 27829 30984 27863
rect 30932 27820 30984 27829
rect 31484 27820 31536 27872
rect 31668 27820 31720 27872
rect 31944 27820 31996 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 50326 27718 50378 27770
rect 50390 27718 50442 27770
rect 50454 27718 50506 27770
rect 50518 27718 50570 27770
rect 1676 27616 1728 27668
rect 2780 27616 2832 27668
rect 5448 27591 5500 27600
rect 2504 27480 2556 27532
rect 3332 27523 3384 27532
rect 3332 27489 3341 27523
rect 3341 27489 3375 27523
rect 3375 27489 3384 27523
rect 3332 27480 3384 27489
rect 5448 27557 5457 27591
rect 5457 27557 5491 27591
rect 5491 27557 5500 27591
rect 5448 27548 5500 27557
rect 7012 27616 7064 27668
rect 12440 27616 12492 27668
rect 13728 27616 13780 27668
rect 16212 27616 16264 27668
rect 18604 27616 18656 27668
rect 18880 27616 18932 27668
rect 20996 27616 21048 27668
rect 21180 27616 21232 27668
rect 9496 27548 9548 27600
rect 9864 27548 9916 27600
rect 5632 27412 5684 27464
rect 6460 27412 6512 27464
rect 7564 27480 7616 27532
rect 7748 27523 7800 27532
rect 7748 27489 7757 27523
rect 7757 27489 7791 27523
rect 7791 27489 7800 27523
rect 7748 27480 7800 27489
rect 8392 27480 8444 27532
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 9772 27523 9824 27532
rect 9772 27489 9781 27523
rect 9781 27489 9815 27523
rect 9815 27489 9824 27523
rect 10048 27523 10100 27532
rect 9772 27480 9824 27489
rect 10048 27489 10057 27523
rect 10057 27489 10091 27523
rect 10091 27489 10100 27523
rect 10048 27480 10100 27489
rect 10968 27548 11020 27600
rect 11152 27480 11204 27532
rect 14648 27480 14700 27532
rect 8116 27412 8168 27464
rect 9956 27455 10008 27464
rect 9956 27421 9965 27455
rect 9965 27421 9999 27455
rect 9999 27421 10008 27455
rect 9956 27412 10008 27421
rect 12624 27412 12676 27464
rect 13728 27455 13780 27464
rect 13728 27421 13737 27455
rect 13737 27421 13771 27455
rect 13771 27421 13780 27455
rect 13728 27412 13780 27421
rect 15476 27548 15528 27600
rect 15384 27523 15436 27532
rect 15384 27489 15393 27523
rect 15393 27489 15427 27523
rect 15427 27489 15436 27523
rect 15384 27480 15436 27489
rect 15568 27523 15620 27532
rect 15568 27489 15577 27523
rect 15577 27489 15611 27523
rect 15611 27489 15620 27523
rect 15568 27480 15620 27489
rect 15292 27412 15344 27464
rect 1400 27276 1452 27328
rect 4712 27276 4764 27328
rect 7288 27276 7340 27328
rect 8208 27276 8260 27328
rect 9496 27319 9548 27328
rect 9496 27285 9505 27319
rect 9505 27285 9539 27319
rect 9539 27285 9548 27319
rect 9496 27276 9548 27285
rect 9680 27276 9732 27328
rect 10968 27276 11020 27328
rect 12532 27344 12584 27396
rect 13820 27344 13872 27396
rect 15476 27387 15528 27396
rect 15476 27353 15485 27387
rect 15485 27353 15519 27387
rect 15519 27353 15528 27387
rect 15476 27344 15528 27353
rect 12256 27276 12308 27328
rect 12348 27276 12400 27328
rect 13544 27319 13596 27328
rect 13544 27285 13553 27319
rect 13553 27285 13587 27319
rect 13587 27285 13596 27319
rect 13544 27276 13596 27285
rect 14556 27276 14608 27328
rect 17040 27480 17092 27532
rect 17132 27412 17184 27464
rect 16488 27344 16540 27396
rect 17408 27480 17460 27532
rect 17592 27523 17644 27532
rect 17592 27489 17601 27523
rect 17601 27489 17635 27523
rect 17635 27489 17644 27523
rect 17592 27480 17644 27489
rect 18052 27480 18104 27532
rect 18604 27480 18656 27532
rect 22284 27548 22336 27600
rect 26884 27616 26936 27668
rect 29092 27659 29144 27668
rect 29092 27625 29101 27659
rect 29101 27625 29135 27659
rect 29135 27625 29144 27659
rect 29092 27616 29144 27625
rect 23572 27591 23624 27600
rect 17868 27412 17920 27464
rect 18512 27455 18564 27464
rect 18512 27421 18521 27455
rect 18521 27421 18555 27455
rect 18555 27421 18564 27455
rect 18512 27412 18564 27421
rect 20168 27480 20220 27532
rect 20444 27523 20496 27532
rect 20444 27489 20458 27523
rect 20458 27489 20492 27523
rect 20492 27489 20496 27523
rect 21180 27523 21232 27532
rect 20444 27480 20496 27489
rect 21180 27489 21189 27523
rect 21189 27489 21223 27523
rect 21223 27489 21232 27523
rect 21180 27480 21232 27489
rect 21364 27523 21416 27532
rect 21364 27489 21373 27523
rect 21373 27489 21407 27523
rect 21407 27489 21416 27523
rect 21364 27480 21416 27489
rect 21272 27455 21324 27464
rect 16120 27276 16172 27328
rect 17040 27319 17092 27328
rect 17040 27285 17049 27319
rect 17049 27285 17083 27319
rect 17083 27285 17092 27319
rect 17040 27276 17092 27285
rect 17592 27344 17644 27396
rect 18052 27319 18104 27328
rect 18052 27285 18061 27319
rect 18061 27285 18095 27319
rect 18095 27285 18104 27319
rect 18052 27276 18104 27285
rect 18144 27276 18196 27328
rect 20444 27276 20496 27328
rect 20628 27319 20680 27328
rect 20628 27285 20637 27319
rect 20637 27285 20671 27319
rect 20671 27285 20680 27319
rect 20628 27276 20680 27285
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 22008 27480 22060 27532
rect 23572 27557 23581 27591
rect 23581 27557 23615 27591
rect 23615 27557 23624 27591
rect 23572 27548 23624 27557
rect 21180 27344 21232 27396
rect 21916 27455 21968 27464
rect 21916 27421 21925 27455
rect 21925 27421 21959 27455
rect 21959 27421 21968 27455
rect 21916 27412 21968 27421
rect 21456 27344 21508 27396
rect 23480 27523 23532 27532
rect 23480 27489 23489 27523
rect 23489 27489 23523 27523
rect 23523 27489 23532 27523
rect 23480 27480 23532 27489
rect 24124 27523 24176 27532
rect 24124 27489 24133 27523
rect 24133 27489 24167 27523
rect 24167 27489 24176 27523
rect 24124 27480 24176 27489
rect 23204 27412 23256 27464
rect 24768 27548 24820 27600
rect 27988 27548 28040 27600
rect 30380 27548 30432 27600
rect 26148 27480 26200 27532
rect 26608 27523 26660 27532
rect 26608 27489 26617 27523
rect 26617 27489 26651 27523
rect 26651 27489 26660 27523
rect 27436 27523 27488 27532
rect 26608 27480 26660 27489
rect 27436 27489 27470 27523
rect 27470 27489 27488 27523
rect 27436 27480 27488 27489
rect 25688 27387 25740 27396
rect 25688 27353 25697 27387
rect 25697 27353 25731 27387
rect 25731 27353 25740 27387
rect 25688 27344 25740 27353
rect 25872 27344 25924 27396
rect 26424 27344 26476 27396
rect 25964 27276 26016 27328
rect 27160 27455 27212 27464
rect 27160 27421 27169 27455
rect 27169 27421 27203 27455
rect 27203 27421 27212 27455
rect 27160 27412 27212 27421
rect 30196 27480 30248 27532
rect 30840 27523 30892 27532
rect 30840 27489 30849 27523
rect 30849 27489 30883 27523
rect 30883 27489 30892 27523
rect 30840 27480 30892 27489
rect 31668 27548 31720 27600
rect 34612 27616 34664 27668
rect 57980 27616 58032 27668
rect 32956 27480 33008 27532
rect 33048 27480 33100 27532
rect 35716 27523 35768 27532
rect 35716 27489 35725 27523
rect 35725 27489 35759 27523
rect 35759 27489 35768 27523
rect 35716 27480 35768 27489
rect 55588 27523 55640 27532
rect 55588 27489 55597 27523
rect 55597 27489 55631 27523
rect 55631 27489 55640 27523
rect 55588 27480 55640 27489
rect 56048 27480 56100 27532
rect 32036 27412 32088 27464
rect 32864 27412 32916 27464
rect 33416 27455 33468 27464
rect 33416 27421 33425 27455
rect 33425 27421 33459 27455
rect 33459 27421 33468 27455
rect 33416 27412 33468 27421
rect 56784 27412 56836 27464
rect 57704 27455 57756 27464
rect 57704 27421 57713 27455
rect 57713 27421 57747 27455
rect 57747 27421 57756 27455
rect 57704 27412 57756 27421
rect 31760 27344 31812 27396
rect 30012 27276 30064 27328
rect 31208 27276 31260 27328
rect 31668 27319 31720 27328
rect 31668 27285 31677 27319
rect 31677 27285 31711 27319
rect 31711 27285 31720 27319
rect 31668 27276 31720 27285
rect 32864 27276 32916 27328
rect 34796 27319 34848 27328
rect 34796 27285 34805 27319
rect 34805 27285 34839 27319
rect 34839 27285 34848 27319
rect 34796 27276 34848 27285
rect 36360 27276 36412 27328
rect 56968 27319 57020 27328
rect 56968 27285 56977 27319
rect 56977 27285 57011 27319
rect 57011 27285 57020 27319
rect 56968 27276 57020 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 1860 27115 1912 27124
rect 1860 27081 1869 27115
rect 1869 27081 1903 27115
rect 1903 27081 1912 27115
rect 1860 27072 1912 27081
rect 5448 27115 5500 27124
rect 5448 27081 5457 27115
rect 5457 27081 5491 27115
rect 5491 27081 5500 27115
rect 5448 27072 5500 27081
rect 5632 27072 5684 27124
rect 10416 27072 10468 27124
rect 11152 27115 11204 27124
rect 11152 27081 11161 27115
rect 11161 27081 11195 27115
rect 11195 27081 11204 27115
rect 11152 27072 11204 27081
rect 8116 27004 8168 27056
rect 9956 27004 10008 27056
rect 3332 26936 3384 26988
rect 5448 26936 5500 26988
rect 6828 26979 6880 26988
rect 6828 26945 6837 26979
rect 6837 26945 6871 26979
rect 6871 26945 6880 26979
rect 6828 26936 6880 26945
rect 7932 26936 7984 26988
rect 9864 26936 9916 26988
rect 3424 26911 3476 26920
rect 3424 26877 3433 26911
rect 3433 26877 3467 26911
rect 3467 26877 3476 26911
rect 3424 26868 3476 26877
rect 4528 26911 4580 26920
rect 4528 26877 4537 26911
rect 4537 26877 4571 26911
rect 4571 26877 4580 26911
rect 4528 26868 4580 26877
rect 4712 26911 4764 26920
rect 4712 26877 4721 26911
rect 4721 26877 4755 26911
rect 4755 26877 4764 26911
rect 4712 26868 4764 26877
rect 5264 26911 5316 26920
rect 5264 26877 5273 26911
rect 5273 26877 5307 26911
rect 5307 26877 5316 26911
rect 7104 26911 7156 26920
rect 5264 26868 5316 26877
rect 5356 26800 5408 26852
rect 7104 26877 7138 26911
rect 7138 26877 7156 26911
rect 7104 26868 7156 26877
rect 8392 26868 8444 26920
rect 10140 26868 10192 26920
rect 10416 26911 10468 26920
rect 10416 26877 10425 26911
rect 10425 26877 10459 26911
rect 10459 26877 10468 26911
rect 10416 26868 10468 26877
rect 11244 27004 11296 27056
rect 14096 27072 14148 27124
rect 17316 27072 17368 27124
rect 17868 27072 17920 27124
rect 17960 27072 18012 27124
rect 21456 27072 21508 27124
rect 24124 27072 24176 27124
rect 24676 27115 24728 27124
rect 24676 27081 24685 27115
rect 24685 27081 24719 27115
rect 24719 27081 24728 27115
rect 24676 27072 24728 27081
rect 11612 27004 11664 27056
rect 8116 26800 8168 26852
rect 8576 26800 8628 26852
rect 10232 26800 10284 26852
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 12348 26936 12400 26988
rect 12624 26936 12676 26988
rect 10968 26868 11020 26877
rect 12440 26868 12492 26920
rect 12716 26911 12768 26920
rect 12716 26877 12725 26911
rect 12725 26877 12759 26911
rect 12759 26877 12768 26911
rect 12716 26868 12768 26877
rect 13360 26868 13412 26920
rect 13544 26911 13596 26920
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 15476 27004 15528 27056
rect 17776 27047 17828 27056
rect 17776 27013 17785 27047
rect 17785 27013 17819 27047
rect 17819 27013 17828 27047
rect 17776 27004 17828 27013
rect 13820 26936 13872 26988
rect 14648 26936 14700 26988
rect 17040 26936 17092 26988
rect 17224 26936 17276 26988
rect 17684 26936 17736 26988
rect 14188 26911 14240 26920
rect 13544 26868 13596 26877
rect 14188 26877 14197 26911
rect 14197 26877 14231 26911
rect 14231 26877 14240 26911
rect 14188 26868 14240 26877
rect 2044 26732 2096 26784
rect 3884 26775 3936 26784
rect 3884 26741 3893 26775
rect 3893 26741 3927 26775
rect 3927 26741 3936 26775
rect 3884 26732 3936 26741
rect 4160 26732 4212 26784
rect 7472 26732 7524 26784
rect 11428 26800 11480 26852
rect 14096 26800 14148 26852
rect 11336 26732 11388 26784
rect 12624 26732 12676 26784
rect 12992 26732 13044 26784
rect 13452 26732 13504 26784
rect 15844 26868 15896 26920
rect 16212 26911 16264 26920
rect 16212 26877 16221 26911
rect 16221 26877 16255 26911
rect 16255 26877 16264 26911
rect 16212 26868 16264 26877
rect 17500 26911 17552 26920
rect 17500 26877 17509 26911
rect 17509 26877 17543 26911
rect 17543 26877 17552 26911
rect 17500 26868 17552 26877
rect 17592 26911 17644 26920
rect 17592 26877 17601 26911
rect 17601 26877 17635 26911
rect 17635 26877 17644 26911
rect 17592 26868 17644 26877
rect 17868 26911 17920 26920
rect 17868 26877 17877 26911
rect 17877 26877 17911 26911
rect 17911 26877 17920 26911
rect 21088 26936 21140 26988
rect 17868 26868 17920 26877
rect 18696 26868 18748 26920
rect 18420 26843 18472 26852
rect 18420 26809 18429 26843
rect 18429 26809 18463 26843
rect 18463 26809 18472 26843
rect 18420 26800 18472 26809
rect 19432 26800 19484 26852
rect 21364 26868 21416 26920
rect 22652 26911 22704 26920
rect 22652 26877 22661 26911
rect 22661 26877 22695 26911
rect 22695 26877 22704 26911
rect 22652 26868 22704 26877
rect 25872 27072 25924 27124
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 26424 27072 26476 27124
rect 27160 27072 27212 27124
rect 27712 27072 27764 27124
rect 26608 27004 26660 27056
rect 29368 27072 29420 27124
rect 33048 27115 33100 27124
rect 25596 26936 25648 26988
rect 26516 26979 26568 26988
rect 25780 26868 25832 26920
rect 26516 26945 26525 26979
rect 26525 26945 26559 26979
rect 26559 26945 26568 26979
rect 32220 27004 32272 27056
rect 33048 27081 33057 27115
rect 33057 27081 33091 27115
rect 33091 27081 33100 27115
rect 33048 27072 33100 27081
rect 35532 27072 35584 27124
rect 56784 27115 56836 27124
rect 56784 27081 56793 27115
rect 56793 27081 56827 27115
rect 56827 27081 56836 27115
rect 56784 27072 56836 27081
rect 57704 27072 57756 27124
rect 33416 27004 33468 27056
rect 26516 26936 26568 26945
rect 32128 26936 32180 26988
rect 26792 26868 26844 26920
rect 27988 26911 28040 26920
rect 27988 26877 27997 26911
rect 27997 26877 28031 26911
rect 28031 26877 28040 26911
rect 27988 26868 28040 26877
rect 29000 26868 29052 26920
rect 19340 26732 19392 26784
rect 20720 26732 20772 26784
rect 21364 26732 21416 26784
rect 23020 26800 23072 26852
rect 24584 26843 24636 26852
rect 24584 26809 24593 26843
rect 24593 26809 24627 26843
rect 24627 26809 24636 26843
rect 24584 26800 24636 26809
rect 25228 26843 25280 26852
rect 25228 26809 25237 26843
rect 25237 26809 25271 26843
rect 25271 26809 25280 26843
rect 25228 26800 25280 26809
rect 29460 26868 29512 26920
rect 30012 26911 30064 26920
rect 30012 26877 30021 26911
rect 30021 26877 30055 26911
rect 30055 26877 30064 26911
rect 30012 26868 30064 26877
rect 30196 26911 30248 26920
rect 30196 26877 30205 26911
rect 30205 26877 30239 26911
rect 30239 26877 30248 26911
rect 30196 26868 30248 26877
rect 30380 26911 30432 26920
rect 30380 26877 30389 26911
rect 30389 26877 30423 26911
rect 30423 26877 30432 26911
rect 30380 26868 30432 26877
rect 22284 26732 22336 26784
rect 28540 26732 28592 26784
rect 30288 26843 30340 26852
rect 30288 26809 30297 26843
rect 30297 26809 30331 26843
rect 30331 26809 30340 26843
rect 30288 26800 30340 26809
rect 31392 26868 31444 26920
rect 31944 26868 31996 26920
rect 33324 26911 33376 26920
rect 33324 26877 33333 26911
rect 33333 26877 33367 26911
rect 33367 26877 33376 26911
rect 33324 26868 33376 26877
rect 33784 26936 33836 26988
rect 34704 26936 34756 26988
rect 56876 26936 56928 26988
rect 33508 26911 33560 26920
rect 33508 26877 33517 26911
rect 33517 26877 33551 26911
rect 33551 26877 33560 26911
rect 33508 26868 33560 26877
rect 33692 26911 33744 26920
rect 33692 26877 33701 26911
rect 33701 26877 33735 26911
rect 33735 26877 33744 26911
rect 33692 26868 33744 26877
rect 57428 26911 57480 26920
rect 31116 26800 31168 26852
rect 33048 26800 33100 26852
rect 57428 26877 57437 26911
rect 57437 26877 57471 26911
rect 57471 26877 57480 26911
rect 57428 26868 57480 26877
rect 37188 26800 37240 26852
rect 55404 26843 55456 26852
rect 55404 26809 55413 26843
rect 55413 26809 55447 26843
rect 55447 26809 55456 26843
rect 55404 26800 55456 26809
rect 55496 26843 55548 26852
rect 55496 26809 55505 26843
rect 55505 26809 55539 26843
rect 55539 26809 55548 26843
rect 57980 26843 58032 26852
rect 55496 26800 55548 26809
rect 57980 26809 57989 26843
rect 57989 26809 58023 26843
rect 58023 26809 58032 26843
rect 57980 26800 58032 26809
rect 31852 26775 31904 26784
rect 31852 26741 31861 26775
rect 31861 26741 31895 26775
rect 31895 26741 31904 26775
rect 31852 26732 31904 26741
rect 32772 26732 32824 26784
rect 35624 26732 35676 26784
rect 58348 26732 58400 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 50326 26630 50378 26682
rect 50390 26630 50442 26682
rect 50454 26630 50506 26682
rect 50518 26630 50570 26682
rect 2504 26571 2556 26580
rect 2504 26537 2513 26571
rect 2513 26537 2547 26571
rect 2547 26537 2556 26571
rect 2504 26528 2556 26537
rect 4528 26528 4580 26580
rect 7748 26528 7800 26580
rect 8484 26571 8536 26580
rect 8484 26537 8493 26571
rect 8493 26537 8527 26571
rect 8527 26537 8536 26571
rect 8484 26528 8536 26537
rect 9680 26528 9732 26580
rect 10876 26528 10928 26580
rect 11244 26528 11296 26580
rect 12348 26528 12400 26580
rect 12440 26528 12492 26580
rect 12624 26528 12676 26580
rect 16212 26528 16264 26580
rect 2044 26435 2096 26444
rect 2044 26401 2053 26435
rect 2053 26401 2087 26435
rect 2087 26401 2096 26435
rect 2044 26392 2096 26401
rect 3056 26435 3108 26444
rect 3056 26401 3065 26435
rect 3065 26401 3099 26435
rect 3099 26401 3108 26435
rect 3056 26392 3108 26401
rect 4712 26435 4764 26444
rect 4712 26401 4721 26435
rect 4721 26401 4755 26435
rect 4755 26401 4764 26435
rect 4712 26392 4764 26401
rect 5356 26435 5408 26444
rect 5356 26401 5365 26435
rect 5365 26401 5399 26435
rect 5399 26401 5408 26435
rect 5356 26392 5408 26401
rect 6184 26435 6236 26444
rect 6184 26401 6193 26435
rect 6193 26401 6227 26435
rect 6227 26401 6236 26435
rect 6184 26392 6236 26401
rect 6920 26392 6972 26444
rect 7012 26435 7064 26444
rect 7012 26401 7021 26435
rect 7021 26401 7055 26435
rect 7055 26401 7064 26435
rect 7472 26435 7524 26444
rect 7012 26392 7064 26401
rect 7472 26401 7481 26435
rect 7481 26401 7515 26435
rect 7515 26401 7524 26435
rect 7472 26392 7524 26401
rect 9496 26460 9548 26512
rect 7196 26256 7248 26308
rect 8208 26324 8260 26376
rect 9864 26392 9916 26444
rect 15016 26503 15068 26512
rect 15016 26469 15050 26503
rect 15050 26469 15068 26503
rect 15016 26460 15068 26469
rect 10324 26435 10376 26444
rect 10324 26401 10333 26435
rect 10333 26401 10367 26435
rect 10367 26401 10376 26435
rect 10324 26392 10376 26401
rect 10416 26392 10468 26444
rect 10784 26392 10836 26444
rect 11152 26435 11204 26444
rect 11152 26401 11161 26435
rect 11161 26401 11195 26435
rect 11195 26401 11204 26435
rect 11152 26392 11204 26401
rect 11428 26392 11480 26444
rect 11520 26435 11572 26444
rect 11520 26401 11529 26435
rect 11529 26401 11563 26435
rect 11563 26401 11572 26435
rect 11520 26392 11572 26401
rect 11980 26392 12032 26444
rect 12348 26435 12400 26444
rect 12348 26401 12357 26435
rect 12357 26401 12391 26435
rect 12391 26401 12400 26435
rect 12348 26392 12400 26401
rect 12440 26435 12492 26444
rect 12440 26401 12449 26435
rect 12449 26401 12483 26435
rect 12483 26401 12492 26435
rect 12716 26435 12768 26444
rect 12440 26392 12492 26401
rect 12716 26401 12725 26435
rect 12725 26401 12759 26435
rect 12759 26401 12768 26435
rect 12716 26392 12768 26401
rect 15476 26392 15528 26444
rect 16948 26528 17000 26580
rect 21364 26528 21416 26580
rect 17040 26460 17092 26512
rect 21824 26528 21876 26580
rect 23388 26528 23440 26580
rect 25596 26528 25648 26580
rect 30288 26528 30340 26580
rect 31944 26528 31996 26580
rect 32128 26571 32180 26580
rect 32128 26537 32137 26571
rect 32137 26537 32171 26571
rect 32171 26537 32180 26571
rect 32128 26528 32180 26537
rect 33692 26528 33744 26580
rect 37188 26571 37240 26580
rect 37188 26537 37197 26571
rect 37197 26537 37231 26571
rect 37231 26537 37240 26571
rect 37188 26528 37240 26537
rect 10232 26324 10284 26376
rect 11336 26367 11388 26376
rect 11336 26333 11345 26367
rect 11345 26333 11379 26367
rect 11379 26333 11388 26367
rect 11336 26324 11388 26333
rect 13176 26324 13228 26376
rect 13452 26324 13504 26376
rect 13820 26367 13872 26376
rect 13820 26333 13829 26367
rect 13829 26333 13863 26367
rect 13863 26333 13872 26367
rect 13820 26324 13872 26333
rect 14372 26324 14424 26376
rect 16212 26324 16264 26376
rect 16948 26392 17000 26444
rect 17500 26392 17552 26444
rect 17592 26392 17644 26444
rect 19340 26392 19392 26444
rect 19892 26392 19944 26444
rect 20812 26435 20864 26444
rect 17868 26367 17920 26376
rect 17868 26333 17877 26367
rect 17877 26333 17911 26367
rect 17911 26333 17920 26367
rect 18328 26367 18380 26376
rect 17868 26324 17920 26333
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 19064 26324 19116 26376
rect 20812 26401 20821 26435
rect 20821 26401 20855 26435
rect 20855 26401 20864 26435
rect 20812 26392 20864 26401
rect 21088 26392 21140 26444
rect 21456 26435 21508 26444
rect 21456 26401 21465 26435
rect 21465 26401 21499 26435
rect 21499 26401 21508 26435
rect 21456 26392 21508 26401
rect 23664 26460 23716 26512
rect 21824 26392 21876 26444
rect 22192 26392 22244 26444
rect 23388 26392 23440 26444
rect 25964 26460 26016 26512
rect 30564 26460 30616 26512
rect 31116 26503 31168 26512
rect 31116 26469 31125 26503
rect 31125 26469 31159 26503
rect 31159 26469 31168 26503
rect 32956 26503 33008 26512
rect 31116 26460 31168 26469
rect 26608 26435 26660 26444
rect 26608 26401 26617 26435
rect 26617 26401 26651 26435
rect 26651 26401 26660 26435
rect 26608 26392 26660 26401
rect 26792 26435 26844 26444
rect 26792 26401 26801 26435
rect 26801 26401 26835 26435
rect 26835 26401 26844 26435
rect 26792 26392 26844 26401
rect 26884 26435 26936 26444
rect 26884 26401 26893 26435
rect 26893 26401 26927 26435
rect 26927 26401 26936 26435
rect 26884 26392 26936 26401
rect 28264 26392 28316 26444
rect 29552 26392 29604 26444
rect 32956 26469 32965 26503
rect 32965 26469 32999 26503
rect 32999 26469 33008 26503
rect 32956 26460 33008 26469
rect 22008 26324 22060 26376
rect 25780 26367 25832 26376
rect 25780 26333 25789 26367
rect 25789 26333 25823 26367
rect 25823 26333 25832 26367
rect 25780 26324 25832 26333
rect 27160 26324 27212 26376
rect 27252 26324 27304 26376
rect 32312 26392 32364 26444
rect 32588 26435 32640 26444
rect 32588 26401 32597 26435
rect 32597 26401 32631 26435
rect 32631 26401 32640 26435
rect 32588 26392 32640 26401
rect 32772 26435 32824 26444
rect 32772 26401 32779 26435
rect 32779 26401 32824 26435
rect 32772 26392 32824 26401
rect 32864 26435 32916 26444
rect 32864 26401 32873 26435
rect 32873 26401 32907 26435
rect 32907 26401 32916 26435
rect 32864 26392 32916 26401
rect 33048 26435 33100 26444
rect 33784 26460 33836 26512
rect 34796 26460 34848 26512
rect 35808 26460 35860 26512
rect 33048 26401 33062 26435
rect 33062 26401 33096 26435
rect 33096 26401 33100 26435
rect 33048 26392 33100 26401
rect 33968 26435 34020 26444
rect 33968 26401 33977 26435
rect 33977 26401 34011 26435
rect 34011 26401 34020 26435
rect 33968 26392 34020 26401
rect 36360 26435 36412 26444
rect 32404 26324 32456 26376
rect 36360 26401 36369 26435
rect 36369 26401 36403 26435
rect 36403 26401 36412 26435
rect 36360 26392 36412 26401
rect 36636 26460 36688 26512
rect 37096 26435 37148 26444
rect 37096 26401 37105 26435
rect 37105 26401 37139 26435
rect 37139 26401 37148 26435
rect 37096 26392 37148 26401
rect 56692 26528 56744 26580
rect 57980 26528 58032 26580
rect 35256 26324 35308 26376
rect 55956 26324 56008 26376
rect 57980 26324 58032 26376
rect 3148 26231 3200 26240
rect 3148 26197 3157 26231
rect 3157 26197 3191 26231
rect 3191 26197 3200 26231
rect 3148 26188 3200 26197
rect 6276 26231 6328 26240
rect 6276 26197 6285 26231
rect 6285 26197 6319 26231
rect 6319 26197 6328 26231
rect 6276 26188 6328 26197
rect 6736 26188 6788 26240
rect 9680 26188 9732 26240
rect 13544 26256 13596 26308
rect 17316 26256 17368 26308
rect 10048 26188 10100 26240
rect 10508 26231 10560 26240
rect 10508 26197 10517 26231
rect 10517 26197 10551 26231
rect 10551 26197 10560 26231
rect 10508 26188 10560 26197
rect 11704 26231 11756 26240
rect 11704 26197 11713 26231
rect 11713 26197 11747 26231
rect 11747 26197 11756 26231
rect 11704 26188 11756 26197
rect 12900 26231 12952 26240
rect 12900 26197 12909 26231
rect 12909 26197 12943 26231
rect 12943 26197 12952 26231
rect 12900 26188 12952 26197
rect 15476 26188 15528 26240
rect 17132 26188 17184 26240
rect 21088 26188 21140 26240
rect 21272 26231 21324 26240
rect 21272 26197 21281 26231
rect 21281 26197 21315 26231
rect 21315 26197 21324 26231
rect 21272 26188 21324 26197
rect 21824 26256 21876 26308
rect 21640 26188 21692 26240
rect 23664 26188 23716 26240
rect 25504 26231 25556 26240
rect 25504 26197 25513 26231
rect 25513 26197 25547 26231
rect 25547 26197 25556 26231
rect 25504 26188 25556 26197
rect 25872 26256 25924 26308
rect 27804 26256 27856 26308
rect 34520 26256 34572 26308
rect 55404 26256 55456 26308
rect 29184 26188 29236 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 3056 25984 3108 26036
rect 4068 25916 4120 25968
rect 3884 25848 3936 25900
rect 3608 25823 3660 25832
rect 3608 25789 3617 25823
rect 3617 25789 3651 25823
rect 3651 25789 3660 25823
rect 3608 25780 3660 25789
rect 3976 25780 4028 25832
rect 6184 25984 6236 26036
rect 7564 25984 7616 26036
rect 25228 25984 25280 26036
rect 25780 25984 25832 26036
rect 29368 26027 29420 26036
rect 8484 25916 8536 25968
rect 10048 25916 10100 25968
rect 19064 25916 19116 25968
rect 19432 25916 19484 25968
rect 21364 25916 21416 25968
rect 26148 25916 26200 25968
rect 29368 25993 29377 26027
rect 29377 25993 29411 26027
rect 29411 25993 29420 26027
rect 29368 25984 29420 25993
rect 30196 25984 30248 26036
rect 32588 25984 32640 26036
rect 33048 26027 33100 26036
rect 33048 25993 33057 26027
rect 33057 25993 33091 26027
rect 33091 25993 33100 26027
rect 33048 25984 33100 25993
rect 35256 25984 35308 26036
rect 55496 25984 55548 26036
rect 55956 26027 56008 26036
rect 55956 25993 55965 26027
rect 55965 25993 55999 26027
rect 55999 25993 56008 26027
rect 55956 25984 56008 25993
rect 6736 25780 6788 25832
rect 18328 25848 18380 25900
rect 19248 25891 19300 25900
rect 19248 25857 19257 25891
rect 19257 25857 19291 25891
rect 19291 25857 19300 25891
rect 19248 25848 19300 25857
rect 31116 25959 31168 25968
rect 31116 25925 31125 25959
rect 31125 25925 31159 25959
rect 31159 25925 31168 25959
rect 31116 25916 31168 25925
rect 33324 25916 33376 25968
rect 33968 25916 34020 25968
rect 34244 25916 34296 25968
rect 35624 25916 35676 25968
rect 7932 25780 7984 25832
rect 8668 25780 8720 25832
rect 10508 25780 10560 25832
rect 10600 25823 10652 25832
rect 10600 25789 10609 25823
rect 10609 25789 10643 25823
rect 10643 25789 10652 25823
rect 10600 25780 10652 25789
rect 11060 25780 11112 25832
rect 12900 25780 12952 25832
rect 15108 25823 15160 25832
rect 5172 25712 5224 25764
rect 7196 25755 7248 25764
rect 7196 25721 7230 25755
rect 7230 25721 7248 25755
rect 7196 25712 7248 25721
rect 7656 25712 7708 25764
rect 2872 25644 2924 25696
rect 4068 25644 4120 25696
rect 9864 25644 9916 25696
rect 10324 25712 10376 25764
rect 13636 25712 13688 25764
rect 14280 25712 14332 25764
rect 15108 25789 15117 25823
rect 15117 25789 15151 25823
rect 15151 25789 15160 25823
rect 15108 25780 15160 25789
rect 15568 25823 15620 25832
rect 15568 25789 15577 25823
rect 15577 25789 15611 25823
rect 15611 25789 15620 25823
rect 15568 25780 15620 25789
rect 16212 25823 16264 25832
rect 16212 25789 16221 25823
rect 16221 25789 16255 25823
rect 16255 25789 16264 25823
rect 16212 25780 16264 25789
rect 17960 25780 18012 25832
rect 18880 25823 18932 25832
rect 18880 25789 18911 25823
rect 18911 25789 18932 25823
rect 18880 25780 18932 25789
rect 18512 25712 18564 25764
rect 18972 25712 19024 25764
rect 12716 25644 12768 25696
rect 15384 25644 15436 25696
rect 16948 25644 17000 25696
rect 17316 25644 17368 25696
rect 18236 25644 18288 25696
rect 18604 25644 18656 25696
rect 18788 25644 18840 25696
rect 20168 25780 20220 25832
rect 20996 25780 21048 25832
rect 21364 25780 21416 25832
rect 21456 25780 21508 25832
rect 22284 25780 22336 25832
rect 22652 25780 22704 25832
rect 23296 25780 23348 25832
rect 25964 25823 26016 25832
rect 25964 25789 25973 25823
rect 25973 25789 26007 25823
rect 26007 25789 26016 25823
rect 25964 25780 26016 25789
rect 26148 25823 26200 25832
rect 26148 25789 26157 25823
rect 26157 25789 26191 25823
rect 26191 25789 26200 25823
rect 26148 25780 26200 25789
rect 26240 25823 26292 25832
rect 26240 25789 26249 25823
rect 26249 25789 26283 25823
rect 26283 25789 26292 25823
rect 26516 25823 26568 25832
rect 26240 25780 26292 25789
rect 26516 25789 26525 25823
rect 26525 25789 26559 25823
rect 26559 25789 26568 25823
rect 26516 25780 26568 25789
rect 28264 25780 28316 25832
rect 30288 25780 30340 25832
rect 32128 25848 32180 25900
rect 32588 25848 32640 25900
rect 34336 25891 34388 25900
rect 22192 25644 22244 25696
rect 24584 25644 24636 25696
rect 29644 25712 29696 25764
rect 29828 25644 29880 25696
rect 30472 25644 30524 25696
rect 31208 25823 31260 25832
rect 31208 25789 31217 25823
rect 31217 25789 31251 25823
rect 31251 25789 31260 25823
rect 31208 25780 31260 25789
rect 31852 25780 31904 25832
rect 32404 25780 32456 25832
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 36636 25891 36688 25900
rect 36636 25857 36645 25891
rect 36645 25857 36679 25891
rect 36679 25857 36688 25891
rect 36636 25848 36688 25857
rect 34060 25823 34112 25832
rect 32680 25712 32732 25764
rect 34060 25789 34069 25823
rect 34069 25789 34103 25823
rect 34103 25789 34112 25823
rect 34796 25823 34848 25832
rect 34060 25780 34112 25789
rect 34796 25789 34805 25823
rect 34805 25789 34839 25823
rect 34839 25789 34848 25823
rect 34796 25780 34848 25789
rect 35624 25823 35676 25832
rect 35624 25789 35633 25823
rect 35633 25789 35667 25823
rect 35667 25789 35676 25823
rect 35624 25780 35676 25789
rect 36360 25823 36412 25832
rect 36360 25789 36369 25823
rect 36369 25789 36403 25823
rect 36403 25789 36412 25823
rect 36360 25780 36412 25789
rect 35992 25712 36044 25764
rect 55680 25780 55732 25832
rect 56508 25780 56560 25832
rect 56876 25780 56928 25832
rect 57612 25780 57664 25832
rect 58256 25780 58308 25832
rect 58164 25755 58216 25764
rect 58164 25721 58173 25755
rect 58173 25721 58207 25755
rect 58207 25721 58216 25755
rect 58164 25712 58216 25721
rect 31300 25644 31352 25696
rect 33140 25644 33192 25696
rect 34428 25644 34480 25696
rect 34520 25644 34572 25696
rect 35808 25644 35860 25696
rect 57060 25644 57112 25696
rect 57428 25687 57480 25696
rect 57428 25653 57437 25687
rect 57437 25653 57471 25687
rect 57471 25653 57480 25687
rect 57428 25644 57480 25653
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 50326 25542 50378 25594
rect 50390 25542 50442 25594
rect 50454 25542 50506 25594
rect 50518 25542 50570 25594
rect 5172 25483 5224 25492
rect 5172 25449 5181 25483
rect 5181 25449 5215 25483
rect 5215 25449 5224 25483
rect 5172 25440 5224 25449
rect 6828 25440 6880 25492
rect 6920 25440 6972 25492
rect 17960 25483 18012 25492
rect 1860 25347 1912 25356
rect 1860 25313 1869 25347
rect 1869 25313 1903 25347
rect 1903 25313 1912 25347
rect 1860 25304 1912 25313
rect 3608 25304 3660 25356
rect 4068 25304 4120 25356
rect 5264 25347 5316 25356
rect 5264 25313 5273 25347
rect 5273 25313 5307 25347
rect 5307 25313 5316 25347
rect 7564 25372 7616 25424
rect 5264 25304 5316 25313
rect 6000 25347 6052 25356
rect 6000 25313 6009 25347
rect 6009 25313 6043 25347
rect 6043 25313 6052 25347
rect 6000 25304 6052 25313
rect 6184 25304 6236 25356
rect 7840 25372 7892 25424
rect 9772 25415 9824 25424
rect 9772 25381 9781 25415
rect 9781 25381 9815 25415
rect 9815 25381 9824 25415
rect 9772 25372 9824 25381
rect 11704 25372 11756 25424
rect 13636 25415 13688 25424
rect 13636 25381 13645 25415
rect 13645 25381 13679 25415
rect 13679 25381 13688 25415
rect 13636 25372 13688 25381
rect 7012 25279 7064 25288
rect 7012 25245 7021 25279
rect 7021 25245 7055 25279
rect 7055 25245 7064 25279
rect 7012 25236 7064 25245
rect 8024 25347 8076 25356
rect 8024 25313 8033 25347
rect 8033 25313 8067 25347
rect 8067 25313 8076 25347
rect 8024 25304 8076 25313
rect 9588 25347 9640 25356
rect 9588 25313 9597 25347
rect 9597 25313 9631 25347
rect 9631 25313 9640 25347
rect 9588 25304 9640 25313
rect 8392 25236 8444 25288
rect 12716 25304 12768 25356
rect 14648 25304 14700 25356
rect 14832 25304 14884 25356
rect 1952 25143 2004 25152
rect 1952 25109 1961 25143
rect 1961 25109 1995 25143
rect 1995 25109 2004 25143
rect 1952 25100 2004 25109
rect 3332 25143 3384 25152
rect 3332 25109 3341 25143
rect 3341 25109 3375 25143
rect 3375 25109 3384 25143
rect 3332 25100 3384 25109
rect 4620 25143 4672 25152
rect 4620 25109 4629 25143
rect 4629 25109 4663 25143
rect 4663 25109 4672 25143
rect 4620 25100 4672 25109
rect 6552 25100 6604 25152
rect 6828 25100 6880 25152
rect 7656 25100 7708 25152
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 11060 25100 11112 25152
rect 11152 25100 11204 25152
rect 15660 25236 15712 25288
rect 17960 25449 17969 25483
rect 17969 25449 18003 25483
rect 18003 25449 18012 25483
rect 17960 25440 18012 25449
rect 18144 25440 18196 25492
rect 21364 25483 21416 25492
rect 16304 25372 16356 25424
rect 16212 25304 16264 25356
rect 16672 25347 16724 25356
rect 16672 25313 16681 25347
rect 16681 25313 16715 25347
rect 16715 25313 16724 25347
rect 16672 25304 16724 25313
rect 16856 25304 16908 25356
rect 17316 25347 17368 25356
rect 17316 25313 17325 25347
rect 17325 25313 17359 25347
rect 17359 25313 17368 25347
rect 17316 25304 17368 25313
rect 18512 25372 18564 25424
rect 20628 25372 20680 25424
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 22192 25440 22244 25492
rect 22836 25440 22888 25492
rect 23480 25440 23532 25492
rect 28264 25483 28316 25492
rect 21640 25372 21692 25424
rect 22376 25372 22428 25424
rect 18420 25347 18472 25356
rect 18420 25313 18434 25347
rect 18434 25313 18468 25347
rect 18468 25313 18472 25347
rect 18420 25304 18472 25313
rect 18880 25304 18932 25356
rect 23572 25304 23624 25356
rect 17500 25236 17552 25288
rect 17592 25236 17644 25288
rect 21548 25236 21600 25288
rect 12164 25143 12216 25152
rect 12164 25109 12173 25143
rect 12173 25109 12207 25143
rect 12207 25109 12216 25143
rect 12164 25100 12216 25109
rect 13452 25100 13504 25152
rect 15568 25168 15620 25220
rect 19892 25168 19944 25220
rect 25504 25347 25556 25356
rect 25504 25313 25513 25347
rect 25513 25313 25547 25347
rect 25547 25313 25556 25347
rect 26516 25372 26568 25424
rect 25504 25304 25556 25313
rect 28264 25449 28273 25483
rect 28273 25449 28307 25483
rect 28307 25449 28316 25483
rect 28264 25440 28316 25449
rect 31208 25440 31260 25492
rect 32312 25483 32364 25492
rect 32312 25449 32321 25483
rect 32321 25449 32355 25483
rect 32355 25449 32364 25483
rect 32312 25440 32364 25449
rect 34336 25483 34388 25492
rect 34336 25449 34345 25483
rect 34345 25449 34379 25483
rect 34379 25449 34388 25483
rect 34336 25440 34388 25449
rect 34428 25440 34480 25492
rect 29920 25372 29972 25424
rect 30564 25372 30616 25424
rect 26792 25236 26844 25288
rect 27988 25304 28040 25356
rect 26516 25168 26568 25220
rect 28724 25236 28776 25288
rect 29276 25304 29328 25356
rect 30472 25347 30524 25356
rect 30472 25313 30481 25347
rect 30481 25313 30515 25347
rect 30515 25313 30524 25347
rect 30472 25304 30524 25313
rect 30932 25304 30984 25356
rect 31300 25347 31352 25356
rect 31300 25313 31309 25347
rect 31309 25313 31343 25347
rect 31343 25313 31352 25347
rect 31300 25304 31352 25313
rect 31852 25304 31904 25356
rect 32404 25304 32456 25356
rect 30380 25236 30432 25288
rect 32588 25279 32640 25288
rect 31300 25168 31352 25220
rect 31760 25168 31812 25220
rect 16120 25100 16172 25152
rect 16856 25100 16908 25152
rect 17408 25143 17460 25152
rect 17408 25109 17417 25143
rect 17417 25109 17451 25143
rect 17451 25109 17460 25143
rect 17408 25100 17460 25109
rect 17500 25100 17552 25152
rect 22100 25100 22152 25152
rect 25780 25100 25832 25152
rect 26056 25100 26108 25152
rect 27988 25100 28040 25152
rect 29368 25100 29420 25152
rect 32036 25100 32088 25152
rect 32588 25245 32597 25279
rect 32597 25245 32631 25279
rect 32631 25245 32640 25279
rect 32588 25236 32640 25245
rect 32680 25279 32732 25288
rect 32680 25245 32689 25279
rect 32689 25245 32723 25279
rect 32723 25245 32732 25279
rect 32680 25236 32732 25245
rect 33140 25304 33192 25356
rect 33692 25304 33744 25356
rect 33968 25347 34020 25356
rect 33968 25313 33977 25347
rect 33977 25313 34011 25347
rect 34011 25313 34020 25347
rect 33968 25304 34020 25313
rect 34060 25347 34112 25356
rect 34060 25313 34069 25347
rect 34069 25313 34103 25347
rect 34103 25313 34112 25347
rect 34060 25304 34112 25313
rect 34244 25304 34296 25356
rect 36452 25347 36504 25356
rect 36452 25313 36461 25347
rect 36461 25313 36495 25347
rect 36495 25313 36504 25347
rect 36452 25304 36504 25313
rect 36544 25347 36596 25356
rect 36544 25313 36553 25347
rect 36553 25313 36587 25347
rect 36587 25313 36596 25347
rect 36544 25304 36596 25313
rect 37096 25304 37148 25356
rect 55588 25440 55640 25492
rect 57980 25483 58032 25492
rect 57980 25449 57989 25483
rect 57989 25449 58023 25483
rect 58023 25449 58032 25483
rect 57980 25440 58032 25449
rect 56324 25372 56376 25424
rect 36728 25279 36780 25288
rect 36728 25245 36737 25279
rect 36737 25245 36771 25279
rect 36771 25245 36780 25279
rect 36728 25236 36780 25245
rect 36084 25168 36136 25220
rect 55680 25304 55732 25356
rect 57428 25304 57480 25356
rect 34612 25100 34664 25152
rect 35900 25100 35952 25152
rect 55404 25143 55456 25152
rect 55404 25109 55413 25143
rect 55413 25109 55447 25143
rect 55447 25109 55456 25143
rect 55404 25100 55456 25109
rect 57244 25143 57296 25152
rect 57244 25109 57253 25143
rect 57253 25109 57287 25143
rect 57287 25109 57296 25143
rect 57244 25100 57296 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 1860 24896 1912 24948
rect 3332 24760 3384 24812
rect 4068 24828 4120 24880
rect 8300 24828 8352 24880
rect 9588 24896 9640 24948
rect 13452 24896 13504 24948
rect 13636 24939 13688 24948
rect 13636 24905 13645 24939
rect 13645 24905 13679 24939
rect 13679 24905 13688 24939
rect 13636 24896 13688 24905
rect 14556 24896 14608 24948
rect 11520 24828 11572 24880
rect 12164 24828 12216 24880
rect 15660 24896 15712 24948
rect 16764 24896 16816 24948
rect 17408 24896 17460 24948
rect 21088 24896 21140 24948
rect 24584 24896 24636 24948
rect 17592 24828 17644 24880
rect 17960 24828 18012 24880
rect 18328 24828 18380 24880
rect 20168 24828 20220 24880
rect 24492 24828 24544 24880
rect 3148 24692 3200 24744
rect 4988 24692 5040 24744
rect 5264 24692 5316 24744
rect 5632 24692 5684 24744
rect 10968 24760 11020 24812
rect 12072 24760 12124 24812
rect 14464 24760 14516 24812
rect 16672 24760 16724 24812
rect 18144 24760 18196 24812
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 21824 24760 21876 24812
rect 22468 24760 22520 24812
rect 26148 24896 26200 24948
rect 26884 24939 26936 24948
rect 26884 24905 26893 24939
rect 26893 24905 26927 24939
rect 26927 24905 26936 24939
rect 26884 24896 26936 24905
rect 30380 24896 30432 24948
rect 32036 24939 32088 24948
rect 32036 24905 32045 24939
rect 32045 24905 32079 24939
rect 32079 24905 32088 24939
rect 32036 24896 32088 24905
rect 32680 24896 32732 24948
rect 27804 24760 27856 24812
rect 8208 24692 8260 24744
rect 6092 24624 6144 24676
rect 7932 24624 7984 24676
rect 8484 24692 8536 24744
rect 10140 24735 10192 24744
rect 10140 24701 10149 24735
rect 10149 24701 10183 24735
rect 10183 24701 10192 24735
rect 10140 24692 10192 24701
rect 10416 24735 10468 24744
rect 10416 24701 10425 24735
rect 10425 24701 10459 24735
rect 10459 24701 10468 24735
rect 10692 24735 10744 24744
rect 10416 24692 10468 24701
rect 10692 24701 10701 24735
rect 10701 24701 10735 24735
rect 10735 24701 10744 24735
rect 10692 24692 10744 24701
rect 12808 24692 12860 24744
rect 11152 24624 11204 24676
rect 11520 24624 11572 24676
rect 11796 24624 11848 24676
rect 14372 24692 14424 24744
rect 15844 24692 15896 24744
rect 16856 24692 16908 24744
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 12992 24624 13044 24676
rect 14740 24624 14792 24676
rect 17132 24624 17184 24676
rect 18604 24735 18656 24744
rect 3884 24599 3936 24608
rect 3884 24565 3893 24599
rect 3893 24565 3927 24599
rect 3927 24565 3936 24599
rect 3884 24556 3936 24565
rect 4804 24599 4856 24608
rect 4804 24565 4813 24599
rect 4813 24565 4847 24599
rect 4847 24565 4856 24599
rect 4804 24556 4856 24565
rect 5264 24556 5316 24608
rect 7104 24556 7156 24608
rect 8024 24556 8076 24608
rect 8300 24556 8352 24608
rect 8576 24556 8628 24608
rect 9680 24556 9732 24608
rect 10876 24599 10928 24608
rect 10876 24565 10885 24599
rect 10885 24565 10919 24599
rect 10919 24565 10928 24599
rect 10876 24556 10928 24565
rect 13452 24556 13504 24608
rect 14004 24556 14056 24608
rect 14648 24556 14700 24608
rect 17776 24556 17828 24608
rect 18604 24701 18638 24735
rect 18638 24701 18656 24735
rect 18604 24692 18656 24701
rect 20812 24692 20864 24744
rect 21456 24692 21508 24744
rect 21732 24692 21784 24744
rect 25504 24735 25556 24744
rect 18696 24624 18748 24676
rect 18788 24556 18840 24608
rect 20076 24556 20128 24608
rect 20996 24624 21048 24676
rect 22008 24624 22060 24676
rect 23388 24667 23440 24676
rect 23388 24633 23397 24667
rect 23397 24633 23431 24667
rect 23431 24633 23440 24667
rect 23388 24624 23440 24633
rect 24584 24624 24636 24676
rect 25504 24701 25513 24735
rect 25513 24701 25547 24735
rect 25547 24701 25556 24735
rect 25504 24692 25556 24701
rect 25780 24735 25832 24744
rect 25780 24701 25814 24735
rect 25814 24701 25832 24735
rect 25780 24692 25832 24701
rect 31300 24760 31352 24812
rect 31668 24760 31720 24812
rect 24400 24556 24452 24608
rect 26148 24624 26200 24676
rect 29368 24735 29420 24744
rect 29368 24701 29402 24735
rect 29402 24701 29420 24735
rect 29368 24692 29420 24701
rect 29736 24692 29788 24744
rect 32588 24692 32640 24744
rect 33324 24828 33376 24880
rect 35992 24896 36044 24948
rect 33968 24760 34020 24812
rect 55404 24760 55456 24812
rect 33692 24692 33744 24744
rect 34428 24692 34480 24744
rect 34704 24692 34756 24744
rect 35900 24692 35952 24744
rect 36452 24735 36504 24744
rect 36452 24701 36461 24735
rect 36461 24701 36495 24735
rect 36495 24701 36504 24735
rect 36452 24692 36504 24701
rect 36636 24735 36688 24744
rect 36636 24701 36645 24735
rect 36645 24701 36679 24735
rect 36679 24701 36688 24735
rect 36636 24692 36688 24701
rect 36728 24692 36780 24744
rect 55772 24735 55824 24744
rect 27988 24599 28040 24608
rect 27988 24565 27997 24599
rect 27997 24565 28031 24599
rect 28031 24565 28040 24599
rect 27988 24556 28040 24565
rect 30840 24556 30892 24608
rect 31392 24556 31444 24608
rect 32404 24624 32456 24676
rect 33324 24624 33376 24676
rect 32680 24556 32732 24608
rect 55772 24701 55781 24735
rect 55781 24701 55815 24735
rect 55815 24701 55824 24735
rect 55772 24692 55824 24701
rect 58072 24760 58124 24812
rect 57060 24735 57112 24744
rect 57060 24701 57069 24735
rect 57069 24701 57103 24735
rect 57103 24701 57112 24735
rect 57060 24692 57112 24701
rect 57428 24692 57480 24744
rect 35808 24556 35860 24608
rect 57336 24624 57388 24676
rect 57980 24556 58032 24608
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 50326 24454 50378 24506
rect 50390 24454 50442 24506
rect 50454 24454 50506 24506
rect 50518 24454 50570 24506
rect 5080 24352 5132 24404
rect 5632 24395 5684 24404
rect 5632 24361 5641 24395
rect 5641 24361 5675 24395
rect 5675 24361 5684 24395
rect 5632 24352 5684 24361
rect 6092 24395 6144 24404
rect 6092 24361 6101 24395
rect 6101 24361 6135 24395
rect 6135 24361 6144 24395
rect 6092 24352 6144 24361
rect 6368 24352 6420 24404
rect 8484 24395 8536 24404
rect 4804 24284 4856 24336
rect 5264 24284 5316 24336
rect 3884 24216 3936 24268
rect 2688 24191 2740 24200
rect 2688 24157 2697 24191
rect 2697 24157 2731 24191
rect 2731 24157 2740 24191
rect 2688 24148 2740 24157
rect 4068 24148 4120 24200
rect 6368 24259 6420 24268
rect 6368 24225 6377 24259
rect 6377 24225 6411 24259
rect 6411 24225 6420 24259
rect 8484 24361 8493 24395
rect 8493 24361 8527 24395
rect 8527 24361 8536 24395
rect 8484 24352 8536 24361
rect 10416 24352 10468 24404
rect 14464 24352 14516 24404
rect 6368 24216 6420 24225
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 7564 24259 7616 24268
rect 7564 24225 7573 24259
rect 7573 24225 7607 24259
rect 7607 24225 7616 24259
rect 7564 24216 7616 24225
rect 8024 24216 8076 24268
rect 8300 24216 8352 24268
rect 9588 24284 9640 24336
rect 10876 24284 10928 24336
rect 10968 24284 11020 24336
rect 10784 24216 10836 24268
rect 11336 24259 11388 24268
rect 11336 24225 11345 24259
rect 11345 24225 11379 24259
rect 11379 24225 11388 24259
rect 11336 24216 11388 24225
rect 11520 24259 11572 24268
rect 11520 24225 11529 24259
rect 11529 24225 11563 24259
rect 11563 24225 11572 24259
rect 11520 24216 11572 24225
rect 12440 24284 12492 24336
rect 16764 24284 16816 24336
rect 11980 24216 12032 24268
rect 12624 24216 12676 24268
rect 14464 24216 14516 24268
rect 14832 24259 14884 24268
rect 14832 24225 14841 24259
rect 14841 24225 14875 24259
rect 14875 24225 14884 24259
rect 14832 24216 14884 24225
rect 14924 24216 14976 24268
rect 24400 24352 24452 24404
rect 29552 24395 29604 24404
rect 29552 24361 29561 24395
rect 29561 24361 29595 24395
rect 29595 24361 29604 24395
rect 29552 24352 29604 24361
rect 30472 24352 30524 24404
rect 31668 24352 31720 24404
rect 32588 24352 32640 24404
rect 35992 24352 36044 24404
rect 55772 24352 55824 24404
rect 19064 24327 19116 24336
rect 19064 24293 19073 24327
rect 19073 24293 19107 24327
rect 19107 24293 19116 24327
rect 19064 24284 19116 24293
rect 11612 24191 11664 24200
rect 3056 24080 3108 24132
rect 7932 24080 7984 24132
rect 8668 24080 8720 24132
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 12348 24148 12400 24200
rect 14188 24148 14240 24200
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 17960 24259 18012 24268
rect 17960 24225 17969 24259
rect 17969 24225 18003 24259
rect 18003 24225 18012 24259
rect 17960 24216 18012 24225
rect 18236 24216 18288 24268
rect 18604 24216 18656 24268
rect 21180 24284 21232 24336
rect 21824 24284 21876 24336
rect 21916 24284 21968 24336
rect 29092 24284 29144 24336
rect 57980 24327 58032 24336
rect 57980 24293 57989 24327
rect 57989 24293 58023 24327
rect 58023 24293 58032 24327
rect 57980 24284 58032 24293
rect 58164 24327 58216 24336
rect 58164 24293 58173 24327
rect 58173 24293 58207 24327
rect 58207 24293 58216 24327
rect 58164 24284 58216 24293
rect 18052 24191 18104 24200
rect 1860 24055 1912 24064
rect 1860 24021 1869 24055
rect 1869 24021 1903 24055
rect 1903 24021 1912 24055
rect 1860 24012 1912 24021
rect 1952 24012 2004 24064
rect 6552 24055 6604 24064
rect 6552 24021 6561 24055
rect 6561 24021 6595 24055
rect 6595 24021 6604 24055
rect 6552 24012 6604 24021
rect 6920 24012 6972 24064
rect 8392 24012 8444 24064
rect 10692 24012 10744 24064
rect 13452 24055 13504 24064
rect 13452 24021 13461 24055
rect 13461 24021 13495 24055
rect 13495 24021 13504 24055
rect 13452 24012 13504 24021
rect 13544 24012 13596 24064
rect 17592 24080 17644 24132
rect 17316 24012 17368 24064
rect 18052 24157 18061 24191
rect 18061 24157 18095 24191
rect 18095 24157 18104 24191
rect 18052 24148 18104 24157
rect 20628 24216 20680 24268
rect 22652 24216 22704 24268
rect 22836 24216 22888 24268
rect 25412 24216 25464 24268
rect 25688 24259 25740 24268
rect 25688 24225 25697 24259
rect 25697 24225 25731 24259
rect 25731 24225 25740 24259
rect 25688 24216 25740 24225
rect 20352 24191 20404 24200
rect 20352 24157 20361 24191
rect 20361 24157 20395 24191
rect 20395 24157 20404 24191
rect 20352 24148 20404 24157
rect 27344 24216 27396 24268
rect 30748 24216 30800 24268
rect 17960 24080 18012 24132
rect 21916 24080 21968 24132
rect 22008 24080 22060 24132
rect 26516 24148 26568 24200
rect 28356 24148 28408 24200
rect 28908 24191 28960 24200
rect 28908 24157 28917 24191
rect 28917 24157 28951 24191
rect 28951 24157 28960 24191
rect 28908 24148 28960 24157
rect 30288 24148 30340 24200
rect 30840 24148 30892 24200
rect 32036 24216 32088 24268
rect 32404 24259 32456 24268
rect 32404 24225 32413 24259
rect 32413 24225 32447 24259
rect 32447 24225 32456 24259
rect 32404 24216 32456 24225
rect 32680 24216 32732 24268
rect 33140 24216 33192 24268
rect 35808 24259 35860 24268
rect 35808 24225 35817 24259
rect 35817 24225 35851 24259
rect 35851 24225 35860 24259
rect 35808 24216 35860 24225
rect 55680 24259 55732 24268
rect 55680 24225 55689 24259
rect 55689 24225 55723 24259
rect 55723 24225 55732 24259
rect 55680 24216 55732 24225
rect 57428 24259 57480 24268
rect 57428 24225 57437 24259
rect 57437 24225 57471 24259
rect 57471 24225 57480 24259
rect 57428 24216 57480 24225
rect 31024 24080 31076 24132
rect 31484 24148 31536 24200
rect 31760 24148 31812 24200
rect 20168 24012 20220 24064
rect 20536 24012 20588 24064
rect 20904 24012 20956 24064
rect 23112 24012 23164 24064
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 25136 24012 25188 24064
rect 28448 24055 28500 24064
rect 28448 24021 28457 24055
rect 28457 24021 28491 24055
rect 28491 24021 28500 24055
rect 28448 24012 28500 24021
rect 30840 24055 30892 24064
rect 30840 24021 30849 24055
rect 30849 24021 30883 24055
rect 30883 24021 30892 24055
rect 30840 24012 30892 24021
rect 34704 24080 34756 24132
rect 34152 24012 34204 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 6552 23808 6604 23860
rect 6828 23808 6880 23860
rect 8668 23808 8720 23860
rect 8852 23851 8904 23860
rect 8852 23817 8861 23851
rect 8861 23817 8895 23851
rect 8895 23817 8904 23851
rect 8852 23808 8904 23817
rect 9128 23808 9180 23860
rect 9864 23808 9916 23860
rect 2964 23740 3016 23792
rect 2872 23672 2924 23724
rect 4620 23672 4672 23724
rect 1952 23604 2004 23656
rect 4436 23604 4488 23656
rect 4988 23604 5040 23656
rect 6000 23672 6052 23724
rect 6368 23672 6420 23724
rect 8208 23740 8260 23792
rect 11980 23808 12032 23860
rect 14004 23851 14056 23860
rect 14004 23817 14013 23851
rect 14013 23817 14047 23851
rect 14047 23817 14056 23851
rect 14004 23808 14056 23817
rect 14832 23808 14884 23860
rect 17040 23808 17092 23860
rect 20352 23851 20404 23860
rect 20352 23817 20361 23851
rect 20361 23817 20395 23851
rect 20395 23817 20404 23851
rect 20352 23808 20404 23817
rect 11244 23740 11296 23792
rect 11888 23740 11940 23792
rect 23388 23808 23440 23860
rect 23572 23808 23624 23860
rect 26148 23808 26200 23860
rect 29368 23808 29420 23860
rect 29736 23808 29788 23860
rect 30564 23808 30616 23860
rect 32220 23808 32272 23860
rect 33140 23808 33192 23860
rect 5908 23647 5960 23656
rect 5908 23613 5917 23647
rect 5917 23613 5951 23647
rect 5951 23613 5960 23647
rect 5908 23604 5960 23613
rect 6828 23647 6880 23656
rect 6828 23613 6837 23647
rect 6837 23613 6871 23647
rect 6871 23613 6880 23647
rect 6828 23604 6880 23613
rect 11980 23672 12032 23724
rect 21548 23740 21600 23792
rect 23296 23740 23348 23792
rect 26516 23740 26568 23792
rect 30932 23740 30984 23792
rect 36636 23808 36688 23860
rect 56048 23851 56100 23860
rect 56048 23817 56057 23851
rect 56057 23817 56091 23851
rect 56091 23817 56100 23851
rect 56048 23808 56100 23817
rect 14188 23715 14240 23724
rect 8484 23604 8536 23656
rect 9680 23604 9732 23656
rect 12072 23647 12124 23656
rect 12072 23613 12081 23647
rect 12081 23613 12115 23647
rect 12115 23613 12124 23647
rect 12348 23647 12400 23656
rect 12072 23604 12124 23613
rect 12348 23613 12382 23647
rect 12382 23613 12400 23647
rect 12348 23604 12400 23613
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 15200 23715 15252 23724
rect 4528 23536 4580 23588
rect 7012 23536 7064 23588
rect 7564 23536 7616 23588
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 4804 23511 4856 23520
rect 2780 23468 2832 23477
rect 4804 23477 4813 23511
rect 4813 23477 4847 23511
rect 4847 23477 4856 23511
rect 4804 23468 4856 23477
rect 7840 23468 7892 23520
rect 14280 23604 14332 23656
rect 14924 23647 14976 23656
rect 14924 23613 14933 23647
rect 14933 23613 14967 23647
rect 14967 23613 14976 23647
rect 14924 23604 14976 23613
rect 15200 23681 15209 23715
rect 15209 23681 15243 23715
rect 15243 23681 15252 23715
rect 15200 23672 15252 23681
rect 15660 23604 15712 23656
rect 16212 23647 16264 23656
rect 16212 23613 16221 23647
rect 16221 23613 16255 23647
rect 16255 23613 16264 23647
rect 16212 23604 16264 23613
rect 16396 23647 16448 23656
rect 16396 23613 16405 23647
rect 16405 23613 16439 23647
rect 16439 23613 16448 23647
rect 16396 23604 16448 23613
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 20076 23647 20128 23656
rect 20076 23613 20085 23647
rect 20085 23613 20119 23647
rect 20119 23613 20128 23647
rect 20076 23604 20128 23613
rect 14464 23536 14516 23588
rect 14188 23511 14240 23520
rect 14188 23477 14197 23511
rect 14197 23477 14231 23511
rect 14231 23477 14240 23511
rect 14188 23468 14240 23477
rect 15384 23468 15436 23520
rect 18512 23511 18564 23520
rect 18512 23477 18521 23511
rect 18521 23477 18555 23511
rect 18555 23477 18564 23511
rect 18512 23468 18564 23477
rect 19432 23536 19484 23588
rect 20352 23536 20404 23588
rect 22192 23604 22244 23656
rect 22284 23604 22336 23656
rect 22836 23647 22888 23656
rect 22836 23613 22845 23647
rect 22845 23613 22879 23647
rect 22879 23613 22888 23647
rect 22836 23604 22888 23613
rect 23296 23604 23348 23656
rect 24216 23604 24268 23656
rect 26608 23672 26660 23724
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 30380 23672 30432 23724
rect 25504 23647 25556 23656
rect 25504 23613 25513 23647
rect 25513 23613 25547 23647
rect 25547 23613 25556 23647
rect 25504 23604 25556 23613
rect 26884 23604 26936 23656
rect 28448 23604 28500 23656
rect 30748 23604 30800 23656
rect 31024 23604 31076 23656
rect 31392 23647 31444 23656
rect 21456 23579 21508 23588
rect 21456 23545 21465 23579
rect 21465 23545 21499 23579
rect 21499 23545 21508 23579
rect 22652 23579 22704 23588
rect 21456 23536 21508 23545
rect 22652 23545 22661 23579
rect 22661 23545 22695 23579
rect 22695 23545 22704 23579
rect 22652 23536 22704 23545
rect 21640 23511 21692 23520
rect 21640 23477 21649 23511
rect 21649 23477 21683 23511
rect 21683 23477 21692 23511
rect 21640 23468 21692 23477
rect 21824 23468 21876 23520
rect 25320 23536 25372 23588
rect 25044 23468 25096 23520
rect 30012 23536 30064 23588
rect 30288 23579 30340 23588
rect 30288 23545 30297 23579
rect 30297 23545 30331 23579
rect 30331 23545 30340 23579
rect 30288 23536 30340 23545
rect 25964 23468 26016 23520
rect 27160 23468 27212 23520
rect 31024 23468 31076 23520
rect 31392 23613 31401 23647
rect 31401 23613 31435 23647
rect 31435 23613 31444 23647
rect 31392 23604 31444 23613
rect 34428 23740 34480 23792
rect 58164 23783 58216 23792
rect 58164 23749 58173 23783
rect 58173 23749 58207 23783
rect 58207 23749 58216 23783
rect 58164 23740 58216 23749
rect 34704 23672 34756 23724
rect 31944 23647 31996 23656
rect 31944 23613 31953 23647
rect 31953 23613 31987 23647
rect 31987 23613 31996 23647
rect 31944 23604 31996 23613
rect 33232 23604 33284 23656
rect 31576 23536 31628 23588
rect 33508 23647 33560 23656
rect 33508 23613 33517 23647
rect 33517 23613 33551 23647
rect 33551 23613 33560 23647
rect 33692 23647 33744 23656
rect 33508 23604 33560 23613
rect 33692 23613 33701 23647
rect 33701 23613 33735 23647
rect 33735 23613 33744 23647
rect 33692 23604 33744 23613
rect 33968 23604 34020 23656
rect 34244 23604 34296 23656
rect 35348 23604 35400 23656
rect 34060 23536 34112 23588
rect 35992 23536 36044 23588
rect 55588 23647 55640 23656
rect 55588 23613 55597 23647
rect 55597 23613 55631 23647
rect 55631 23613 55640 23647
rect 55588 23604 55640 23613
rect 56508 23604 56560 23656
rect 57336 23604 57388 23656
rect 58072 23536 58124 23588
rect 31392 23468 31444 23520
rect 31944 23468 31996 23520
rect 34520 23468 34572 23520
rect 36176 23511 36228 23520
rect 36176 23477 36185 23511
rect 36185 23477 36219 23511
rect 36219 23477 36228 23511
rect 36176 23468 36228 23477
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 55220 23511 55272 23520
rect 55220 23477 55229 23511
rect 55229 23477 55263 23511
rect 55263 23477 55272 23511
rect 55220 23468 55272 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 50326 23366 50378 23418
rect 50390 23366 50442 23418
rect 50454 23366 50506 23418
rect 50518 23366 50570 23418
rect 3148 23307 3200 23316
rect 3148 23273 3157 23307
rect 3157 23273 3191 23307
rect 3191 23273 3200 23307
rect 3148 23264 3200 23273
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 10140 23264 10192 23316
rect 10968 23264 11020 23316
rect 11152 23264 11204 23316
rect 54300 23264 54352 23316
rect 55588 23264 55640 23316
rect 1860 23239 1912 23248
rect 1860 23205 1869 23239
rect 1869 23205 1903 23239
rect 1903 23205 1912 23239
rect 1860 23196 1912 23205
rect 4804 23196 4856 23248
rect 2596 23128 2648 23180
rect 3424 23128 3476 23180
rect 4068 23128 4120 23180
rect 6920 23171 6972 23180
rect 6920 23137 6929 23171
rect 6929 23137 6963 23171
rect 6963 23137 6972 23171
rect 6920 23128 6972 23137
rect 7196 23128 7248 23180
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 9680 23128 9732 23180
rect 10324 23128 10376 23180
rect 11152 23171 11204 23180
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 12072 23196 12124 23248
rect 14556 23196 14608 23248
rect 11520 23171 11572 23180
rect 11520 23137 11529 23171
rect 11529 23137 11563 23171
rect 11563 23137 11572 23171
rect 11520 23128 11572 23137
rect 11796 23128 11848 23180
rect 12348 23128 12400 23180
rect 16212 23196 16264 23248
rect 7932 23060 7984 23112
rect 11704 23060 11756 23112
rect 14096 23060 14148 23112
rect 1952 22967 2004 22976
rect 1952 22933 1961 22967
rect 1961 22933 1995 22967
rect 1995 22933 2004 22967
rect 1952 22924 2004 22933
rect 5724 22924 5776 22976
rect 8024 22924 8076 22976
rect 8576 22924 8628 22976
rect 11244 22924 11296 22976
rect 12164 22924 12216 22976
rect 14004 22924 14056 22976
rect 15292 23128 15344 23180
rect 17040 23171 17092 23180
rect 17040 23137 17049 23171
rect 17049 23137 17083 23171
rect 17083 23137 17092 23171
rect 17040 23128 17092 23137
rect 17776 23128 17828 23180
rect 18512 23196 18564 23248
rect 20076 23128 20128 23180
rect 20168 23171 20220 23180
rect 20168 23137 20177 23171
rect 20177 23137 20211 23171
rect 20211 23137 20220 23171
rect 20168 23128 20220 23137
rect 20720 23128 20772 23180
rect 21732 23128 21784 23180
rect 16120 22967 16172 22976
rect 16120 22933 16129 22967
rect 16129 22933 16163 22967
rect 16163 22933 16172 22967
rect 16120 22924 16172 22933
rect 17040 22924 17092 22976
rect 19984 23060 20036 23112
rect 20444 23103 20496 23112
rect 20444 23069 20470 23103
rect 20470 23069 20496 23103
rect 20444 23060 20496 23069
rect 21548 23060 21600 23112
rect 24860 23196 24912 23248
rect 25872 23196 25924 23248
rect 26332 23196 26384 23248
rect 22836 23128 22888 23180
rect 23848 23171 23900 23180
rect 23848 23137 23857 23171
rect 23857 23137 23891 23171
rect 23891 23137 23900 23171
rect 23848 23128 23900 23137
rect 24216 23128 24268 23180
rect 24308 23171 24360 23180
rect 24308 23137 24317 23171
rect 24317 23137 24351 23171
rect 24351 23137 24360 23171
rect 24308 23128 24360 23137
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 18788 22992 18840 23044
rect 26516 23128 26568 23180
rect 28816 23128 28868 23180
rect 25596 23060 25648 23112
rect 30840 23196 30892 23248
rect 31760 23239 31812 23248
rect 31760 23205 31769 23239
rect 31769 23205 31803 23239
rect 31803 23205 31812 23239
rect 31760 23196 31812 23205
rect 29460 23128 29512 23180
rect 31024 23171 31076 23180
rect 31024 23137 31033 23171
rect 31033 23137 31067 23171
rect 31067 23137 31076 23171
rect 31024 23128 31076 23137
rect 31208 23171 31260 23180
rect 31208 23137 31217 23171
rect 31217 23137 31251 23171
rect 31251 23137 31260 23171
rect 31208 23128 31260 23137
rect 31576 23171 31628 23180
rect 31576 23137 31585 23171
rect 31585 23137 31619 23171
rect 31619 23137 31628 23171
rect 31576 23128 31628 23137
rect 32220 23171 32272 23180
rect 32220 23137 32229 23171
rect 32229 23137 32263 23171
rect 32263 23137 32272 23171
rect 32220 23128 32272 23137
rect 32404 23171 32456 23180
rect 32404 23137 32411 23171
rect 32411 23137 32456 23171
rect 32404 23128 32456 23137
rect 27344 23035 27396 23044
rect 27344 23001 27353 23035
rect 27353 23001 27387 23035
rect 27387 23001 27396 23035
rect 27344 22992 27396 23001
rect 29276 23060 29328 23112
rect 30380 23060 30432 23112
rect 31300 23103 31352 23112
rect 31300 23069 31309 23103
rect 31309 23069 31343 23103
rect 31343 23069 31352 23103
rect 31300 23060 31352 23069
rect 31392 23103 31444 23112
rect 31392 23069 31401 23103
rect 31401 23069 31435 23103
rect 31435 23069 31444 23103
rect 31392 23060 31444 23069
rect 31760 23060 31812 23112
rect 34152 23171 34204 23180
rect 34152 23137 34161 23171
rect 34161 23137 34195 23171
rect 34195 23137 34204 23171
rect 34152 23128 34204 23137
rect 34520 23171 34572 23180
rect 34520 23137 34529 23171
rect 34529 23137 34563 23171
rect 34563 23137 34572 23171
rect 34520 23128 34572 23137
rect 36176 23196 36228 23248
rect 36544 23128 36596 23180
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 19156 22924 19208 22976
rect 21364 22924 21416 22976
rect 24216 22924 24268 22976
rect 25688 22924 25740 22976
rect 26884 22924 26936 22976
rect 28264 22924 28316 22976
rect 29552 22992 29604 23044
rect 32312 22924 32364 22976
rect 36728 23060 36780 23112
rect 33692 22992 33744 23044
rect 34428 23035 34480 23044
rect 34428 23001 34437 23035
rect 34437 23001 34471 23035
rect 34471 23001 34480 23035
rect 34428 22992 34480 23001
rect 36544 22992 36596 23044
rect 55404 23128 55456 23180
rect 57980 23171 58032 23180
rect 57980 23137 57989 23171
rect 57989 23137 58023 23171
rect 58023 23137 58032 23171
rect 57980 23128 58032 23137
rect 55680 22992 55732 23044
rect 58164 23035 58216 23044
rect 58164 23001 58173 23035
rect 58173 23001 58207 23035
rect 58207 23001 58216 23035
rect 58164 22992 58216 23001
rect 57520 22924 57572 22976
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 2136 22695 2188 22704
rect 2136 22661 2145 22695
rect 2145 22661 2179 22695
rect 2179 22661 2188 22695
rect 2136 22652 2188 22661
rect 6920 22720 6972 22772
rect 2872 22652 2924 22704
rect 4896 22584 4948 22636
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 2044 22516 2096 22568
rect 3516 22559 3568 22568
rect 3516 22525 3525 22559
rect 3525 22525 3559 22559
rect 3559 22525 3568 22559
rect 3516 22516 3568 22525
rect 5724 22559 5776 22568
rect 5724 22525 5733 22559
rect 5733 22525 5767 22559
rect 5767 22525 5776 22559
rect 5724 22516 5776 22525
rect 7472 22559 7524 22568
rect 7472 22525 7481 22559
rect 7481 22525 7515 22559
rect 7515 22525 7524 22559
rect 7472 22516 7524 22525
rect 10508 22652 10560 22704
rect 14188 22720 14240 22772
rect 14004 22695 14056 22704
rect 14004 22661 14013 22695
rect 14013 22661 14047 22695
rect 14047 22661 14056 22695
rect 15660 22763 15712 22772
rect 15660 22729 15669 22763
rect 15669 22729 15703 22763
rect 15703 22729 15712 22763
rect 15660 22720 15712 22729
rect 19800 22720 19852 22772
rect 19984 22763 20036 22772
rect 19984 22729 19993 22763
rect 19993 22729 20027 22763
rect 20027 22729 20036 22763
rect 19984 22720 20036 22729
rect 20168 22720 20220 22772
rect 20352 22763 20404 22772
rect 20352 22729 20361 22763
rect 20361 22729 20395 22763
rect 20395 22729 20404 22763
rect 20352 22720 20404 22729
rect 21732 22720 21784 22772
rect 24032 22720 24084 22772
rect 24492 22720 24544 22772
rect 25872 22720 25924 22772
rect 28908 22720 28960 22772
rect 29000 22720 29052 22772
rect 14004 22652 14056 22661
rect 10968 22584 11020 22636
rect 11060 22584 11112 22636
rect 11612 22584 11664 22636
rect 14096 22584 14148 22636
rect 18696 22652 18748 22704
rect 18788 22652 18840 22704
rect 19340 22652 19392 22704
rect 19524 22695 19576 22704
rect 19524 22661 19533 22695
rect 19533 22661 19567 22695
rect 19567 22661 19576 22695
rect 19524 22652 19576 22661
rect 30932 22720 30984 22772
rect 31208 22763 31260 22772
rect 31208 22729 31217 22763
rect 31217 22729 31251 22763
rect 31251 22729 31260 22763
rect 31208 22720 31260 22729
rect 31392 22720 31444 22772
rect 32404 22720 32456 22772
rect 35348 22720 35400 22772
rect 35992 22763 36044 22772
rect 35992 22729 36001 22763
rect 36001 22729 36035 22763
rect 36035 22729 36044 22763
rect 35992 22720 36044 22729
rect 57980 22763 58032 22772
rect 57980 22729 57989 22763
rect 57989 22729 58023 22763
rect 58023 22729 58032 22763
rect 57980 22720 58032 22729
rect 10048 22516 10100 22568
rect 10324 22559 10376 22568
rect 10324 22525 10333 22559
rect 10333 22525 10367 22559
rect 10367 22525 10376 22559
rect 10324 22516 10376 22525
rect 10416 22516 10468 22568
rect 10784 22516 10836 22568
rect 11428 22516 11480 22568
rect 12164 22516 12216 22568
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 2596 22380 2648 22432
rect 4804 22448 4856 22500
rect 4988 22491 5040 22500
rect 4988 22457 4997 22491
rect 4997 22457 5031 22491
rect 5031 22457 5040 22491
rect 4988 22448 5040 22457
rect 5448 22448 5500 22500
rect 5908 22380 5960 22432
rect 6276 22380 6328 22432
rect 7288 22380 7340 22432
rect 8116 22380 8168 22432
rect 11704 22448 11756 22500
rect 16120 22516 16172 22568
rect 17408 22516 17460 22568
rect 19064 22584 19116 22636
rect 18972 22559 19024 22568
rect 16396 22448 16448 22500
rect 17960 22448 18012 22500
rect 11520 22380 11572 22432
rect 14188 22423 14240 22432
rect 14188 22389 14197 22423
rect 14197 22389 14231 22423
rect 14231 22389 14240 22423
rect 14188 22380 14240 22389
rect 14280 22380 14332 22432
rect 17684 22423 17736 22432
rect 17684 22389 17693 22423
rect 17693 22389 17727 22423
rect 17727 22389 17736 22423
rect 18604 22448 18656 22500
rect 18972 22525 18981 22559
rect 18981 22525 19015 22559
rect 19015 22525 19024 22559
rect 18972 22516 19024 22525
rect 19340 22559 19392 22568
rect 19340 22525 19349 22559
rect 19349 22525 19383 22559
rect 19383 22525 19392 22559
rect 19340 22516 19392 22525
rect 19524 22516 19576 22568
rect 20076 22516 20128 22568
rect 20444 22559 20496 22568
rect 20444 22525 20453 22559
rect 20453 22525 20487 22559
rect 20487 22525 20496 22559
rect 20444 22516 20496 22525
rect 20996 22559 21048 22568
rect 20996 22525 21005 22559
rect 21005 22525 21039 22559
rect 21039 22525 21048 22559
rect 20996 22516 21048 22525
rect 21088 22559 21140 22568
rect 21088 22525 21098 22559
rect 21098 22525 21132 22559
rect 21132 22525 21140 22559
rect 21088 22516 21140 22525
rect 21456 22516 21508 22568
rect 21640 22516 21692 22568
rect 22652 22559 22704 22568
rect 22652 22525 22661 22559
rect 22661 22525 22695 22559
rect 22695 22525 22704 22559
rect 22652 22516 22704 22525
rect 23940 22559 23992 22568
rect 20352 22448 20404 22500
rect 21364 22491 21416 22500
rect 21364 22457 21373 22491
rect 21373 22457 21407 22491
rect 21407 22457 21416 22491
rect 23940 22525 23949 22559
rect 23949 22525 23983 22559
rect 23983 22525 23992 22559
rect 23940 22516 23992 22525
rect 24400 22516 24452 22568
rect 24584 22559 24636 22568
rect 24584 22525 24593 22559
rect 24593 22525 24627 22559
rect 24627 22525 24636 22559
rect 24584 22516 24636 22525
rect 24676 22559 24728 22568
rect 24676 22525 24686 22559
rect 24686 22525 24720 22559
rect 24720 22525 24728 22559
rect 24676 22516 24728 22525
rect 25780 22516 25832 22568
rect 25872 22516 25924 22568
rect 24860 22491 24912 22500
rect 21364 22448 21416 22457
rect 17684 22380 17736 22389
rect 18788 22380 18840 22432
rect 18972 22380 19024 22432
rect 20720 22380 20772 22432
rect 23848 22380 23900 22432
rect 24860 22457 24869 22491
rect 24869 22457 24903 22491
rect 24903 22457 24912 22491
rect 24860 22448 24912 22457
rect 24952 22491 25004 22500
rect 24952 22457 24961 22491
rect 24961 22457 24995 22491
rect 24995 22457 25004 22491
rect 24952 22448 25004 22457
rect 25136 22380 25188 22432
rect 25688 22423 25740 22432
rect 25688 22389 25697 22423
rect 25697 22389 25731 22423
rect 25731 22389 25740 22423
rect 25688 22380 25740 22389
rect 26148 22559 26200 22568
rect 26148 22525 26157 22559
rect 26157 22525 26191 22559
rect 26191 22525 26200 22559
rect 26424 22584 26476 22636
rect 26148 22516 26200 22525
rect 27344 22516 27396 22568
rect 28540 22516 28592 22568
rect 28632 22559 28684 22568
rect 28632 22525 28641 22559
rect 28641 22525 28675 22559
rect 28675 22525 28684 22559
rect 28632 22516 28684 22525
rect 29000 22516 29052 22568
rect 29276 22559 29328 22568
rect 29276 22525 29285 22559
rect 29285 22525 29319 22559
rect 29319 22525 29328 22559
rect 29276 22516 29328 22525
rect 29460 22559 29512 22568
rect 29460 22525 29469 22559
rect 29469 22525 29503 22559
rect 29503 22525 29512 22559
rect 29460 22516 29512 22525
rect 29368 22491 29420 22500
rect 29368 22457 29377 22491
rect 29377 22457 29411 22491
rect 29411 22457 29420 22491
rect 29368 22448 29420 22457
rect 27620 22380 27672 22432
rect 27896 22423 27948 22432
rect 27896 22389 27905 22423
rect 27905 22389 27939 22423
rect 27939 22389 27948 22423
rect 27896 22380 27948 22389
rect 30564 22584 30616 22636
rect 31576 22584 31628 22636
rect 34520 22652 34572 22704
rect 32220 22584 32272 22636
rect 33600 22584 33652 22636
rect 30288 22516 30340 22568
rect 31208 22516 31260 22568
rect 30380 22448 30432 22500
rect 31760 22448 31812 22500
rect 33232 22516 33284 22568
rect 34152 22559 34204 22568
rect 34152 22525 34161 22559
rect 34161 22525 34195 22559
rect 34195 22525 34204 22559
rect 34152 22516 34204 22525
rect 35348 22559 35400 22568
rect 35348 22525 35357 22559
rect 35357 22525 35391 22559
rect 35391 22525 35400 22559
rect 35348 22516 35400 22525
rect 35992 22559 36044 22568
rect 35992 22525 36001 22559
rect 36001 22525 36035 22559
rect 36035 22525 36044 22559
rect 35992 22516 36044 22525
rect 57520 22627 57572 22636
rect 57520 22593 57529 22627
rect 57529 22593 57563 22627
rect 57563 22593 57572 22627
rect 57520 22584 57572 22593
rect 55036 22559 55088 22568
rect 55036 22525 55045 22559
rect 55045 22525 55079 22559
rect 55079 22525 55088 22559
rect 55036 22516 55088 22525
rect 55496 22559 55548 22568
rect 55496 22525 55505 22559
rect 55505 22525 55539 22559
rect 55539 22525 55548 22559
rect 55496 22516 55548 22525
rect 56416 22516 56468 22568
rect 32404 22448 32456 22500
rect 34612 22448 34664 22500
rect 57060 22491 57112 22500
rect 57060 22457 57069 22491
rect 57069 22457 57103 22491
rect 57103 22457 57112 22491
rect 57060 22448 57112 22457
rect 31944 22380 31996 22432
rect 32036 22423 32088 22432
rect 32036 22389 32045 22423
rect 32045 22389 32079 22423
rect 32079 22389 32088 22423
rect 32036 22380 32088 22389
rect 32312 22380 32364 22432
rect 35440 22423 35492 22432
rect 35440 22389 35449 22423
rect 35449 22389 35483 22423
rect 35483 22389 35492 22423
rect 35440 22380 35492 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 50326 22278 50378 22330
rect 50390 22278 50442 22330
rect 50454 22278 50506 22330
rect 50518 22278 50570 22330
rect 10324 22176 10376 22228
rect 10968 22176 11020 22228
rect 6736 22108 6788 22160
rect 3424 22040 3476 22092
rect 5540 22083 5592 22092
rect 5540 22049 5549 22083
rect 5549 22049 5583 22083
rect 5583 22049 5592 22083
rect 5540 22040 5592 22049
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 6644 22083 6696 22092
rect 6644 22049 6653 22083
rect 6653 22049 6687 22083
rect 6687 22049 6696 22083
rect 6644 22040 6696 22049
rect 8208 22108 8260 22160
rect 7564 22083 7616 22092
rect 7564 22049 7573 22083
rect 7573 22049 7607 22083
rect 7607 22049 7616 22083
rect 7564 22040 7616 22049
rect 4068 21972 4120 22024
rect 9680 22040 9732 22092
rect 10048 22040 10100 22092
rect 10416 22108 10468 22160
rect 11152 22108 11204 22160
rect 13912 22176 13964 22228
rect 32220 22176 32272 22228
rect 11428 22151 11480 22160
rect 11428 22117 11437 22151
rect 11437 22117 11471 22151
rect 11471 22117 11480 22151
rect 11980 22151 12032 22160
rect 11428 22108 11480 22117
rect 11980 22117 11989 22151
rect 11989 22117 12023 22151
rect 12023 22117 12032 22151
rect 11980 22108 12032 22117
rect 10324 22083 10376 22092
rect 10324 22049 10333 22083
rect 10333 22049 10367 22083
rect 10367 22049 10376 22083
rect 10324 22040 10376 22049
rect 10508 22083 10560 22092
rect 10508 22049 10517 22083
rect 10517 22049 10551 22083
rect 10551 22049 10560 22083
rect 10508 22040 10560 22049
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 12072 22040 12124 22092
rect 12348 22040 12400 22092
rect 15016 22040 15068 22092
rect 15384 22040 15436 22092
rect 15844 22040 15896 22092
rect 18236 22083 18288 22092
rect 18236 22049 18245 22083
rect 18245 22049 18279 22083
rect 18279 22049 18288 22083
rect 18512 22083 18564 22092
rect 18236 22040 18288 22049
rect 18512 22049 18521 22083
rect 18521 22049 18555 22083
rect 18555 22049 18564 22083
rect 18512 22040 18564 22049
rect 3056 21947 3108 21956
rect 2320 21879 2372 21888
rect 2320 21845 2329 21879
rect 2329 21845 2363 21879
rect 2363 21845 2372 21879
rect 2320 21836 2372 21845
rect 3056 21913 3065 21947
rect 3065 21913 3099 21947
rect 3099 21913 3108 21947
rect 3056 21904 3108 21913
rect 4896 21947 4948 21956
rect 4896 21913 4905 21947
rect 4905 21913 4939 21947
rect 4939 21913 4948 21947
rect 4896 21904 4948 21913
rect 14188 21972 14240 22024
rect 15936 21972 15988 22024
rect 18328 21972 18380 22024
rect 11520 21904 11572 21956
rect 12440 21904 12492 21956
rect 12992 21904 13044 21956
rect 14280 21904 14332 21956
rect 15292 21904 15344 21956
rect 22192 22108 22244 22160
rect 23940 22151 23992 22160
rect 23940 22117 23949 22151
rect 23949 22117 23983 22151
rect 23983 22117 23992 22151
rect 23940 22108 23992 22117
rect 25136 22108 25188 22160
rect 25320 22151 25372 22160
rect 25320 22117 25329 22151
rect 25329 22117 25363 22151
rect 25363 22117 25372 22151
rect 25320 22108 25372 22117
rect 25688 22108 25740 22160
rect 20076 22083 20128 22092
rect 20076 22049 20085 22083
rect 20085 22049 20119 22083
rect 20119 22049 20128 22083
rect 20076 22040 20128 22049
rect 21824 22040 21876 22092
rect 22560 22083 22612 22092
rect 22560 22049 22569 22083
rect 22569 22049 22603 22083
rect 22603 22049 22612 22083
rect 22560 22040 22612 22049
rect 25228 22040 25280 22092
rect 25504 22083 25556 22092
rect 25504 22049 25513 22083
rect 25513 22049 25547 22083
rect 25547 22049 25556 22083
rect 25504 22040 25556 22049
rect 27896 22108 27948 22160
rect 30840 22108 30892 22160
rect 19708 21972 19760 22024
rect 20444 21972 20496 22024
rect 20720 21972 20772 22024
rect 22836 22015 22888 22024
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 25596 21972 25648 22024
rect 29184 22040 29236 22092
rect 30748 22083 30800 22092
rect 30748 22049 30757 22083
rect 30757 22049 30791 22083
rect 30791 22049 30800 22083
rect 30748 22040 30800 22049
rect 31392 22108 31444 22160
rect 32312 22151 32364 22160
rect 32312 22117 32321 22151
rect 32321 22117 32355 22151
rect 32355 22117 32364 22151
rect 32312 22108 32364 22117
rect 33232 22176 33284 22228
rect 33600 22176 33652 22228
rect 35440 22176 35492 22228
rect 38752 22176 38804 22228
rect 33324 22108 33376 22160
rect 27804 21972 27856 22024
rect 31300 22040 31352 22092
rect 32036 22083 32088 22092
rect 32036 22049 32045 22083
rect 32045 22049 32079 22083
rect 32079 22049 32088 22083
rect 32036 22040 32088 22049
rect 32220 22083 32272 22092
rect 32220 22049 32227 22083
rect 32227 22049 32272 22083
rect 32220 22040 32272 22049
rect 32496 22083 32548 22092
rect 32496 22049 32510 22083
rect 32510 22049 32544 22083
rect 32544 22049 32548 22083
rect 32496 22040 32548 22049
rect 33324 21972 33376 22024
rect 33692 22040 33744 22092
rect 33784 22083 33836 22092
rect 33784 22049 33793 22083
rect 33793 22049 33827 22083
rect 33827 22049 33836 22083
rect 33784 22040 33836 22049
rect 36084 22083 36136 22092
rect 36084 22049 36093 22083
rect 36093 22049 36127 22083
rect 36127 22049 36136 22083
rect 36084 22040 36136 22049
rect 36268 22083 36320 22092
rect 36268 22049 36277 22083
rect 36277 22049 36311 22083
rect 36311 22049 36320 22083
rect 36268 22040 36320 22049
rect 55220 22176 55272 22228
rect 39120 22108 39172 22160
rect 55496 22108 55548 22160
rect 23572 21904 23624 21956
rect 27620 21947 27672 21956
rect 27620 21913 27629 21947
rect 27629 21913 27663 21947
rect 27663 21913 27672 21947
rect 27620 21904 27672 21913
rect 31116 21947 31168 21956
rect 31116 21913 31125 21947
rect 31125 21913 31159 21947
rect 31159 21913 31168 21947
rect 31116 21904 31168 21913
rect 8208 21836 8260 21888
rect 8852 21836 8904 21888
rect 11980 21836 12032 21888
rect 15200 21836 15252 21888
rect 15384 21836 15436 21888
rect 16120 21836 16172 21888
rect 17500 21879 17552 21888
rect 17500 21845 17509 21879
rect 17509 21845 17543 21879
rect 17543 21845 17552 21879
rect 17500 21836 17552 21845
rect 17592 21836 17644 21888
rect 18144 21836 18196 21888
rect 20168 21836 20220 21888
rect 20352 21836 20404 21888
rect 20904 21836 20956 21888
rect 23020 21836 23072 21888
rect 24400 21836 24452 21888
rect 29092 21836 29144 21888
rect 29460 21836 29512 21888
rect 31300 21836 31352 21888
rect 32956 21836 33008 21888
rect 33140 21879 33192 21888
rect 33140 21845 33149 21879
rect 33149 21845 33183 21879
rect 33183 21845 33192 21879
rect 33140 21836 33192 21845
rect 35440 21904 35492 21956
rect 55036 22040 55088 22092
rect 55772 22083 55824 22092
rect 55772 22049 55781 22083
rect 55781 22049 55815 22083
rect 55815 22049 55824 22083
rect 55772 22040 55824 22049
rect 57980 22083 58032 22092
rect 57980 22049 57989 22083
rect 57989 22049 58023 22083
rect 58023 22049 58032 22083
rect 57980 22040 58032 22049
rect 48044 21972 48096 22024
rect 58072 21972 58124 22024
rect 58164 21947 58216 21956
rect 58164 21913 58173 21947
rect 58173 21913 58207 21947
rect 58207 21913 58216 21947
rect 58164 21904 58216 21913
rect 33784 21836 33836 21888
rect 34520 21836 34572 21888
rect 55864 21836 55916 21888
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 1952 21675 2004 21684
rect 1952 21641 1961 21675
rect 1961 21641 1995 21675
rect 1995 21641 2004 21675
rect 1952 21632 2004 21641
rect 2688 21632 2740 21684
rect 4804 21632 4856 21684
rect 5448 21632 5500 21684
rect 6736 21632 6788 21684
rect 15844 21632 15896 21684
rect 16120 21632 16172 21684
rect 6000 21564 6052 21616
rect 10600 21564 10652 21616
rect 3424 21496 3476 21548
rect 4068 21496 4120 21548
rect 2872 21360 2924 21412
rect 3424 21403 3476 21412
rect 3424 21369 3433 21403
rect 3433 21369 3467 21403
rect 3467 21369 3476 21403
rect 3424 21360 3476 21369
rect 4068 21403 4120 21412
rect 4068 21369 4077 21403
rect 4077 21369 4111 21403
rect 4111 21369 4120 21403
rect 4068 21360 4120 21369
rect 4804 21292 4856 21344
rect 6644 21496 6696 21548
rect 7564 21539 7616 21548
rect 7564 21505 7573 21539
rect 7573 21505 7607 21539
rect 7607 21505 7616 21539
rect 7564 21496 7616 21505
rect 8208 21496 8260 21548
rect 12440 21564 12492 21616
rect 13728 21496 13780 21548
rect 5632 21471 5684 21480
rect 5632 21437 5641 21471
rect 5641 21437 5675 21471
rect 5675 21437 5684 21471
rect 5632 21428 5684 21437
rect 6368 21428 6420 21480
rect 7932 21428 7984 21480
rect 8576 21471 8628 21480
rect 8576 21437 8585 21471
rect 8585 21437 8619 21471
rect 8619 21437 8628 21471
rect 8576 21428 8628 21437
rect 8852 21471 8904 21480
rect 8852 21437 8886 21471
rect 8886 21437 8904 21471
rect 8852 21428 8904 21437
rect 10140 21428 10192 21480
rect 7932 21335 7984 21344
rect 7932 21301 7941 21335
rect 7941 21301 7975 21335
rect 7975 21301 7984 21335
rect 7932 21292 7984 21301
rect 10324 21360 10376 21412
rect 10876 21428 10928 21480
rect 11336 21428 11388 21480
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 12440 21471 12492 21480
rect 12440 21437 12449 21471
rect 12449 21437 12483 21471
rect 12483 21437 12492 21471
rect 12440 21428 12492 21437
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 13544 21471 13596 21480
rect 13544 21437 13553 21471
rect 13553 21437 13587 21471
rect 13587 21437 13596 21471
rect 13544 21428 13596 21437
rect 13820 21428 13872 21480
rect 15200 21496 15252 21548
rect 15384 21496 15436 21548
rect 17960 21632 18012 21684
rect 18788 21632 18840 21684
rect 19340 21632 19392 21684
rect 20444 21632 20496 21684
rect 24032 21632 24084 21684
rect 24400 21632 24452 21684
rect 27252 21632 27304 21684
rect 27344 21632 27396 21684
rect 29000 21632 29052 21684
rect 31392 21632 31444 21684
rect 33232 21632 33284 21684
rect 33600 21675 33652 21684
rect 33600 21641 33609 21675
rect 33609 21641 33643 21675
rect 33643 21641 33652 21675
rect 33600 21632 33652 21641
rect 33692 21632 33744 21684
rect 35348 21632 35400 21684
rect 56416 21632 56468 21684
rect 57980 21675 58032 21684
rect 57980 21641 57989 21675
rect 57989 21641 58023 21675
rect 58023 21641 58032 21675
rect 57980 21632 58032 21641
rect 15016 21428 15068 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 15568 21471 15620 21480
rect 15568 21437 15577 21471
rect 15577 21437 15611 21471
rect 15611 21437 15620 21471
rect 15568 21428 15620 21437
rect 15844 21471 15896 21480
rect 15844 21437 15853 21471
rect 15853 21437 15887 21471
rect 15887 21437 15896 21471
rect 17776 21471 17828 21480
rect 15844 21428 15896 21437
rect 17776 21437 17785 21471
rect 17785 21437 17819 21471
rect 17819 21437 17828 21471
rect 17776 21428 17828 21437
rect 18328 21428 18380 21480
rect 12992 21360 13044 21412
rect 13728 21360 13780 21412
rect 10508 21292 10560 21344
rect 11152 21335 11204 21344
rect 11152 21301 11161 21335
rect 11161 21301 11195 21335
rect 11195 21301 11204 21335
rect 11152 21292 11204 21301
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 17040 21292 17092 21344
rect 22560 21564 22612 21616
rect 25228 21564 25280 21616
rect 19340 21496 19392 21548
rect 19708 21496 19760 21548
rect 23020 21496 23072 21548
rect 19984 21428 20036 21480
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 20628 21428 20680 21480
rect 20812 21471 20864 21480
rect 20812 21437 20821 21471
rect 20821 21437 20855 21471
rect 20855 21437 20864 21471
rect 20812 21428 20864 21437
rect 21364 21428 21416 21480
rect 22928 21471 22980 21480
rect 22928 21437 22937 21471
rect 22937 21437 22971 21471
rect 22971 21437 22980 21471
rect 22928 21428 22980 21437
rect 23112 21471 23164 21480
rect 23112 21437 23121 21471
rect 23121 21437 23155 21471
rect 23155 21437 23164 21471
rect 23112 21428 23164 21437
rect 23848 21496 23900 21548
rect 24400 21539 24452 21548
rect 24400 21505 24409 21539
rect 24409 21505 24443 21539
rect 24443 21505 24452 21539
rect 24400 21496 24452 21505
rect 23480 21471 23532 21480
rect 23480 21437 23489 21471
rect 23489 21437 23523 21471
rect 23523 21437 23532 21471
rect 23480 21428 23532 21437
rect 24216 21428 24268 21480
rect 25136 21471 25188 21480
rect 25136 21437 25145 21471
rect 25145 21437 25179 21471
rect 25179 21437 25188 21471
rect 25136 21428 25188 21437
rect 26700 21496 26752 21548
rect 30748 21496 30800 21548
rect 20260 21360 20312 21412
rect 24860 21360 24912 21412
rect 25412 21360 25464 21412
rect 26792 21471 26844 21480
rect 26792 21437 26813 21471
rect 26813 21437 26844 21471
rect 26792 21428 26844 21437
rect 27068 21428 27120 21480
rect 27620 21428 27672 21480
rect 26976 21360 27028 21412
rect 28540 21428 28592 21480
rect 29092 21471 29144 21480
rect 29092 21437 29101 21471
rect 29101 21437 29135 21471
rect 29135 21437 29144 21471
rect 29092 21428 29144 21437
rect 30564 21471 30616 21480
rect 29000 21360 29052 21412
rect 30564 21437 30573 21471
rect 30573 21437 30607 21471
rect 30607 21437 30616 21471
rect 30564 21428 30616 21437
rect 30656 21471 30708 21480
rect 30656 21437 30665 21471
rect 30665 21437 30699 21471
rect 30699 21437 30708 21471
rect 30656 21428 30708 21437
rect 19984 21292 20036 21344
rect 20076 21292 20128 21344
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 24400 21335 24452 21344
rect 24400 21301 24409 21335
rect 24409 21301 24443 21335
rect 24443 21301 24452 21335
rect 24400 21292 24452 21301
rect 25504 21335 25556 21344
rect 25504 21301 25513 21335
rect 25513 21301 25547 21335
rect 25547 21301 25556 21335
rect 25504 21292 25556 21301
rect 26608 21292 26660 21344
rect 26884 21292 26936 21344
rect 27252 21292 27304 21344
rect 29092 21292 29144 21344
rect 30380 21335 30432 21344
rect 30380 21301 30389 21335
rect 30389 21301 30423 21335
rect 30423 21301 30432 21335
rect 30380 21292 30432 21301
rect 30932 21564 30984 21616
rect 31484 21496 31536 21548
rect 32220 21564 32272 21616
rect 34152 21564 34204 21616
rect 58256 21564 58308 21616
rect 55864 21539 55916 21548
rect 31208 21428 31260 21480
rect 33324 21471 33376 21480
rect 33324 21437 33333 21471
rect 33333 21437 33367 21471
rect 33367 21437 33376 21471
rect 33324 21428 33376 21437
rect 33600 21428 33652 21480
rect 33876 21428 33928 21480
rect 55864 21505 55873 21539
rect 55873 21505 55907 21539
rect 55907 21505 55916 21539
rect 55864 21496 55916 21505
rect 36084 21471 36136 21480
rect 31484 21403 31536 21412
rect 31484 21369 31493 21403
rect 31493 21369 31527 21403
rect 31527 21369 31536 21403
rect 31484 21360 31536 21369
rect 33048 21360 33100 21412
rect 34244 21360 34296 21412
rect 34612 21360 34664 21412
rect 36084 21437 36093 21471
rect 36093 21437 36127 21471
rect 36127 21437 36136 21471
rect 36084 21428 36136 21437
rect 55220 21471 55272 21480
rect 55220 21437 55229 21471
rect 55229 21437 55263 21471
rect 55263 21437 55272 21471
rect 55680 21471 55732 21480
rect 55220 21428 55272 21437
rect 55680 21437 55689 21471
rect 55689 21437 55723 21471
rect 55723 21437 55732 21471
rect 55680 21428 55732 21437
rect 56876 21471 56928 21480
rect 56876 21437 56885 21471
rect 56885 21437 56919 21471
rect 56919 21437 56928 21471
rect 56876 21428 56928 21437
rect 57520 21471 57572 21480
rect 57520 21437 57529 21471
rect 57529 21437 57563 21471
rect 57563 21437 57572 21471
rect 57520 21428 57572 21437
rect 57704 21471 57756 21480
rect 57704 21437 57713 21471
rect 57713 21437 57747 21471
rect 57747 21437 57756 21471
rect 57704 21428 57756 21437
rect 48044 21360 48096 21412
rect 33968 21292 34020 21344
rect 34060 21292 34112 21344
rect 34520 21292 34572 21344
rect 55220 21292 55272 21344
rect 57428 21292 57480 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 50326 21190 50378 21242
rect 50390 21190 50442 21242
rect 50454 21190 50506 21242
rect 50518 21190 50570 21242
rect 3516 21088 3568 21140
rect 4712 21088 4764 21140
rect 4804 21088 4856 21140
rect 2780 21020 2832 21072
rect 2596 20952 2648 21004
rect 2688 20952 2740 21004
rect 5632 21020 5684 21072
rect 7196 21063 7248 21072
rect 7196 21029 7205 21063
rect 7205 21029 7239 21063
rect 7239 21029 7248 21063
rect 7196 21020 7248 21029
rect 11152 21020 11204 21072
rect 12808 21020 12860 21072
rect 5448 20952 5500 21004
rect 6368 20995 6420 21004
rect 6368 20961 6377 20995
rect 6377 20961 6411 20995
rect 6411 20961 6420 20995
rect 6368 20952 6420 20961
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 8392 20995 8444 21004
rect 8392 20961 8401 20995
rect 8401 20961 8435 20995
rect 8435 20961 8444 20995
rect 8392 20952 8444 20961
rect 8484 20952 8536 21004
rect 11612 20995 11664 21004
rect 11612 20961 11621 20995
rect 11621 20961 11655 20995
rect 11655 20961 11664 20995
rect 11612 20952 11664 20961
rect 15108 21088 15160 21140
rect 15200 21088 15252 21140
rect 17592 21088 17644 21140
rect 17868 21131 17920 21140
rect 17868 21097 17877 21131
rect 17877 21097 17911 21131
rect 17911 21097 17920 21131
rect 17868 21088 17920 21097
rect 20076 21088 20128 21140
rect 20260 21131 20312 21140
rect 20260 21097 20269 21131
rect 20269 21097 20303 21131
rect 20303 21097 20312 21131
rect 20260 21088 20312 21097
rect 20812 21088 20864 21140
rect 23112 21088 23164 21140
rect 17684 21020 17736 21072
rect 14832 20952 14884 21004
rect 15476 20952 15528 21004
rect 3792 20884 3844 20936
rect 7380 20927 7432 20936
rect 7380 20893 7389 20927
rect 7389 20893 7423 20927
rect 7423 20893 7432 20927
rect 7380 20884 7432 20893
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 14556 20884 14608 20936
rect 4620 20816 4672 20868
rect 1952 20791 2004 20800
rect 1952 20757 1961 20791
rect 1961 20757 1995 20791
rect 1995 20757 2004 20791
rect 1952 20748 2004 20757
rect 2688 20791 2740 20800
rect 2688 20757 2697 20791
rect 2697 20757 2731 20791
rect 2731 20757 2740 20791
rect 2688 20748 2740 20757
rect 5632 20748 5684 20800
rect 10784 20748 10836 20800
rect 10968 20748 11020 20800
rect 12624 20748 12676 20800
rect 17040 20995 17092 21004
rect 17040 20961 17049 20995
rect 17049 20961 17083 20995
rect 17083 20961 17092 20995
rect 17040 20952 17092 20961
rect 17960 20995 18012 21004
rect 17960 20961 17969 20995
rect 17969 20961 18003 20995
rect 18003 20961 18012 20995
rect 17960 20952 18012 20961
rect 19248 20952 19300 21004
rect 21548 21020 21600 21072
rect 23664 21020 23716 21072
rect 23848 21088 23900 21140
rect 25412 21131 25464 21140
rect 25412 21097 25421 21131
rect 25421 21097 25455 21131
rect 25455 21097 25464 21131
rect 25412 21088 25464 21097
rect 31024 21088 31076 21140
rect 31484 21088 31536 21140
rect 32956 21088 33008 21140
rect 34152 21088 34204 21140
rect 28908 21020 28960 21072
rect 19156 20884 19208 20936
rect 19708 20884 19760 20936
rect 20352 20884 20404 20936
rect 20444 20884 20496 20936
rect 24952 20952 25004 21004
rect 25320 20995 25372 21004
rect 25320 20961 25329 20995
rect 25329 20961 25363 20995
rect 25363 20961 25372 20995
rect 25320 20952 25372 20961
rect 25872 20952 25924 21004
rect 26516 20995 26568 21004
rect 26516 20961 26525 20995
rect 26525 20961 26559 20995
rect 26559 20961 26568 20995
rect 26516 20952 26568 20961
rect 26608 20995 26660 21004
rect 26608 20961 26617 20995
rect 26617 20961 26651 20995
rect 26651 20961 26660 20995
rect 26608 20952 26660 20961
rect 27620 20952 27672 21004
rect 26884 20927 26936 20936
rect 26884 20893 26893 20927
rect 26893 20893 26927 20927
rect 26927 20893 26936 20927
rect 28724 20952 28776 21004
rect 30380 21020 30432 21072
rect 33324 21020 33376 21072
rect 29276 20952 29328 21004
rect 31208 20995 31260 21004
rect 31208 20961 31217 20995
rect 31217 20961 31251 20995
rect 31251 20961 31260 20995
rect 31208 20952 31260 20961
rect 31392 20952 31444 21004
rect 31576 20995 31628 21004
rect 31576 20961 31585 20995
rect 31585 20961 31619 20995
rect 31619 20961 31628 20995
rect 31576 20952 31628 20961
rect 32588 20995 32640 21004
rect 32588 20961 32597 20995
rect 32597 20961 32631 20995
rect 32631 20961 32640 20995
rect 32588 20952 32640 20961
rect 33968 21020 34020 21072
rect 35716 21020 35768 21072
rect 26884 20884 26936 20893
rect 19800 20816 19852 20868
rect 20076 20859 20128 20868
rect 20076 20825 20085 20859
rect 20085 20825 20119 20859
rect 20119 20825 20128 20859
rect 20076 20816 20128 20825
rect 20720 20816 20772 20868
rect 30932 20884 30984 20936
rect 34336 20995 34388 21004
rect 34336 20961 34345 20995
rect 34345 20961 34379 20995
rect 34379 20961 34388 20995
rect 34336 20952 34388 20961
rect 36084 20995 36136 21004
rect 36084 20961 36093 20995
rect 36093 20961 36127 20995
rect 36127 20961 36136 20995
rect 36084 20952 36136 20961
rect 57704 21088 57756 21140
rect 57520 21020 57572 21072
rect 33692 20927 33744 20936
rect 33692 20893 33701 20927
rect 33701 20893 33735 20927
rect 33735 20893 33744 20927
rect 33692 20884 33744 20893
rect 28540 20816 28592 20868
rect 29000 20816 29052 20868
rect 32496 20816 32548 20868
rect 33968 20884 34020 20936
rect 55220 20952 55272 21004
rect 56048 20952 56100 21004
rect 58164 20995 58216 21004
rect 58164 20961 58173 20995
rect 58173 20961 58207 20995
rect 58207 20961 58216 20995
rect 58164 20952 58216 20961
rect 36452 20884 36504 20936
rect 15476 20748 15528 20800
rect 15936 20748 15988 20800
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 16212 20748 16264 20800
rect 17408 20748 17460 20800
rect 19708 20748 19760 20800
rect 26700 20748 26752 20800
rect 29736 20748 29788 20800
rect 31944 20748 31996 20800
rect 36084 20748 36136 20800
rect 55680 20816 55732 20868
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 2044 20544 2096 20596
rect 7196 20544 7248 20596
rect 10324 20544 10376 20596
rect 11796 20544 11848 20596
rect 12256 20587 12308 20596
rect 12256 20553 12265 20587
rect 12265 20553 12299 20587
rect 12299 20553 12308 20587
rect 12256 20544 12308 20553
rect 13268 20587 13320 20596
rect 13268 20553 13277 20587
rect 13277 20553 13311 20587
rect 13311 20553 13320 20587
rect 13268 20544 13320 20553
rect 14096 20544 14148 20596
rect 14832 20587 14884 20596
rect 14832 20553 14841 20587
rect 14841 20553 14875 20587
rect 14875 20553 14884 20587
rect 14832 20544 14884 20553
rect 6000 20476 6052 20528
rect 2688 20340 2740 20392
rect 5080 20383 5132 20392
rect 3056 20315 3108 20324
rect 3056 20281 3065 20315
rect 3065 20281 3099 20315
rect 3099 20281 3108 20315
rect 3608 20315 3660 20324
rect 3056 20272 3108 20281
rect 3608 20281 3617 20315
rect 3617 20281 3651 20315
rect 3651 20281 3660 20315
rect 3608 20272 3660 20281
rect 5080 20349 5089 20383
rect 5089 20349 5123 20383
rect 5123 20349 5132 20383
rect 5080 20340 5132 20349
rect 5356 20272 5408 20324
rect 5632 20272 5684 20324
rect 5448 20204 5500 20256
rect 5540 20204 5592 20256
rect 7012 20315 7064 20324
rect 7012 20281 7021 20315
rect 7021 20281 7055 20315
rect 7055 20281 7064 20315
rect 7564 20315 7616 20324
rect 7012 20272 7064 20281
rect 7564 20281 7573 20315
rect 7573 20281 7607 20315
rect 7607 20281 7616 20315
rect 7564 20272 7616 20281
rect 8484 20340 8536 20392
rect 8852 20383 8904 20392
rect 8024 20272 8076 20324
rect 8852 20349 8861 20383
rect 8861 20349 8895 20383
rect 8895 20349 8904 20383
rect 8852 20340 8904 20349
rect 13912 20476 13964 20528
rect 22928 20544 22980 20596
rect 23020 20587 23072 20596
rect 23020 20553 23029 20587
rect 23029 20553 23063 20587
rect 23063 20553 23072 20587
rect 23020 20544 23072 20553
rect 10600 20408 10652 20460
rect 13544 20408 13596 20460
rect 14280 20408 14332 20460
rect 9128 20340 9180 20392
rect 10140 20383 10192 20392
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 10692 20383 10744 20392
rect 10692 20349 10701 20383
rect 10701 20349 10735 20383
rect 10735 20349 10744 20383
rect 10692 20340 10744 20349
rect 12072 20383 12124 20392
rect 12072 20349 12081 20383
rect 12081 20349 12115 20383
rect 12115 20349 12124 20383
rect 12072 20340 12124 20349
rect 13820 20340 13872 20392
rect 15292 20408 15344 20460
rect 16028 20408 16080 20460
rect 15016 20383 15068 20392
rect 12348 20272 12400 20324
rect 15016 20349 15025 20383
rect 15025 20349 15059 20383
rect 15059 20349 15068 20383
rect 15016 20340 15068 20349
rect 16120 20340 16172 20392
rect 17500 20340 17552 20392
rect 17684 20383 17736 20392
rect 17684 20349 17693 20383
rect 17693 20349 17727 20383
rect 17727 20349 17736 20383
rect 17684 20340 17736 20349
rect 18880 20408 18932 20460
rect 19524 20476 19576 20528
rect 20996 20476 21048 20528
rect 21272 20476 21324 20528
rect 23480 20544 23532 20596
rect 23940 20544 23992 20596
rect 25412 20587 25464 20596
rect 25412 20553 25436 20587
rect 25436 20553 25464 20587
rect 25412 20544 25464 20553
rect 25872 20587 25924 20596
rect 25872 20553 25881 20587
rect 25881 20553 25915 20587
rect 25915 20553 25924 20587
rect 25872 20544 25924 20553
rect 26516 20544 26568 20596
rect 29000 20544 29052 20596
rect 30656 20544 30708 20596
rect 33324 20544 33376 20596
rect 34612 20544 34664 20596
rect 56048 20544 56100 20596
rect 56876 20587 56928 20596
rect 56876 20553 56885 20587
rect 56885 20553 56919 20587
rect 56919 20553 56928 20587
rect 56876 20544 56928 20553
rect 19984 20408 20036 20460
rect 18512 20340 18564 20392
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 19616 20340 19668 20392
rect 20536 20408 20588 20460
rect 20628 20408 20680 20460
rect 20168 20340 20220 20392
rect 20904 20383 20956 20392
rect 20904 20349 20913 20383
rect 20913 20349 20947 20383
rect 20947 20349 20956 20383
rect 20904 20340 20956 20349
rect 21548 20408 21600 20460
rect 24032 20476 24084 20528
rect 27712 20476 27764 20528
rect 30932 20476 30984 20528
rect 25596 20451 25648 20460
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 10876 20247 10928 20256
rect 10876 20213 10885 20247
rect 10885 20213 10919 20247
rect 10919 20213 10928 20247
rect 10876 20204 10928 20213
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 15568 20204 15620 20256
rect 15844 20204 15896 20256
rect 21180 20272 21232 20324
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23572 20383 23624 20392
rect 23296 20340 23348 20349
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 25596 20417 25605 20451
rect 25605 20417 25639 20451
rect 25639 20417 25648 20451
rect 25596 20408 25648 20417
rect 27804 20451 27856 20460
rect 27804 20417 27813 20451
rect 27813 20417 27847 20451
rect 27847 20417 27856 20451
rect 27804 20408 27856 20417
rect 23572 20340 23624 20349
rect 23664 20272 23716 20324
rect 25504 20340 25556 20392
rect 26424 20315 26476 20324
rect 20076 20204 20128 20256
rect 20628 20204 20680 20256
rect 20904 20204 20956 20256
rect 21272 20204 21324 20256
rect 22192 20204 22244 20256
rect 24584 20204 24636 20256
rect 26424 20281 26433 20315
rect 26433 20281 26467 20315
rect 26467 20281 26476 20315
rect 26424 20272 26476 20281
rect 29276 20272 29328 20324
rect 29736 20340 29788 20392
rect 31576 20408 31628 20460
rect 31484 20340 31536 20392
rect 31944 20451 31996 20460
rect 31944 20417 31953 20451
rect 31953 20417 31987 20451
rect 31987 20417 31996 20451
rect 31944 20408 31996 20417
rect 32864 20408 32916 20460
rect 34520 20408 34572 20460
rect 36452 20451 36504 20460
rect 33048 20383 33100 20392
rect 30932 20272 30984 20324
rect 33048 20349 33057 20383
rect 33057 20349 33091 20383
rect 33091 20349 33100 20383
rect 33048 20340 33100 20349
rect 33140 20340 33192 20392
rect 36452 20417 36461 20451
rect 36461 20417 36495 20451
rect 36495 20417 36504 20451
rect 36452 20408 36504 20417
rect 36084 20383 36136 20392
rect 32588 20272 32640 20324
rect 36084 20349 36093 20383
rect 36093 20349 36127 20383
rect 36127 20349 36136 20383
rect 36084 20340 36136 20349
rect 36268 20383 36320 20392
rect 36268 20349 36277 20383
rect 36277 20349 36311 20383
rect 36311 20349 36320 20383
rect 36268 20340 36320 20349
rect 26884 20204 26936 20256
rect 29368 20204 29420 20256
rect 29644 20204 29696 20256
rect 35992 20272 36044 20324
rect 55220 20383 55272 20392
rect 55220 20349 55229 20383
rect 55229 20349 55263 20383
rect 55263 20349 55272 20383
rect 55220 20340 55272 20349
rect 55404 20340 55456 20392
rect 56048 20340 56100 20392
rect 56968 20340 57020 20392
rect 57704 20383 57756 20392
rect 57704 20349 57713 20383
rect 57713 20349 57747 20383
rect 57747 20349 57756 20383
rect 57704 20340 57756 20349
rect 56508 20272 56560 20324
rect 56784 20315 56836 20324
rect 56784 20281 56793 20315
rect 56793 20281 56827 20315
rect 56827 20281 56836 20315
rect 56784 20272 56836 20281
rect 55220 20204 55272 20256
rect 55772 20204 55824 20256
rect 56140 20204 56192 20256
rect 57980 20204 58032 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 50326 20102 50378 20154
rect 50390 20102 50442 20154
rect 50454 20102 50506 20154
rect 50518 20102 50570 20154
rect 2964 20000 3016 20052
rect 2504 19975 2556 19984
rect 2504 19941 2513 19975
rect 2513 19941 2547 19975
rect 2547 19941 2556 19975
rect 2504 19932 2556 19941
rect 7932 20000 7984 20052
rect 4620 19932 4672 19984
rect 10876 19932 10928 19984
rect 5724 19864 5776 19916
rect 8484 19907 8536 19916
rect 8484 19873 8493 19907
rect 8493 19873 8527 19907
rect 8527 19873 8536 19907
rect 8484 19864 8536 19873
rect 8576 19864 8628 19916
rect 11336 19864 11388 19916
rect 12256 20000 12308 20052
rect 12348 20000 12400 20052
rect 50988 20000 51040 20052
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 14188 19932 14240 19984
rect 21456 19932 21508 19984
rect 12072 19864 12124 19916
rect 12256 19864 12308 19916
rect 13360 19907 13412 19916
rect 4804 19839 4856 19848
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 2964 19771 3016 19780
rect 2964 19737 2973 19771
rect 2973 19737 3007 19771
rect 3007 19737 3016 19771
rect 2964 19728 3016 19737
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 7288 19796 7340 19848
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 6368 19728 6420 19780
rect 12440 19796 12492 19848
rect 12900 19796 12952 19848
rect 13360 19873 13369 19907
rect 13369 19873 13403 19907
rect 13403 19873 13412 19907
rect 13360 19864 13412 19873
rect 14924 19864 14976 19916
rect 15016 19907 15068 19916
rect 15016 19873 15025 19907
rect 15025 19873 15059 19907
rect 15059 19873 15068 19907
rect 15752 19907 15804 19916
rect 15016 19864 15068 19873
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 15752 19864 15804 19873
rect 13176 19839 13228 19848
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 16212 19864 16264 19916
rect 18880 19907 18932 19916
rect 13176 19796 13228 19805
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 20812 19864 20864 19916
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 22192 19932 22244 19984
rect 14188 19728 14240 19780
rect 15476 19728 15528 19780
rect 20628 19796 20680 19848
rect 5816 19703 5868 19712
rect 5816 19669 5825 19703
rect 5825 19669 5859 19703
rect 5859 19669 5868 19703
rect 5816 19660 5868 19669
rect 10692 19660 10744 19712
rect 12440 19660 12492 19712
rect 13544 19703 13596 19712
rect 13544 19669 13553 19703
rect 13553 19669 13587 19703
rect 13587 19669 13596 19703
rect 13544 19660 13596 19669
rect 14832 19703 14884 19712
rect 14832 19669 14841 19703
rect 14841 19669 14875 19703
rect 14875 19669 14884 19703
rect 14832 19660 14884 19669
rect 15016 19660 15068 19712
rect 19984 19728 20036 19780
rect 18236 19660 18288 19712
rect 18972 19703 19024 19712
rect 18972 19669 18981 19703
rect 18981 19669 19015 19703
rect 19015 19669 19024 19703
rect 18972 19660 19024 19669
rect 19064 19660 19116 19712
rect 19892 19660 19944 19712
rect 20720 19728 20772 19780
rect 21272 19728 21324 19780
rect 21456 19728 21508 19780
rect 21732 19864 21784 19916
rect 21916 19907 21968 19916
rect 21916 19873 21925 19907
rect 21925 19873 21959 19907
rect 21959 19873 21968 19907
rect 21916 19864 21968 19873
rect 24124 19932 24176 19984
rect 24492 19932 24544 19984
rect 26608 19975 26660 19984
rect 26608 19941 26617 19975
rect 26617 19941 26651 19975
rect 26651 19941 26660 19975
rect 26608 19932 26660 19941
rect 27712 19975 27764 19984
rect 27712 19941 27721 19975
rect 27721 19941 27755 19975
rect 27755 19941 27764 19975
rect 27712 19932 27764 19941
rect 28356 19975 28408 19984
rect 28356 19941 28365 19975
rect 28365 19941 28399 19975
rect 28399 19941 28408 19975
rect 28356 19932 28408 19941
rect 28724 19932 28776 19984
rect 36268 19932 36320 19984
rect 23020 19907 23072 19916
rect 23020 19873 23029 19907
rect 23029 19873 23063 19907
rect 23063 19873 23072 19907
rect 23020 19864 23072 19873
rect 23204 19864 23256 19916
rect 23572 19864 23624 19916
rect 24032 19907 24084 19916
rect 24032 19873 24041 19907
rect 24041 19873 24075 19907
rect 24075 19873 24084 19907
rect 24032 19864 24084 19873
rect 24216 19864 24268 19916
rect 24584 19864 24636 19916
rect 25320 19907 25372 19916
rect 25320 19873 25330 19907
rect 25330 19873 25364 19907
rect 25364 19873 25372 19907
rect 25504 19907 25556 19916
rect 25320 19864 25372 19873
rect 25504 19873 25513 19907
rect 25513 19873 25547 19907
rect 25547 19873 25556 19907
rect 25504 19864 25556 19873
rect 25136 19796 25188 19848
rect 26700 19864 26752 19916
rect 26976 19864 27028 19916
rect 27620 19907 27672 19916
rect 25780 19796 25832 19848
rect 27068 19839 27120 19848
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 27620 19873 27629 19907
rect 27629 19873 27663 19907
rect 27663 19873 27672 19907
rect 27620 19864 27672 19873
rect 28264 19907 28316 19916
rect 28264 19873 28273 19907
rect 28273 19873 28307 19907
rect 28307 19873 28316 19907
rect 28264 19864 28316 19873
rect 28632 19864 28684 19916
rect 28816 19864 28868 19916
rect 31024 19864 31076 19916
rect 32588 19864 32640 19916
rect 32864 19907 32916 19916
rect 32864 19873 32873 19907
rect 32873 19873 32907 19907
rect 32907 19873 32916 19907
rect 32864 19864 32916 19873
rect 33968 19864 34020 19916
rect 53748 19907 53800 19916
rect 53748 19873 53757 19907
rect 53757 19873 53791 19907
rect 53791 19873 53800 19907
rect 56784 19932 56836 19984
rect 57980 19975 58032 19984
rect 57980 19941 57989 19975
rect 57989 19941 58023 19975
rect 58023 19941 58032 19975
rect 57980 19932 58032 19941
rect 58164 19907 58216 19916
rect 53748 19864 53800 19873
rect 58164 19873 58173 19907
rect 58173 19873 58207 19907
rect 58207 19873 58216 19907
rect 58164 19864 58216 19873
rect 27896 19796 27948 19848
rect 30932 19839 30984 19848
rect 30932 19805 30941 19839
rect 30941 19805 30975 19839
rect 30975 19805 30984 19839
rect 30932 19796 30984 19805
rect 25688 19728 25740 19780
rect 54300 19839 54352 19848
rect 54300 19805 54309 19839
rect 54309 19805 54343 19839
rect 54343 19805 54352 19839
rect 54300 19796 54352 19805
rect 56692 19839 56744 19848
rect 56692 19805 56701 19839
rect 56701 19805 56735 19839
rect 56735 19805 56744 19839
rect 56692 19796 56744 19805
rect 56876 19839 56928 19848
rect 56876 19805 56885 19839
rect 56885 19805 56919 19839
rect 56919 19805 56928 19839
rect 56876 19796 56928 19805
rect 22652 19703 22704 19712
rect 22652 19669 22661 19703
rect 22661 19669 22695 19703
rect 22695 19669 22704 19703
rect 22652 19660 22704 19669
rect 23480 19660 23532 19712
rect 24676 19660 24728 19712
rect 26148 19660 26200 19712
rect 57980 19660 58032 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 2504 19456 2556 19508
rect 5080 19456 5132 19508
rect 7012 19456 7064 19508
rect 5448 19388 5500 19440
rect 14004 19456 14056 19508
rect 14188 19499 14240 19508
rect 14188 19465 14197 19499
rect 14197 19465 14231 19499
rect 14231 19465 14240 19499
rect 14188 19456 14240 19465
rect 14924 19456 14976 19508
rect 15752 19456 15804 19508
rect 19064 19499 19116 19508
rect 19064 19465 19073 19499
rect 19073 19465 19107 19499
rect 19107 19465 19116 19499
rect 19064 19456 19116 19465
rect 20076 19456 20128 19508
rect 20720 19456 20772 19508
rect 20812 19456 20864 19508
rect 21732 19456 21784 19508
rect 23296 19456 23348 19508
rect 24676 19499 24728 19508
rect 14096 19431 14148 19440
rect 14096 19397 14105 19431
rect 14105 19397 14139 19431
rect 14139 19397 14148 19431
rect 14096 19388 14148 19397
rect 15384 19388 15436 19440
rect 9680 19320 9732 19372
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 20444 19388 20496 19440
rect 24676 19465 24685 19499
rect 24685 19465 24719 19499
rect 24719 19465 24728 19499
rect 24676 19456 24728 19465
rect 25504 19456 25556 19508
rect 27068 19456 27120 19508
rect 28724 19499 28776 19508
rect 28724 19465 28733 19499
rect 28733 19465 28767 19499
rect 28767 19465 28776 19499
rect 28724 19456 28776 19465
rect 29920 19499 29972 19508
rect 29920 19465 29929 19499
rect 29929 19465 29963 19499
rect 29963 19465 29972 19499
rect 29920 19456 29972 19465
rect 30932 19456 30984 19508
rect 33048 19456 33100 19508
rect 56968 19456 57020 19508
rect 57704 19456 57756 19508
rect 27620 19388 27672 19440
rect 2596 19295 2648 19304
rect 2596 19261 2605 19295
rect 2605 19261 2639 19295
rect 2639 19261 2648 19295
rect 2596 19252 2648 19261
rect 3792 19295 3844 19304
rect 3792 19261 3801 19295
rect 3801 19261 3835 19295
rect 3835 19261 3844 19295
rect 3792 19252 3844 19261
rect 4712 19295 4764 19304
rect 3148 19184 3200 19236
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 5356 19295 5408 19304
rect 5356 19261 5365 19295
rect 5365 19261 5399 19295
rect 5399 19261 5408 19295
rect 5356 19252 5408 19261
rect 10784 19295 10836 19304
rect 5264 19184 5316 19236
rect 4528 19116 4580 19168
rect 5632 19116 5684 19168
rect 8024 19227 8076 19236
rect 8024 19193 8033 19227
rect 8033 19193 8067 19227
rect 8067 19193 8076 19227
rect 8944 19227 8996 19236
rect 8024 19184 8076 19193
rect 8944 19193 8953 19227
rect 8953 19193 8987 19227
rect 8987 19193 8996 19227
rect 8944 19184 8996 19193
rect 10784 19261 10793 19295
rect 10793 19261 10827 19295
rect 10827 19261 10836 19295
rect 10784 19252 10836 19261
rect 11152 19252 11204 19304
rect 11612 19252 11664 19304
rect 12164 19295 12216 19304
rect 12164 19261 12173 19295
rect 12173 19261 12207 19295
rect 12207 19261 12216 19295
rect 12164 19252 12216 19261
rect 12440 19295 12492 19304
rect 12440 19261 12474 19295
rect 12474 19261 12492 19295
rect 12440 19252 12492 19261
rect 15016 19252 15068 19304
rect 12072 19184 12124 19236
rect 10048 19116 10100 19168
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10508 19116 10560 19168
rect 12992 19184 13044 19236
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 16396 19252 16448 19304
rect 16488 19252 16540 19304
rect 17684 19320 17736 19372
rect 17868 19295 17920 19304
rect 16672 19184 16724 19236
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18880 19252 18932 19304
rect 19340 19295 19392 19304
rect 19340 19261 19379 19295
rect 19379 19261 19392 19295
rect 19340 19252 19392 19261
rect 19524 19184 19576 19236
rect 16488 19116 16540 19168
rect 17684 19116 17736 19168
rect 18972 19116 19024 19168
rect 19156 19116 19208 19168
rect 19892 19252 19944 19304
rect 24216 19320 24268 19372
rect 20904 19252 20956 19304
rect 21456 19252 21508 19304
rect 21916 19252 21968 19304
rect 22836 19252 22888 19304
rect 23480 19295 23532 19304
rect 23480 19261 23489 19295
rect 23489 19261 23523 19295
rect 23523 19261 23532 19295
rect 23480 19252 23532 19261
rect 23848 19252 23900 19304
rect 23756 19227 23808 19236
rect 23756 19193 23765 19227
rect 23765 19193 23799 19227
rect 23799 19193 23808 19227
rect 23756 19184 23808 19193
rect 21180 19116 21232 19168
rect 26976 19320 27028 19372
rect 27160 19320 27212 19372
rect 26608 19295 26660 19304
rect 24676 19184 24728 19236
rect 26608 19261 26617 19295
rect 26617 19261 26651 19295
rect 26651 19261 26660 19295
rect 26608 19252 26660 19261
rect 26700 19252 26752 19304
rect 26976 19184 27028 19236
rect 28908 19252 28960 19304
rect 29092 19252 29144 19304
rect 29552 19252 29604 19304
rect 29828 19252 29880 19304
rect 31208 19252 31260 19304
rect 31484 19295 31536 19304
rect 31484 19261 31493 19295
rect 31493 19261 31527 19295
rect 31527 19261 31536 19295
rect 31484 19252 31536 19261
rect 56140 19295 56192 19304
rect 56140 19261 56149 19295
rect 56149 19261 56183 19295
rect 56183 19261 56192 19295
rect 56140 19252 56192 19261
rect 57428 19295 57480 19304
rect 57428 19261 57437 19295
rect 57437 19261 57471 19295
rect 57471 19261 57480 19295
rect 57428 19252 57480 19261
rect 57980 19295 58032 19304
rect 57980 19261 57989 19295
rect 57989 19261 58023 19295
rect 58023 19261 58032 19295
rect 57980 19252 58032 19261
rect 58164 19295 58216 19304
rect 58164 19261 58173 19295
rect 58173 19261 58207 19295
rect 58207 19261 58216 19295
rect 58164 19252 58216 19261
rect 30564 19184 30616 19236
rect 26516 19116 26568 19168
rect 27896 19159 27948 19168
rect 27896 19125 27905 19159
rect 27905 19125 27939 19159
rect 27939 19125 27948 19159
rect 27896 19116 27948 19125
rect 28632 19116 28684 19168
rect 31116 19116 31168 19168
rect 31576 19159 31628 19168
rect 31576 19125 31585 19159
rect 31585 19125 31619 19159
rect 31619 19125 31628 19159
rect 31576 19116 31628 19125
rect 56876 19116 56928 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 50326 19014 50378 19066
rect 50390 19014 50442 19066
rect 50454 19014 50506 19066
rect 50518 19014 50570 19066
rect 3056 18912 3108 18964
rect 4712 18912 4764 18964
rect 6368 18955 6420 18964
rect 2044 18887 2096 18896
rect 2044 18853 2053 18887
rect 2053 18853 2087 18887
rect 2087 18853 2096 18887
rect 2044 18844 2096 18853
rect 6368 18921 6377 18955
rect 6377 18921 6411 18955
rect 6411 18921 6420 18955
rect 6368 18912 6420 18921
rect 6920 18912 6972 18964
rect 8024 18912 8076 18964
rect 10048 18912 10100 18964
rect 5908 18844 5960 18896
rect 2136 18776 2188 18828
rect 3148 18776 3200 18828
rect 6092 18776 6144 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 7012 18776 7064 18828
rect 8852 18844 8904 18896
rect 12440 18912 12492 18964
rect 12532 18955 12584 18964
rect 12532 18921 12541 18955
rect 12541 18921 12575 18955
rect 12575 18921 12584 18955
rect 12532 18912 12584 18921
rect 13360 18912 13412 18964
rect 13452 18912 13504 18964
rect 8116 18776 8168 18828
rect 9680 18776 9732 18828
rect 3424 18708 3476 18760
rect 13544 18844 13596 18896
rect 14832 18844 14884 18896
rect 15200 18844 15252 18896
rect 15476 18844 15528 18896
rect 12992 18819 13044 18828
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 12992 18785 13001 18819
rect 13001 18785 13035 18819
rect 13035 18785 13044 18819
rect 12992 18776 13044 18785
rect 13636 18819 13688 18828
rect 12532 18640 12584 18692
rect 12900 18640 12952 18692
rect 13360 18640 13412 18692
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 15292 18776 15344 18828
rect 8484 18572 8536 18624
rect 12992 18615 13044 18624
rect 12992 18581 13001 18615
rect 13001 18581 13035 18615
rect 13035 18581 13044 18615
rect 12992 18572 13044 18581
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 14924 18572 14976 18624
rect 16672 18955 16724 18964
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 19340 18912 19392 18964
rect 20076 18955 20128 18964
rect 16396 18844 16448 18896
rect 19248 18844 19300 18896
rect 17776 18776 17828 18828
rect 18972 18776 19024 18828
rect 20076 18921 20085 18955
rect 20085 18921 20119 18955
rect 20119 18921 20128 18955
rect 20076 18912 20128 18921
rect 20996 18912 21048 18964
rect 28908 18955 28960 18964
rect 28908 18921 28917 18955
rect 28917 18921 28951 18955
rect 28951 18921 28960 18955
rect 28908 18912 28960 18921
rect 29184 18912 29236 18964
rect 31024 18955 31076 18964
rect 31024 18921 31033 18955
rect 31033 18921 31067 18955
rect 31067 18921 31076 18955
rect 31024 18912 31076 18921
rect 16856 18708 16908 18760
rect 21180 18776 21232 18828
rect 21916 18776 21968 18828
rect 22652 18844 22704 18896
rect 23756 18844 23808 18896
rect 56692 18844 56744 18896
rect 23480 18776 23532 18828
rect 23848 18776 23900 18828
rect 24124 18776 24176 18828
rect 20996 18751 21048 18760
rect 20996 18717 21005 18751
rect 21005 18717 21039 18751
rect 21039 18717 21048 18751
rect 20996 18708 21048 18717
rect 21640 18708 21692 18760
rect 22008 18751 22060 18760
rect 20076 18640 20128 18692
rect 21548 18640 21600 18692
rect 20260 18572 20312 18624
rect 22008 18717 22017 18751
rect 22017 18717 22051 18751
rect 22051 18717 22060 18751
rect 22008 18708 22060 18717
rect 25964 18819 26016 18828
rect 25964 18785 25994 18819
rect 25994 18785 26016 18819
rect 26148 18819 26200 18828
rect 25964 18776 26016 18785
rect 26148 18785 26157 18819
rect 26157 18785 26191 18819
rect 26191 18785 26200 18819
rect 26148 18776 26200 18785
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 26976 18776 27028 18828
rect 28356 18776 28408 18828
rect 29368 18819 29420 18828
rect 29368 18785 29377 18819
rect 29377 18785 29411 18819
rect 29411 18785 29420 18819
rect 29368 18776 29420 18785
rect 30472 18776 30524 18828
rect 30932 18819 30984 18828
rect 30932 18785 30941 18819
rect 30941 18785 30975 18819
rect 30975 18785 30984 18819
rect 30932 18776 30984 18785
rect 31116 18819 31168 18828
rect 31116 18785 31125 18819
rect 31125 18785 31159 18819
rect 31159 18785 31168 18819
rect 31116 18776 31168 18785
rect 55588 18819 55640 18828
rect 55588 18785 55597 18819
rect 55597 18785 55631 18819
rect 55631 18785 55640 18819
rect 55588 18776 55640 18785
rect 57980 18819 58032 18828
rect 57980 18785 57989 18819
rect 57989 18785 58023 18819
rect 58023 18785 58032 18819
rect 57980 18776 58032 18785
rect 26516 18708 26568 18760
rect 26148 18640 26200 18692
rect 28724 18708 28776 18760
rect 31944 18708 31996 18760
rect 58164 18683 58216 18692
rect 58164 18649 58173 18683
rect 58173 18649 58207 18683
rect 58207 18649 58216 18683
rect 58164 18640 58216 18649
rect 21824 18572 21876 18624
rect 23020 18572 23072 18624
rect 24216 18572 24268 18624
rect 25504 18615 25556 18624
rect 25504 18581 25513 18615
rect 25513 18581 25547 18615
rect 25547 18581 25556 18615
rect 25504 18572 25556 18581
rect 26424 18572 26476 18624
rect 57520 18572 57572 18624
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 5724 18411 5776 18420
rect 5724 18377 5733 18411
rect 5733 18377 5767 18411
rect 5767 18377 5776 18411
rect 5724 18368 5776 18377
rect 6092 18368 6144 18420
rect 12440 18368 12492 18420
rect 12532 18368 12584 18420
rect 16764 18368 16816 18420
rect 18972 18411 19024 18420
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 12256 18300 12308 18352
rect 12624 18300 12676 18352
rect 13636 18300 13688 18352
rect 6184 18232 6236 18284
rect 7840 18232 7892 18284
rect 9680 18232 9732 18284
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 10692 18164 10744 18216
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 12900 18164 12952 18216
rect 13820 18232 13872 18284
rect 8484 18139 8536 18148
rect 8484 18105 8493 18139
rect 8493 18105 8527 18139
rect 8527 18105 8536 18139
rect 12440 18139 12492 18148
rect 8484 18096 8536 18105
rect 12440 18105 12449 18139
rect 12449 18105 12483 18139
rect 12483 18105 12492 18139
rect 12440 18096 12492 18105
rect 10140 18028 10192 18080
rect 10324 18071 10376 18080
rect 10324 18037 10333 18071
rect 10333 18037 10367 18071
rect 10367 18037 10376 18071
rect 10324 18028 10376 18037
rect 11244 18028 11296 18080
rect 13912 18096 13964 18148
rect 15568 18300 15620 18352
rect 18420 18300 18472 18352
rect 21364 18368 21416 18420
rect 23664 18368 23716 18420
rect 21456 18343 21508 18352
rect 21456 18309 21465 18343
rect 21465 18309 21499 18343
rect 21499 18309 21508 18343
rect 21456 18300 21508 18309
rect 22008 18300 22060 18352
rect 26332 18368 26384 18420
rect 28356 18368 28408 18420
rect 29276 18411 29328 18420
rect 29276 18377 29285 18411
rect 29285 18377 29319 18411
rect 29319 18377 29328 18411
rect 29276 18368 29328 18377
rect 57980 18411 58032 18420
rect 57980 18377 57989 18411
rect 57989 18377 58023 18411
rect 58023 18377 58032 18411
rect 57980 18368 58032 18377
rect 14924 18232 14976 18284
rect 14648 18096 14700 18148
rect 16028 18164 16080 18216
rect 17776 18232 17828 18284
rect 19984 18232 20036 18284
rect 20260 18232 20312 18284
rect 17316 18207 17368 18216
rect 17316 18173 17325 18207
rect 17325 18173 17359 18207
rect 17359 18173 17368 18207
rect 17316 18164 17368 18173
rect 17960 18164 18012 18216
rect 18236 18164 18288 18216
rect 19156 18207 19208 18216
rect 17868 18096 17920 18148
rect 19156 18173 19165 18207
rect 19165 18173 19199 18207
rect 19199 18173 19208 18207
rect 19156 18164 19208 18173
rect 21364 18232 21416 18284
rect 14188 18028 14240 18080
rect 16120 18028 16172 18080
rect 20168 18028 20220 18080
rect 21824 18232 21876 18284
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 22836 18207 22888 18216
rect 20996 18096 21048 18148
rect 22836 18173 22845 18207
rect 22845 18173 22879 18207
rect 22879 18173 22888 18207
rect 22836 18164 22888 18173
rect 26148 18232 26200 18284
rect 28540 18232 28592 18284
rect 57520 18275 57572 18284
rect 26056 18207 26108 18216
rect 21640 18096 21692 18148
rect 26056 18173 26065 18207
rect 26065 18173 26099 18207
rect 26099 18173 26108 18207
rect 26056 18164 26108 18173
rect 26792 18164 26844 18216
rect 26884 18164 26936 18216
rect 28632 18207 28684 18216
rect 24768 18096 24820 18148
rect 25780 18096 25832 18148
rect 28632 18173 28641 18207
rect 28641 18173 28675 18207
rect 28675 18173 28684 18207
rect 28632 18164 28684 18173
rect 57520 18241 57529 18275
rect 57529 18241 57563 18275
rect 57563 18241 57572 18275
rect 57520 18232 57572 18241
rect 56232 18207 56284 18216
rect 56232 18173 56241 18207
rect 56241 18173 56275 18207
rect 56275 18173 56284 18207
rect 56232 18164 56284 18173
rect 57060 18207 57112 18216
rect 57060 18173 57069 18207
rect 57069 18173 57103 18207
rect 57103 18173 57112 18207
rect 57060 18164 57112 18173
rect 57428 18164 57480 18216
rect 30932 18096 30984 18148
rect 21916 18028 21968 18080
rect 24032 18028 24084 18080
rect 24676 18028 24728 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 50326 17926 50378 17978
rect 50390 17926 50442 17978
rect 50454 17926 50506 17978
rect 50518 17926 50570 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 14004 17824 14056 17876
rect 15200 17824 15252 17876
rect 20076 17824 20128 17876
rect 21364 17867 21416 17876
rect 2320 17756 2372 17808
rect 10600 17799 10652 17808
rect 10600 17765 10609 17799
rect 10609 17765 10643 17799
rect 10643 17765 10652 17799
rect 10600 17756 10652 17765
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 14004 17688 14056 17740
rect 15660 17756 15712 17808
rect 20168 17756 20220 17808
rect 21364 17833 21373 17867
rect 21373 17833 21407 17867
rect 21407 17833 21416 17867
rect 21364 17824 21416 17833
rect 21916 17867 21968 17876
rect 21916 17833 21925 17867
rect 21925 17833 21959 17867
rect 21959 17833 21968 17867
rect 21916 17824 21968 17833
rect 23480 17824 23532 17876
rect 25320 17867 25372 17876
rect 25320 17833 25329 17867
rect 25329 17833 25363 17867
rect 25363 17833 25372 17867
rect 25320 17824 25372 17833
rect 26608 17824 26660 17876
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 16304 17688 16356 17740
rect 19984 17731 20036 17740
rect 19984 17697 19993 17731
rect 19993 17697 20027 17731
rect 20027 17697 20036 17731
rect 19984 17688 20036 17697
rect 21824 17731 21876 17740
rect 21824 17697 21833 17731
rect 21833 17697 21867 17731
rect 21867 17697 21876 17731
rect 21824 17688 21876 17697
rect 22836 17731 22888 17740
rect 22836 17697 22845 17731
rect 22845 17697 22879 17731
rect 22879 17697 22888 17731
rect 22836 17688 22888 17697
rect 23388 17756 23440 17808
rect 24032 17731 24084 17740
rect 24032 17697 24041 17731
rect 24041 17697 24075 17731
rect 24075 17697 24084 17731
rect 24032 17688 24084 17697
rect 25136 17688 25188 17740
rect 25504 17756 25556 17808
rect 58164 17799 58216 17808
rect 58164 17765 58173 17799
rect 58173 17765 58207 17799
rect 58207 17765 58216 17799
rect 58164 17756 58216 17765
rect 10508 17663 10560 17672
rect 10508 17629 10517 17663
rect 10517 17629 10551 17663
rect 10551 17629 10560 17663
rect 10508 17620 10560 17629
rect 1768 17552 1820 17604
rect 25780 17620 25832 17672
rect 12164 17552 12216 17604
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 13820 17484 13872 17536
rect 55404 17620 55456 17672
rect 26148 17484 26200 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 14004 17280 14056 17332
rect 21640 17280 21692 17332
rect 24768 17323 24820 17332
rect 24768 17289 24777 17323
rect 24777 17289 24811 17323
rect 24811 17289 24820 17323
rect 24768 17280 24820 17289
rect 25780 17280 25832 17332
rect 55220 17280 55272 17332
rect 55404 17323 55456 17332
rect 55404 17289 55413 17323
rect 55413 17289 55447 17323
rect 55447 17289 55456 17323
rect 55404 17280 55456 17289
rect 56324 17255 56376 17264
rect 56324 17221 56333 17255
rect 56333 17221 56367 17255
rect 56367 17221 56376 17255
rect 56324 17212 56376 17221
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10416 17144 10468 17196
rect 12992 17144 13044 17196
rect 14188 17144 14240 17196
rect 20352 17144 20404 17196
rect 23388 17187 23440 17196
rect 5540 17076 5592 17128
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 9772 17076 9824 17085
rect 2044 17051 2096 17060
rect 2044 17017 2053 17051
rect 2053 17017 2087 17051
rect 2087 17017 2096 17051
rect 2044 17008 2096 17017
rect 12256 17051 12308 17060
rect 12256 17017 12265 17051
rect 12265 17017 12299 17051
rect 12299 17017 12308 17051
rect 13176 17051 13228 17060
rect 12256 17008 12308 17017
rect 13176 17017 13185 17051
rect 13185 17017 13219 17051
rect 13219 17017 13228 17051
rect 13176 17008 13228 17017
rect 13820 17051 13872 17060
rect 13820 17017 13829 17051
rect 13829 17017 13863 17051
rect 13863 17017 13872 17051
rect 13820 17008 13872 17017
rect 9680 16940 9732 16992
rect 14740 17008 14792 17060
rect 21364 17076 21416 17128
rect 22836 17119 22888 17128
rect 22836 17085 22845 17119
rect 22845 17085 22879 17119
rect 22879 17085 22888 17119
rect 22836 17076 22888 17085
rect 23388 17153 23397 17187
rect 23397 17153 23431 17187
rect 23431 17153 23440 17187
rect 23388 17144 23440 17153
rect 24124 17119 24176 17128
rect 24124 17085 24133 17119
rect 24133 17085 24167 17119
rect 24167 17085 24176 17119
rect 24124 17076 24176 17085
rect 55772 17076 55824 17128
rect 57060 17119 57112 17128
rect 57060 17085 57069 17119
rect 57069 17085 57103 17119
rect 57103 17085 57112 17119
rect 57060 17076 57112 17085
rect 57520 17119 57572 17128
rect 57520 17085 57529 17119
rect 57529 17085 57563 17119
rect 57563 17085 57572 17119
rect 57520 17076 57572 17085
rect 53748 17008 53800 17060
rect 57980 16940 58032 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 50326 16838 50378 16890
rect 50390 16838 50442 16890
rect 50454 16838 50506 16890
rect 50518 16838 50570 16890
rect 1860 16736 1912 16788
rect 9680 16736 9732 16788
rect 10600 16779 10652 16788
rect 10600 16745 10609 16779
rect 10609 16745 10643 16779
rect 10643 16745 10652 16779
rect 10600 16736 10652 16745
rect 13912 16736 13964 16788
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 2136 16668 2188 16720
rect 10416 16668 10468 16720
rect 21548 16668 21600 16720
rect 9772 16600 9824 16652
rect 12072 16600 12124 16652
rect 22836 16643 22888 16652
rect 22836 16609 22845 16643
rect 22845 16609 22879 16643
rect 22879 16609 22888 16643
rect 22836 16600 22888 16609
rect 24216 16643 24268 16652
rect 24216 16609 24225 16643
rect 24225 16609 24259 16643
rect 24259 16609 24268 16643
rect 24216 16600 24268 16609
rect 26056 16600 26108 16652
rect 55772 16643 55824 16652
rect 55772 16609 55781 16643
rect 55781 16609 55815 16643
rect 55815 16609 55824 16643
rect 55772 16600 55824 16609
rect 57980 16711 58032 16720
rect 57980 16677 57989 16711
rect 57989 16677 58023 16711
rect 58023 16677 58032 16711
rect 57980 16668 58032 16677
rect 58164 16711 58216 16720
rect 58164 16677 58173 16711
rect 58173 16677 58207 16711
rect 58207 16677 58216 16711
rect 58164 16668 58216 16677
rect 57980 16532 58032 16584
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 56600 16192 56652 16244
rect 57520 16124 57572 16176
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 4712 16056 4764 16108
rect 4988 16056 5040 16108
rect 5816 15988 5868 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 55588 15988 55640 16040
rect 56324 15988 56376 16040
rect 15016 15963 15068 15972
rect 15016 15929 15025 15963
rect 15025 15929 15059 15963
rect 15059 15929 15068 15963
rect 15016 15920 15068 15929
rect 57060 15920 57112 15972
rect 58164 15920 58216 15972
rect 56324 15895 56376 15904
rect 56324 15861 56333 15895
rect 56333 15861 56367 15895
rect 56367 15861 56376 15895
rect 56324 15852 56376 15861
rect 58072 15895 58124 15904
rect 58072 15861 58081 15895
rect 58081 15861 58115 15895
rect 58115 15861 58124 15895
rect 58072 15852 58124 15861
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 50326 15750 50378 15802
rect 50390 15750 50442 15802
rect 50454 15750 50506 15802
rect 50518 15750 50570 15802
rect 58164 15691 58216 15700
rect 58164 15657 58173 15691
rect 58173 15657 58207 15691
rect 58207 15657 58216 15691
rect 58164 15648 58216 15657
rect 56324 15512 56376 15564
rect 56692 15512 56744 15564
rect 56876 15555 56928 15564
rect 56876 15521 56885 15555
rect 56885 15521 56919 15555
rect 56919 15521 56928 15555
rect 56876 15512 56928 15521
rect 56968 15351 57020 15360
rect 56968 15317 56977 15351
rect 56977 15317 57011 15351
rect 57011 15317 57020 15351
rect 56968 15308 57020 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 1952 15147 2004 15156
rect 1952 15113 1961 15147
rect 1961 15113 1995 15147
rect 1995 15113 2004 15147
rect 1952 15104 2004 15113
rect 55220 15104 55272 15156
rect 56876 15104 56928 15156
rect 58256 15036 58308 15088
rect 7380 14900 7432 14952
rect 55772 14900 55824 14952
rect 56140 14943 56192 14952
rect 56140 14909 56149 14943
rect 56149 14909 56183 14943
rect 56183 14909 56192 14943
rect 56140 14900 56192 14909
rect 57980 14943 58032 14952
rect 57980 14909 57989 14943
rect 57989 14909 58023 14943
rect 58023 14909 58032 14943
rect 57980 14900 58032 14909
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 50326 14662 50378 14714
rect 50390 14662 50442 14714
rect 50454 14662 50506 14714
rect 50518 14662 50570 14714
rect 7564 14492 7616 14544
rect 55588 14467 55640 14476
rect 55588 14433 55597 14467
rect 55597 14433 55631 14467
rect 55631 14433 55640 14467
rect 55588 14424 55640 14433
rect 56600 14424 56652 14476
rect 55772 14356 55824 14408
rect 53840 14288 53892 14340
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 55772 14059 55824 14068
rect 55772 14025 55781 14059
rect 55781 14025 55815 14059
rect 55815 14025 55824 14059
rect 55772 14016 55824 14025
rect 56784 13948 56836 14000
rect 56140 13812 56192 13864
rect 56692 13812 56744 13864
rect 57152 13812 57204 13864
rect 57520 13855 57572 13864
rect 57520 13821 57529 13855
rect 57529 13821 57563 13855
rect 57563 13821 57572 13855
rect 57520 13812 57572 13821
rect 58164 13719 58216 13728
rect 58164 13685 58173 13719
rect 58173 13685 58207 13719
rect 58207 13685 58216 13719
rect 58164 13676 58216 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 50326 13574 50378 13626
rect 50390 13574 50442 13626
rect 50454 13574 50506 13626
rect 50518 13574 50570 13626
rect 58072 13515 58124 13524
rect 58072 13481 58081 13515
rect 58081 13481 58115 13515
rect 58115 13481 58124 13515
rect 58072 13472 58124 13481
rect 7472 13404 7524 13456
rect 57520 13404 57572 13456
rect 58164 13404 58216 13456
rect 56784 13336 56836 13388
rect 2044 13243 2096 13252
rect 2044 13209 2053 13243
rect 2053 13209 2087 13243
rect 2087 13209 2096 13243
rect 2044 13200 2096 13209
rect 23388 13200 23440 13252
rect 57244 13175 57296 13184
rect 57244 13141 57253 13175
rect 57253 13141 57287 13175
rect 57287 13141 57296 13175
rect 57244 13132 57296 13141
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 56140 12928 56192 12980
rect 57336 12971 57388 12980
rect 57336 12937 57345 12971
rect 57345 12937 57379 12971
rect 57379 12937 57388 12971
rect 57336 12928 57388 12937
rect 55404 12767 55456 12776
rect 55404 12733 55413 12767
rect 55413 12733 55447 12767
rect 55447 12733 55456 12767
rect 55404 12724 55456 12733
rect 56048 12767 56100 12776
rect 56048 12733 56057 12767
rect 56057 12733 56091 12767
rect 56091 12733 56100 12767
rect 56048 12724 56100 12733
rect 57244 12767 57296 12776
rect 57244 12733 57253 12767
rect 57253 12733 57287 12767
rect 57287 12733 57296 12767
rect 57244 12724 57296 12733
rect 57980 12699 58032 12708
rect 57980 12665 57989 12699
rect 57989 12665 58023 12699
rect 58023 12665 58032 12699
rect 57980 12656 58032 12665
rect 57888 12588 57940 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 50326 12486 50378 12538
rect 50390 12486 50442 12538
rect 50454 12486 50506 12538
rect 50518 12486 50570 12538
rect 1952 12427 2004 12436
rect 1952 12393 1961 12427
rect 1961 12393 1995 12427
rect 1995 12393 2004 12427
rect 1952 12384 2004 12393
rect 57980 12384 58032 12436
rect 4896 12316 4948 12368
rect 56876 12291 56928 12300
rect 56876 12257 56885 12291
rect 56885 12257 56919 12291
rect 56919 12257 56928 12291
rect 56876 12248 56928 12257
rect 55588 12180 55640 12232
rect 57704 12223 57756 12232
rect 57704 12189 57713 12223
rect 57713 12189 57747 12223
rect 57747 12189 57756 12223
rect 57704 12180 57756 12189
rect 56508 12044 56560 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 55588 11883 55640 11892
rect 55588 11849 55597 11883
rect 55597 11849 55631 11883
rect 55631 11849 55640 11883
rect 55588 11840 55640 11849
rect 56876 11840 56928 11892
rect 4804 11636 4856 11688
rect 56140 11636 56192 11688
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 50326 11398 50378 11450
rect 50390 11398 50442 11450
rect 50454 11398 50506 11450
rect 50518 11398 50570 11450
rect 57704 11296 57756 11348
rect 55588 11203 55640 11212
rect 55588 11169 55597 11203
rect 55597 11169 55631 11203
rect 55631 11169 55640 11203
rect 55588 11160 55640 11169
rect 57152 11160 57204 11212
rect 57980 11203 58032 11212
rect 57980 11169 57989 11203
rect 57989 11169 58023 11203
rect 58023 11169 58032 11203
rect 57980 11160 58032 11169
rect 57888 11024 57940 11076
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 57980 10795 58032 10804
rect 57980 10761 57989 10795
rect 57989 10761 58023 10795
rect 58023 10761 58032 10795
rect 57980 10752 58032 10761
rect 3608 10548 3660 10600
rect 57152 10548 57204 10600
rect 57244 10548 57296 10600
rect 2044 10523 2096 10532
rect 2044 10489 2053 10523
rect 2053 10489 2087 10523
rect 2087 10489 2096 10523
rect 2044 10480 2096 10489
rect 57704 10412 57756 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 50326 10310 50378 10362
rect 50390 10310 50442 10362
rect 50454 10310 50506 10362
rect 50518 10310 50570 10362
rect 57244 10251 57296 10260
rect 57244 10217 57253 10251
rect 57253 10217 57287 10251
rect 57287 10217 57296 10251
rect 57244 10208 57296 10217
rect 55588 10115 55640 10124
rect 55588 10081 55597 10115
rect 55597 10081 55631 10115
rect 55631 10081 55640 10115
rect 55588 10072 55640 10081
rect 57152 10072 57204 10124
rect 57612 10072 57664 10124
rect 58164 9979 58216 9988
rect 58164 9945 58173 9979
rect 58173 9945 58207 9979
rect 58207 9945 58216 9979
rect 58164 9936 58216 9945
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 57612 9639 57664 9648
rect 57612 9605 57621 9639
rect 57621 9605 57655 9639
rect 57655 9605 57664 9639
rect 57612 9596 57664 9605
rect 4068 9460 4120 9512
rect 55680 9503 55732 9512
rect 55680 9469 55689 9503
rect 55689 9469 55723 9503
rect 55723 9469 55732 9503
rect 55680 9460 55732 9469
rect 56784 9460 56836 9512
rect 56968 9503 57020 9512
rect 56968 9469 56977 9503
rect 56977 9469 57011 9503
rect 57011 9469 57020 9503
rect 56968 9460 57020 9469
rect 57152 9503 57204 9512
rect 57152 9469 57161 9503
rect 57161 9469 57195 9503
rect 57195 9469 57204 9503
rect 57152 9460 57204 9469
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 50326 9222 50378 9274
rect 50390 9222 50442 9274
rect 50454 9222 50506 9274
rect 50518 9222 50570 9274
rect 57152 9120 57204 9172
rect 2964 9052 3016 9104
rect 56140 9052 56192 9104
rect 56968 8984 57020 9036
rect 57704 9027 57756 9036
rect 57704 8993 57713 9027
rect 57713 8993 57747 9027
rect 57747 8993 57756 9027
rect 57704 8984 57756 8993
rect 1952 8823 2004 8832
rect 1952 8789 1961 8823
rect 1961 8789 1995 8823
rect 1995 8789 2004 8823
rect 1952 8780 2004 8789
rect 57980 8823 58032 8832
rect 57980 8789 57989 8823
rect 57989 8789 58023 8823
rect 58023 8789 58032 8823
rect 57980 8780 58032 8789
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 56140 8619 56192 8628
rect 56140 8585 56149 8619
rect 56149 8585 56183 8619
rect 56183 8585 56192 8619
rect 56140 8576 56192 8585
rect 57336 8508 57388 8560
rect 58164 8551 58216 8560
rect 58164 8517 58173 8551
rect 58173 8517 58207 8551
rect 58207 8517 58216 8551
rect 58164 8508 58216 8517
rect 56416 8440 56468 8492
rect 57428 8483 57480 8492
rect 57428 8449 57437 8483
rect 57437 8449 57471 8483
rect 57471 8449 57480 8483
rect 57428 8440 57480 8449
rect 56048 8372 56100 8424
rect 57980 8415 58032 8424
rect 57980 8381 57989 8415
rect 57989 8381 58023 8415
rect 58023 8381 58032 8415
rect 57980 8372 58032 8381
rect 55772 8304 55824 8356
rect 56140 8304 56192 8356
rect 57520 8304 57572 8356
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 50326 8134 50378 8186
rect 50390 8134 50442 8186
rect 50454 8134 50506 8186
rect 50518 8134 50570 8186
rect 1860 8007 1912 8016
rect 1860 7973 1869 8007
rect 1869 7973 1903 8007
rect 1903 7973 1912 8007
rect 1860 7964 1912 7973
rect 55128 7896 55180 7948
rect 56784 7896 56836 7948
rect 57336 7939 57388 7948
rect 57336 7905 57345 7939
rect 57345 7905 57379 7939
rect 57379 7905 57388 7939
rect 57336 7896 57388 7905
rect 2044 7803 2096 7812
rect 2044 7769 2053 7803
rect 2053 7769 2087 7803
rect 2087 7769 2096 7803
rect 2044 7760 2096 7769
rect 57336 7760 57388 7812
rect 57520 7803 57572 7812
rect 57520 7769 57529 7803
rect 57529 7769 57563 7803
rect 57563 7769 57572 7803
rect 57520 7760 57572 7769
rect 55680 7692 55732 7744
rect 56232 7692 56284 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 52552 7488 52604 7540
rect 55220 7352 55272 7404
rect 55404 7284 55456 7336
rect 55588 7284 55640 7336
rect 56416 7327 56468 7336
rect 56048 7216 56100 7268
rect 56416 7293 56425 7327
rect 56425 7293 56459 7327
rect 56459 7293 56468 7327
rect 56416 7284 56468 7293
rect 57704 7327 57756 7336
rect 57704 7293 57713 7327
rect 57713 7293 57747 7327
rect 57747 7293 57756 7327
rect 57704 7284 57756 7293
rect 57244 7216 57296 7268
rect 55680 7148 55732 7200
rect 56508 7148 56560 7200
rect 57980 7148 58032 7200
rect 58072 7148 58124 7200
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 50326 7046 50378 7098
rect 50390 7046 50442 7098
rect 50454 7046 50506 7098
rect 50518 7046 50570 7098
rect 53748 6876 53800 6928
rect 57060 6944 57112 6996
rect 14648 6808 14700 6860
rect 52552 6851 52604 6860
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 52552 6817 52561 6851
rect 52561 6817 52595 6851
rect 52595 6817 52604 6851
rect 52552 6808 52604 6817
rect 55772 6851 55824 6860
rect 55772 6817 55781 6851
rect 55781 6817 55815 6851
rect 55815 6817 55824 6851
rect 55772 6808 55824 6817
rect 57980 6851 58032 6860
rect 57980 6817 57989 6851
rect 57989 6817 58023 6851
rect 58023 6817 58032 6851
rect 57980 6808 58032 6817
rect 58164 6851 58216 6860
rect 58164 6817 58173 6851
rect 58173 6817 58207 6851
rect 58207 6817 58216 6851
rect 58164 6808 58216 6817
rect 55496 6672 55548 6724
rect 54300 6604 54352 6656
rect 54484 6647 54536 6656
rect 54484 6613 54493 6647
rect 54493 6613 54527 6647
rect 54527 6613 54536 6647
rect 54484 6604 54536 6613
rect 55864 6604 55916 6656
rect 56140 6604 56192 6656
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 57704 6400 57756 6452
rect 52460 6332 52512 6384
rect 52368 6196 52420 6248
rect 55496 6264 55548 6316
rect 56416 6332 56468 6384
rect 56600 6332 56652 6384
rect 57428 6332 57480 6384
rect 54024 6196 54076 6248
rect 54944 6239 54996 6248
rect 54944 6205 54953 6239
rect 54953 6205 54987 6239
rect 54987 6205 54996 6239
rect 54944 6196 54996 6205
rect 55588 6239 55640 6248
rect 55588 6205 55597 6239
rect 55597 6205 55631 6239
rect 55631 6205 55640 6239
rect 55588 6196 55640 6205
rect 56140 6239 56192 6248
rect 56140 6205 56149 6239
rect 56149 6205 56183 6239
rect 56183 6205 56192 6239
rect 56140 6196 56192 6205
rect 56508 6264 56560 6316
rect 56968 6239 57020 6248
rect 56692 6128 56744 6180
rect 56968 6205 56977 6239
rect 56977 6205 57011 6239
rect 57011 6205 57020 6239
rect 56968 6196 57020 6205
rect 57152 6128 57204 6180
rect 54760 6103 54812 6112
rect 54760 6069 54769 6103
rect 54769 6069 54803 6103
rect 54803 6069 54812 6103
rect 54760 6060 54812 6069
rect 55864 6060 55916 6112
rect 57244 6060 57296 6112
rect 57888 6060 57940 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 50326 5958 50378 6010
rect 50390 5958 50442 6010
rect 50454 5958 50506 6010
rect 50518 5958 50570 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 56968 5856 57020 5908
rect 1860 5831 1912 5840
rect 1860 5797 1869 5831
rect 1869 5797 1903 5831
rect 1903 5797 1912 5831
rect 1860 5788 1912 5797
rect 29552 5720 29604 5772
rect 52460 5763 52512 5772
rect 52460 5729 52469 5763
rect 52469 5729 52503 5763
rect 52503 5729 52512 5763
rect 52460 5720 52512 5729
rect 53748 5763 53800 5772
rect 53748 5729 53757 5763
rect 53757 5729 53791 5763
rect 53791 5729 53800 5763
rect 53748 5720 53800 5729
rect 55680 5788 55732 5840
rect 57612 5788 57664 5840
rect 58164 5831 58216 5840
rect 58164 5797 58173 5831
rect 58173 5797 58207 5831
rect 58207 5797 58216 5831
rect 58164 5788 58216 5797
rect 56508 5720 56560 5772
rect 56692 5763 56744 5772
rect 56692 5729 56701 5763
rect 56701 5729 56735 5763
rect 56735 5729 56744 5763
rect 56692 5720 56744 5729
rect 58072 5720 58124 5772
rect 56784 5652 56836 5704
rect 14740 5516 14792 5568
rect 15016 5516 15068 5568
rect 29552 5516 29604 5568
rect 53104 5559 53156 5568
rect 53104 5525 53113 5559
rect 53113 5525 53147 5559
rect 53147 5525 53156 5559
rect 53104 5516 53156 5525
rect 56876 5516 56928 5568
rect 57060 5559 57112 5568
rect 57060 5525 57069 5559
rect 57069 5525 57103 5559
rect 57103 5525 57112 5559
rect 57060 5516 57112 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 53196 5312 53248 5364
rect 54944 5312 54996 5364
rect 50988 5176 51040 5228
rect 2136 5108 2188 5160
rect 49976 5108 50028 5160
rect 50620 5151 50672 5160
rect 50620 5117 50629 5151
rect 50629 5117 50663 5151
rect 50663 5117 50672 5151
rect 50620 5108 50672 5117
rect 51632 5151 51684 5160
rect 51632 5117 51641 5151
rect 51641 5117 51675 5151
rect 51675 5117 51684 5151
rect 51632 5108 51684 5117
rect 52460 5151 52512 5160
rect 52460 5117 52469 5151
rect 52469 5117 52503 5151
rect 52503 5117 52512 5151
rect 52460 5108 52512 5117
rect 51908 5040 51960 5092
rect 55956 5176 56008 5228
rect 57336 5176 57388 5228
rect 57060 5108 57112 5160
rect 57704 5151 57756 5160
rect 57704 5117 57713 5151
rect 57713 5117 57747 5151
rect 57747 5117 57756 5151
rect 57704 5108 57756 5117
rect 55864 5083 55916 5092
rect 55864 5049 55873 5083
rect 55873 5049 55907 5083
rect 55907 5049 55916 5083
rect 55864 5040 55916 5049
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 53288 4972 53340 5024
rect 55772 4972 55824 5024
rect 57060 4972 57112 5024
rect 58164 5015 58216 5024
rect 58164 4981 58173 5015
rect 58173 4981 58207 5015
rect 58207 4981 58216 5015
rect 58164 4972 58216 4981
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 50326 4870 50378 4922
rect 50390 4870 50442 4922
rect 50454 4870 50506 4922
rect 50518 4870 50570 4922
rect 56692 4768 56744 4820
rect 56416 4700 56468 4752
rect 58164 4700 58216 4752
rect 37372 4632 37424 4684
rect 49148 4632 49200 4684
rect 51908 4675 51960 4684
rect 51908 4641 51917 4675
rect 51917 4641 51951 4675
rect 51951 4641 51960 4675
rect 51908 4632 51960 4641
rect 53196 4675 53248 4684
rect 53196 4641 53205 4675
rect 53205 4641 53239 4675
rect 53239 4641 53248 4675
rect 53196 4632 53248 4641
rect 54576 4632 54628 4684
rect 56600 4632 56652 4684
rect 54300 4564 54352 4616
rect 56784 4564 56836 4616
rect 46940 4496 46992 4548
rect 55036 4496 55088 4548
rect 33600 4428 33652 4480
rect 36268 4428 36320 4480
rect 37280 4428 37332 4480
rect 38384 4428 38436 4480
rect 38568 4471 38620 4480
rect 38568 4437 38577 4471
rect 38577 4437 38611 4471
rect 38611 4437 38620 4471
rect 38568 4428 38620 4437
rect 39396 4428 39448 4480
rect 39488 4428 39540 4480
rect 41512 4471 41564 4480
rect 41512 4437 41521 4471
rect 41521 4437 41555 4471
rect 41555 4437 41564 4471
rect 41512 4428 41564 4437
rect 42340 4471 42392 4480
rect 42340 4437 42349 4471
rect 42349 4437 42383 4471
rect 42383 4437 42392 4471
rect 42340 4428 42392 4437
rect 43444 4471 43496 4480
rect 43444 4437 43453 4471
rect 43453 4437 43487 4471
rect 43487 4437 43496 4471
rect 43444 4428 43496 4437
rect 47032 4471 47084 4480
rect 47032 4437 47041 4471
rect 47041 4437 47075 4471
rect 47075 4437 47084 4471
rect 47032 4428 47084 4437
rect 48044 4471 48096 4480
rect 48044 4437 48053 4471
rect 48053 4437 48087 4471
rect 48087 4437 48096 4471
rect 48044 4428 48096 4437
rect 48964 4428 49016 4480
rect 49056 4428 49108 4480
rect 49700 4428 49752 4480
rect 51724 4471 51776 4480
rect 51724 4437 51733 4471
rect 51733 4437 51767 4471
rect 51767 4437 51776 4471
rect 51724 4428 51776 4437
rect 53748 4428 53800 4480
rect 54392 4428 54444 4480
rect 55312 4428 55364 4480
rect 55588 4471 55640 4480
rect 55588 4437 55597 4471
rect 55597 4437 55631 4471
rect 55631 4437 55640 4471
rect 55588 4428 55640 4437
rect 56968 4471 57020 4480
rect 56968 4437 56977 4471
rect 56977 4437 57011 4471
rect 57011 4437 57020 4471
rect 56968 4428 57020 4437
rect 57980 4471 58032 4480
rect 57980 4437 57989 4471
rect 57989 4437 58023 4471
rect 58023 4437 58032 4471
rect 57980 4428 58032 4437
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 34796 4199 34848 4208
rect 34796 4165 34805 4199
rect 34805 4165 34839 4199
rect 34839 4165 34848 4199
rect 34796 4156 34848 4165
rect 44272 4156 44324 4208
rect 45744 4199 45796 4208
rect 45744 4165 45753 4199
rect 45753 4165 45787 4199
rect 45787 4165 45796 4199
rect 45744 4156 45796 4165
rect 54392 4156 54444 4208
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 2044 4088 2096 4097
rect 30012 4020 30064 4072
rect 33048 4020 33100 4072
rect 13176 3952 13228 4004
rect 35256 4020 35308 4072
rect 36084 4063 36136 4072
rect 36084 4029 36093 4063
rect 36093 4029 36127 4063
rect 36127 4029 36136 4063
rect 36084 4020 36136 4029
rect 37372 4063 37424 4072
rect 37372 4029 37381 4063
rect 37381 4029 37415 4063
rect 37415 4029 37424 4063
rect 37372 4020 37424 4029
rect 41236 4063 41288 4072
rect 41236 4029 41245 4063
rect 41245 4029 41279 4063
rect 41279 4029 41288 4063
rect 41236 4020 41288 4029
rect 42432 4020 42484 4072
rect 43904 4020 43956 4072
rect 47676 4063 47728 4072
rect 47676 4029 47685 4063
rect 47685 4029 47719 4063
rect 47719 4029 47728 4063
rect 47676 4020 47728 4029
rect 49148 4063 49200 4072
rect 49148 4029 49157 4063
rect 49157 4029 49191 4063
rect 49191 4029 49200 4063
rect 49148 4020 49200 4029
rect 47216 3952 47268 4004
rect 33784 3884 33836 3936
rect 34520 3884 34572 3936
rect 34888 3884 34940 3936
rect 37556 3884 37608 3936
rect 39580 3884 39632 3936
rect 39764 3927 39816 3936
rect 39764 3893 39773 3927
rect 39773 3893 39807 3927
rect 39807 3893 39816 3927
rect 39764 3884 39816 3893
rect 40408 3927 40460 3936
rect 40408 3893 40417 3927
rect 40417 3893 40451 3927
rect 40451 3893 40460 3927
rect 40408 3884 40460 3893
rect 41880 3927 41932 3936
rect 41880 3893 41889 3927
rect 41889 3893 41923 3927
rect 41923 3893 41932 3927
rect 41880 3884 41932 3893
rect 43720 3884 43772 3936
rect 44456 3884 44508 3936
rect 47124 3884 47176 3936
rect 49792 4020 49844 4072
rect 55036 4088 55088 4140
rect 56508 4088 56560 4140
rect 58532 4088 58584 4140
rect 50988 4020 51040 4072
rect 51908 4020 51960 4072
rect 53196 4020 53248 4072
rect 54576 4020 54628 4072
rect 55680 4020 55732 4072
rect 56232 4063 56284 4072
rect 56232 4029 56241 4063
rect 56241 4029 56275 4063
rect 56275 4029 56284 4063
rect 56232 4020 56284 4029
rect 57980 4063 58032 4072
rect 57980 4029 57989 4063
rect 57989 4029 58023 4063
rect 58023 4029 58032 4063
rect 57980 4020 58032 4029
rect 54116 3995 54168 4004
rect 49884 3884 49936 3936
rect 51540 3884 51592 3936
rect 52000 3884 52052 3936
rect 52828 3884 52880 3936
rect 54116 3961 54125 3995
rect 54125 3961 54159 3995
rect 54159 3961 54168 3995
rect 54116 3952 54168 3961
rect 54668 3952 54720 4004
rect 58164 3995 58216 4004
rect 58164 3961 58173 3995
rect 58173 3961 58207 3995
rect 58207 3961 58216 3995
rect 58164 3952 58216 3961
rect 53932 3884 53984 3936
rect 54852 3884 54904 3936
rect 56600 3884 56652 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 50326 3782 50378 3834
rect 50390 3782 50442 3834
rect 50454 3782 50506 3834
rect 50518 3782 50570 3834
rect 7840 3612 7892 3664
rect 11244 3655 11296 3664
rect 11244 3621 11253 3655
rect 11253 3621 11287 3655
rect 11287 3621 11296 3655
rect 11244 3612 11296 3621
rect 37372 3680 37424 3732
rect 43904 3723 43956 3732
rect 43904 3689 43913 3723
rect 43913 3689 43947 3723
rect 43947 3689 43956 3723
rect 43904 3680 43956 3689
rect 54116 3680 54168 3732
rect 57704 3680 57756 3732
rect 2320 3544 2372 3596
rect 14740 3544 14792 3596
rect 30656 3587 30708 3596
rect 30656 3553 30665 3587
rect 30665 3553 30699 3587
rect 30699 3553 30708 3587
rect 30656 3544 30708 3553
rect 33416 3544 33468 3596
rect 33968 3544 34020 3596
rect 34336 3544 34388 3596
rect 34888 3544 34940 3596
rect 35440 3544 35492 3596
rect 36084 3544 36136 3596
rect 11060 3476 11112 3528
rect 37740 3544 37792 3596
rect 38660 3544 38712 3596
rect 39304 3587 39356 3596
rect 39304 3553 39313 3587
rect 39313 3553 39347 3587
rect 39347 3553 39356 3587
rect 39304 3544 39356 3553
rect 41052 3587 41104 3596
rect 41052 3553 41061 3587
rect 41061 3553 41095 3587
rect 41095 3553 41104 3587
rect 41052 3544 41104 3553
rect 42432 3587 42484 3596
rect 42432 3553 42441 3587
rect 42441 3553 42475 3587
rect 42475 3553 42484 3587
rect 42432 3544 42484 3553
rect 43076 3544 43128 3596
rect 55588 3655 55640 3664
rect 55588 3621 55597 3655
rect 55597 3621 55631 3655
rect 55631 3621 55640 3655
rect 55588 3612 55640 3621
rect 55680 3612 55732 3664
rect 47216 3544 47268 3596
rect 47584 3587 47636 3596
rect 47584 3553 47593 3587
rect 47593 3553 47627 3587
rect 47627 3553 47636 3587
rect 47584 3544 47636 3553
rect 48504 3587 48556 3596
rect 48504 3553 48513 3587
rect 48513 3553 48547 3587
rect 48547 3553 48556 3587
rect 48504 3544 48556 3553
rect 49884 3544 49936 3596
rect 50160 3544 50212 3596
rect 51448 3544 51500 3596
rect 52644 3544 52696 3596
rect 53104 3587 53156 3596
rect 53104 3553 53113 3587
rect 53113 3553 53147 3587
rect 53147 3553 53156 3587
rect 53104 3544 53156 3553
rect 53288 3587 53340 3596
rect 53288 3553 53297 3587
rect 53297 3553 53331 3587
rect 53331 3553 53340 3587
rect 53288 3544 53340 3553
rect 54300 3587 54352 3596
rect 54300 3553 54309 3587
rect 54309 3553 54343 3587
rect 54343 3553 54352 3587
rect 54300 3544 54352 3553
rect 55312 3544 55364 3596
rect 56784 3544 56836 3596
rect 56968 3544 57020 3596
rect 47676 3476 47728 3528
rect 57428 3476 57480 3528
rect 47216 3408 47268 3460
rect 55956 3408 56008 3460
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 2044 3340 2096 3392
rect 8300 3340 8352 3392
rect 29092 3340 29144 3392
rect 30196 3340 30248 3392
rect 30932 3340 30984 3392
rect 32128 3383 32180 3392
rect 32128 3349 32137 3383
rect 32137 3349 32171 3383
rect 32171 3349 32180 3383
rect 32128 3340 32180 3349
rect 32772 3340 32824 3392
rect 33692 3340 33744 3392
rect 34612 3383 34664 3392
rect 34612 3349 34621 3383
rect 34621 3349 34655 3383
rect 34655 3349 34664 3383
rect 34612 3340 34664 3349
rect 35532 3340 35584 3392
rect 37372 3340 37424 3392
rect 38292 3340 38344 3392
rect 39212 3340 39264 3392
rect 40132 3340 40184 3392
rect 42800 3340 42852 3392
rect 42892 3340 42944 3392
rect 45560 3340 45612 3392
rect 47400 3340 47452 3392
rect 47492 3340 47544 3392
rect 48412 3340 48464 3392
rect 49608 3383 49660 3392
rect 49608 3349 49617 3383
rect 49617 3349 49651 3383
rect 49651 3349 49660 3383
rect 49608 3340 49660 3349
rect 50068 3340 50120 3392
rect 51172 3340 51224 3392
rect 52092 3340 52144 3392
rect 53012 3340 53064 3392
rect 57980 3383 58032 3392
rect 57980 3349 57989 3383
rect 57989 3349 58023 3383
rect 58023 3349 58032 3383
rect 57980 3340 58032 3349
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 1676 3136 1728 3188
rect 2044 3136 2096 3188
rect 3056 3179 3108 3188
rect 3056 3145 3065 3179
rect 3065 3145 3099 3179
rect 3099 3145 3108 3179
rect 3056 3136 3108 3145
rect 33416 3179 33468 3188
rect 33416 3145 33425 3179
rect 33425 3145 33459 3179
rect 33459 3145 33468 3179
rect 33416 3136 33468 3145
rect 35440 3179 35492 3188
rect 35440 3145 35449 3179
rect 35449 3145 35483 3179
rect 35483 3145 35492 3179
rect 35440 3136 35492 3145
rect 38660 3179 38712 3188
rect 38660 3145 38669 3179
rect 38669 3145 38703 3179
rect 38703 3145 38712 3179
rect 38660 3136 38712 3145
rect 39304 3136 39356 3188
rect 47584 3179 47636 3188
rect 47584 3145 47593 3179
rect 47593 3145 47627 3179
rect 47627 3145 47636 3179
rect 47584 3136 47636 3145
rect 51448 3179 51500 3188
rect 51448 3145 51457 3179
rect 51457 3145 51491 3179
rect 51491 3145 51500 3179
rect 51448 3136 51500 3145
rect 54300 3136 54352 3188
rect 54668 3179 54720 3188
rect 54668 3145 54677 3179
rect 54677 3145 54711 3179
rect 54711 3145 54720 3179
rect 54668 3136 54720 3145
rect 55864 3136 55916 3188
rect 56416 3136 56468 3188
rect 4712 3068 4764 3120
rect 30656 3068 30708 3120
rect 49608 3068 49660 3120
rect 480 2932 532 2984
rect 8944 3000 8996 3052
rect 30012 3043 30064 3052
rect 30012 3009 30021 3043
rect 30021 3009 30055 3043
rect 30055 3009 30064 3043
rect 30012 3000 30064 3009
rect 30196 3043 30248 3052
rect 30196 3009 30205 3043
rect 30205 3009 30239 3043
rect 30239 3009 30248 3043
rect 30196 3000 30248 3009
rect 2780 2864 2832 2916
rect 1400 2796 1452 2848
rect 28080 2975 28132 2984
rect 3240 2864 3292 2916
rect 28080 2941 28089 2975
rect 28089 2941 28123 2975
rect 28123 2941 28132 2975
rect 28080 2932 28132 2941
rect 29000 2932 29052 2984
rect 29552 2975 29604 2984
rect 29552 2941 29561 2975
rect 29561 2941 29595 2975
rect 29595 2941 29604 2975
rect 29552 2932 29604 2941
rect 32128 3000 32180 3052
rect 34612 3000 34664 3052
rect 38568 3000 38620 3052
rect 39396 3043 39448 3052
rect 39396 3009 39405 3043
rect 39405 3009 39439 3043
rect 39439 3009 39448 3043
rect 39396 3000 39448 3009
rect 39580 3043 39632 3052
rect 39580 3009 39589 3043
rect 39589 3009 39623 3043
rect 39623 3009 39632 3043
rect 39580 3000 39632 3009
rect 39764 3000 39816 3052
rect 43444 3000 43496 3052
rect 43720 3043 43772 3052
rect 43720 3009 43729 3043
rect 43729 3009 43763 3043
rect 43763 3009 43772 3043
rect 43720 3000 43772 3009
rect 44732 3000 44784 3052
rect 47124 3043 47176 3052
rect 47124 3009 47133 3043
rect 47133 3009 47167 3043
rect 47167 3009 47176 3043
rect 47124 3000 47176 3009
rect 48964 3043 49016 3052
rect 48964 3009 48973 3043
rect 48973 3009 49007 3043
rect 49007 3009 49016 3043
rect 48964 3000 49016 3009
rect 50620 3000 50672 3052
rect 52000 3068 52052 3120
rect 52460 3000 52512 3052
rect 54024 3043 54076 3052
rect 54024 3009 54033 3043
rect 54033 3009 54067 3043
rect 54067 3009 54076 3043
rect 54024 3000 54076 3009
rect 54760 3068 54812 3120
rect 54484 3000 54536 3052
rect 55404 3000 55456 3052
rect 56600 3068 56652 3120
rect 57244 3000 57296 3052
rect 33048 2975 33100 2984
rect 33048 2941 33057 2975
rect 33057 2941 33091 2975
rect 33091 2941 33100 2975
rect 33048 2932 33100 2941
rect 34336 2975 34388 2984
rect 34336 2941 34345 2975
rect 34345 2941 34379 2975
rect 34379 2941 34388 2975
rect 34336 2932 34388 2941
rect 35256 2932 35308 2984
rect 31760 2864 31812 2916
rect 31944 2907 31996 2916
rect 31944 2873 31953 2907
rect 31953 2873 31987 2907
rect 31987 2873 31996 2907
rect 31944 2864 31996 2873
rect 34612 2864 34664 2916
rect 38384 2932 38436 2984
rect 41236 2932 41288 2984
rect 47032 2932 47084 2984
rect 49056 2932 49108 2984
rect 51724 2932 51776 2984
rect 53748 2932 53800 2984
rect 57152 2932 57204 2984
rect 35992 2907 36044 2916
rect 35992 2873 36001 2907
rect 36001 2873 36035 2907
rect 36035 2873 36044 2907
rect 35992 2864 36044 2873
rect 36728 2907 36780 2916
rect 36728 2873 36737 2907
rect 36737 2873 36771 2907
rect 36771 2873 36780 2907
rect 36728 2864 36780 2873
rect 42432 2907 42484 2916
rect 42432 2873 42441 2907
rect 42441 2873 42475 2907
rect 42475 2873 42484 2907
rect 42432 2864 42484 2873
rect 45468 2907 45520 2916
rect 45468 2873 45477 2907
rect 45477 2873 45511 2907
rect 45511 2873 45520 2907
rect 45468 2864 45520 2873
rect 46204 2907 46256 2916
rect 46204 2873 46213 2907
rect 46213 2873 46247 2907
rect 46247 2873 46256 2907
rect 46204 2864 46256 2873
rect 55220 2864 55272 2916
rect 59452 2864 59504 2916
rect 6460 2796 6512 2848
rect 29368 2839 29420 2848
rect 29368 2805 29377 2839
rect 29377 2805 29411 2839
rect 29411 2805 29420 2839
rect 29368 2796 29420 2805
rect 31116 2839 31168 2848
rect 31116 2805 31125 2839
rect 31125 2805 31159 2839
rect 31159 2805 31168 2839
rect 31116 2796 31168 2805
rect 31852 2796 31904 2848
rect 34980 2796 35032 2848
rect 36452 2796 36504 2848
rect 40960 2796 41012 2848
rect 41972 2796 42024 2848
rect 43812 2796 43864 2848
rect 45652 2796 45704 2848
rect 49332 2796 49384 2848
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 50326 2694 50378 2746
rect 50390 2694 50442 2746
rect 50454 2694 50506 2746
rect 50518 2694 50570 2746
rect 31944 2592 31996 2644
rect 35992 2592 36044 2644
rect 36728 2592 36780 2644
rect 41052 2592 41104 2644
rect 42432 2592 42484 2644
rect 45468 2592 45520 2644
rect 46204 2592 46256 2644
rect 48504 2592 48556 2644
rect 50160 2592 50212 2644
rect 56692 2635 56744 2644
rect 56692 2601 56701 2635
rect 56701 2601 56735 2635
rect 56735 2601 56744 2635
rect 56692 2592 56744 2601
rect 11060 2524 11112 2576
rect 31760 2524 31812 2576
rect 53840 2567 53892 2576
rect 53840 2533 53849 2567
rect 53849 2533 53883 2567
rect 53883 2533 53892 2567
rect 53840 2524 53892 2533
rect 55220 2524 55272 2576
rect 56600 2524 56652 2576
rect 57980 2567 58032 2576
rect 57980 2533 57989 2567
rect 57989 2533 58023 2567
rect 58023 2533 58032 2567
rect 57980 2524 58032 2533
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 4160 2456 4212 2508
rect 5080 2499 5132 2508
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 6000 2456 6052 2508
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 7840 2499 7892 2508
rect 6920 2456 6972 2465
rect 7840 2465 7849 2499
rect 7849 2465 7883 2499
rect 7883 2465 7892 2499
rect 7840 2456 7892 2465
rect 8760 2456 8812 2508
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 11520 2456 11572 2508
rect 12440 2456 12492 2508
rect 13360 2456 13412 2508
rect 14280 2456 14332 2508
rect 15200 2456 15252 2508
rect 16120 2456 16172 2508
rect 17040 2456 17092 2508
rect 17960 2456 18012 2508
rect 18880 2499 18932 2508
rect 18880 2465 18889 2499
rect 18889 2465 18923 2499
rect 18923 2465 18932 2499
rect 18880 2456 18932 2465
rect 19800 2456 19852 2508
rect 20720 2456 20772 2508
rect 21640 2499 21692 2508
rect 21640 2465 21649 2499
rect 21649 2465 21683 2499
rect 21683 2465 21692 2499
rect 21640 2456 21692 2465
rect 22560 2456 22612 2508
rect 23480 2456 23532 2508
rect 24400 2499 24452 2508
rect 24400 2465 24409 2499
rect 24409 2465 24443 2499
rect 24443 2465 24452 2499
rect 24400 2456 24452 2465
rect 25320 2456 25372 2508
rect 26240 2499 26292 2508
rect 26240 2465 26249 2499
rect 26249 2465 26283 2499
rect 26283 2465 26292 2499
rect 27160 2499 27212 2508
rect 26240 2456 26292 2465
rect 27160 2465 27169 2499
rect 27169 2465 27203 2499
rect 27203 2465 27212 2499
rect 27160 2456 27212 2465
rect 29092 2499 29144 2508
rect 29092 2465 29101 2499
rect 29101 2465 29135 2499
rect 29135 2465 29144 2499
rect 29092 2456 29144 2465
rect 29368 2456 29420 2508
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 31116 2499 31168 2508
rect 31116 2465 31125 2499
rect 31125 2465 31159 2499
rect 31159 2465 31168 2499
rect 31116 2456 31168 2465
rect 33600 2499 33652 2508
rect 33600 2465 33609 2499
rect 33609 2465 33643 2499
rect 33643 2465 33652 2499
rect 33600 2456 33652 2465
rect 33784 2499 33836 2508
rect 33784 2465 33793 2499
rect 33793 2465 33827 2499
rect 33827 2465 33836 2499
rect 33784 2456 33836 2465
rect 34796 2456 34848 2508
rect 34980 2456 35032 2508
rect 37280 2456 37332 2508
rect 37556 2499 37608 2508
rect 37556 2465 37565 2499
rect 37565 2465 37599 2499
rect 37599 2465 37608 2499
rect 37556 2456 37608 2465
rect 39488 2499 39540 2508
rect 39488 2465 39497 2499
rect 39497 2465 39531 2499
rect 39531 2465 39540 2499
rect 39488 2456 39540 2465
rect 40408 2456 40460 2508
rect 41512 2456 41564 2508
rect 41880 2456 41932 2508
rect 42340 2456 42392 2508
rect 42800 2456 42852 2508
rect 44272 2499 44324 2508
rect 44272 2465 44281 2499
rect 44281 2465 44315 2499
rect 44315 2465 44324 2499
rect 44272 2456 44324 2465
rect 44456 2499 44508 2508
rect 44456 2465 44465 2499
rect 44465 2465 44499 2499
rect 44499 2465 44508 2499
rect 44456 2456 44508 2465
rect 45744 2456 45796 2508
rect 46940 2499 46992 2508
rect 46940 2465 46949 2499
rect 46949 2465 46983 2499
rect 46983 2465 46992 2499
rect 46940 2456 46992 2465
rect 47216 2456 47268 2508
rect 48044 2499 48096 2508
rect 48044 2465 48053 2499
rect 48053 2465 48087 2499
rect 48087 2465 48096 2499
rect 48044 2456 48096 2465
rect 49792 2499 49844 2508
rect 49792 2465 49801 2499
rect 49801 2465 49835 2499
rect 49835 2465 49844 2499
rect 49792 2456 49844 2465
rect 51632 2456 51684 2508
rect 56048 2499 56100 2508
rect 56048 2465 56057 2499
rect 56057 2465 56091 2499
rect 56091 2465 56100 2499
rect 56048 2456 56100 2465
rect 34520 2388 34572 2440
rect 36268 2431 36320 2440
rect 36268 2397 36277 2431
rect 36277 2397 36311 2431
rect 36311 2397 36320 2431
rect 36268 2388 36320 2397
rect 45560 2431 45612 2440
rect 45560 2397 45569 2431
rect 45569 2397 45603 2431
rect 45603 2397 45612 2431
rect 45560 2388 45612 2397
rect 47400 2388 47452 2440
rect 49700 2388 49752 2440
rect 51540 2388 51592 2440
rect 52828 2388 52880 2440
rect 2872 2295 2924 2304
rect 2872 2261 2881 2295
rect 2881 2261 2915 2295
rect 2915 2261 2924 2295
rect 2872 2252 2924 2261
rect 29920 2320 29972 2372
rect 33968 2363 34020 2372
rect 33968 2329 33977 2363
rect 33977 2329 34011 2363
rect 34011 2329 34020 2363
rect 33968 2320 34020 2329
rect 37740 2363 37792 2372
rect 37740 2329 37749 2363
rect 37749 2329 37783 2363
rect 37783 2329 37792 2363
rect 37740 2320 37792 2329
rect 43076 2363 43128 2372
rect 43076 2329 43085 2363
rect 43085 2329 43119 2363
rect 43119 2329 43128 2363
rect 43076 2320 43128 2329
rect 52644 2363 52696 2372
rect 52644 2329 52653 2363
rect 52653 2329 52687 2363
rect 52687 2329 52696 2363
rect 52644 2320 52696 2329
rect 55588 2363 55640 2372
rect 55588 2329 55597 2363
rect 55597 2329 55631 2363
rect 55631 2329 55640 2363
rect 55588 2320 55640 2329
rect 19432 2252 19484 2304
rect 30932 2252 30984 2304
rect 46572 2252 46624 2304
rect 57888 2252 57940 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 49976 1708 50028 1760
rect 56508 1708 56560 1760
rect 52368 756 52420 808
rect 56324 756 56376 808
<< metal2 >>
rect 386 59200 442 60000
rect 1122 59200 1178 60000
rect 1950 59200 2006 60000
rect 2686 59200 2742 60000
rect 2778 59528 2834 59537
rect 2778 59463 2834 59472
rect 400 56506 428 59200
rect 388 56500 440 56506
rect 388 56442 440 56448
rect 1136 56370 1164 59200
rect 1214 58576 1270 58585
rect 1214 58511 1270 58520
rect 1124 56364 1176 56370
rect 1124 56306 1176 56312
rect 1228 56302 1256 58511
rect 1860 57316 1912 57322
rect 1860 57258 1912 57264
rect 1400 56908 1452 56914
rect 1400 56850 1452 56856
rect 1412 56681 1440 56850
rect 1398 56672 1454 56681
rect 1398 56607 1454 56616
rect 1308 56500 1360 56506
rect 1308 56442 1360 56448
rect 1216 56296 1268 56302
rect 1216 56238 1268 56244
rect 1320 37738 1348 56442
rect 1398 55856 1454 55865
rect 1398 55791 1400 55800
rect 1452 55791 1454 55800
rect 1400 55762 1452 55768
rect 1872 55758 1900 57258
rect 1964 55826 1992 59200
rect 2134 57624 2190 57633
rect 2134 57559 2190 57568
rect 2148 56914 2176 57559
rect 2136 56908 2188 56914
rect 2136 56850 2188 56856
rect 2700 56302 2728 59200
rect 2792 57526 2820 59463
rect 3514 59200 3570 60000
rect 4250 59200 4306 60000
rect 5078 59200 5134 60000
rect 5906 59200 5962 60000
rect 6642 59200 6698 60000
rect 7470 59200 7526 60000
rect 8206 59200 8262 60000
rect 9034 59200 9090 60000
rect 9770 59200 9826 60000
rect 10598 59200 10654 60000
rect 11426 59200 11482 60000
rect 12162 59200 12218 60000
rect 12990 59200 13046 60000
rect 13726 59200 13782 60000
rect 14554 59200 14610 60000
rect 15382 59200 15438 60000
rect 16118 59200 16174 60000
rect 16946 59200 17002 60000
rect 17682 59200 17738 60000
rect 18510 59200 18566 60000
rect 19246 59200 19302 60000
rect 20074 59200 20130 60000
rect 20902 59200 20958 60000
rect 21638 59200 21694 60000
rect 22466 59200 22522 60000
rect 23202 59200 23258 60000
rect 24030 59200 24086 60000
rect 24766 59200 24822 60000
rect 25594 59200 25650 60000
rect 26422 59200 26478 60000
rect 27158 59200 27214 60000
rect 27986 59200 28042 60000
rect 28722 59200 28778 60000
rect 29550 59200 29606 60000
rect 30378 59200 30434 60000
rect 31114 59200 31170 60000
rect 31942 59200 31998 60000
rect 32678 59200 32734 60000
rect 33506 59200 33562 60000
rect 34242 59200 34298 60000
rect 35070 59200 35126 60000
rect 35898 59200 35954 60000
rect 36634 59200 36690 60000
rect 37462 59200 37518 60000
rect 38198 59200 38254 60000
rect 39026 59200 39082 60000
rect 39762 59200 39818 60000
rect 40590 59200 40646 60000
rect 41418 59200 41474 60000
rect 42154 59200 42210 60000
rect 42982 59200 43038 60000
rect 43718 59200 43774 60000
rect 44546 59200 44602 60000
rect 45374 59200 45430 60000
rect 46110 59200 46166 60000
rect 46938 59200 46994 60000
rect 47674 59200 47730 60000
rect 48502 59200 48558 60000
rect 49238 59200 49294 60000
rect 50066 59200 50122 60000
rect 50894 59200 50950 60000
rect 51630 59200 51686 60000
rect 52458 59200 52514 60000
rect 53194 59200 53250 60000
rect 54022 59200 54078 60000
rect 54758 59200 54814 60000
rect 55586 59200 55642 60000
rect 56414 59200 56470 60000
rect 56506 59664 56562 59673
rect 56506 59599 56562 59608
rect 2780 57520 2832 57526
rect 2780 57462 2832 57468
rect 3148 56908 3200 56914
rect 3148 56850 3200 56856
rect 3332 56908 3384 56914
rect 3332 56850 3384 56856
rect 2688 56296 2740 56302
rect 2688 56238 2740 56244
rect 3160 55962 3188 56850
rect 3240 56704 3292 56710
rect 3240 56646 3292 56652
rect 3252 56506 3280 56646
rect 3240 56500 3292 56506
rect 3240 56442 3292 56448
rect 3344 56438 3372 56850
rect 3332 56432 3384 56438
rect 3332 56374 3384 56380
rect 3148 55956 3200 55962
rect 3148 55898 3200 55904
rect 3528 55826 3556 59200
rect 4264 57882 4292 59200
rect 4080 57854 4292 57882
rect 4080 57594 4108 57854
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4068 57588 4120 57594
rect 4068 57530 4120 57536
rect 4620 57588 4672 57594
rect 4620 57530 4672 57536
rect 4252 57384 4304 57390
rect 4252 57326 4304 57332
rect 4264 57050 4292 57326
rect 4252 57044 4304 57050
rect 4252 56986 4304 56992
rect 4632 56846 4660 57530
rect 5092 57390 5120 59200
rect 5920 57390 5948 59200
rect 6656 57458 6684 59200
rect 6644 57452 6696 57458
rect 6644 57394 6696 57400
rect 4804 57384 4856 57390
rect 4804 57326 4856 57332
rect 5080 57384 5132 57390
rect 5080 57326 5132 57332
rect 5908 57384 5960 57390
rect 5908 57326 5960 57332
rect 4620 56840 4672 56846
rect 4620 56782 4672 56788
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 4252 56432 4304 56438
rect 4252 56374 4304 56380
rect 4160 56160 4212 56166
rect 4160 56102 4212 56108
rect 4172 55962 4200 56102
rect 4160 55956 4212 55962
rect 4160 55898 4212 55904
rect 1952 55820 2004 55826
rect 1952 55762 2004 55768
rect 3516 55820 3568 55826
rect 3516 55762 3568 55768
rect 1860 55752 1912 55758
rect 1860 55694 1912 55700
rect 4264 55690 4292 56374
rect 4632 56370 4660 56782
rect 4816 56506 4844 57326
rect 7484 57322 7512 59200
rect 7472 57316 7524 57322
rect 7472 57258 7524 57264
rect 5540 57248 5592 57254
rect 5540 57190 5592 57196
rect 4804 56500 4856 56506
rect 4804 56442 4856 56448
rect 4620 56364 4672 56370
rect 4620 56306 4672 56312
rect 5264 56296 5316 56302
rect 5264 56238 5316 56244
rect 4252 55684 4304 55690
rect 4252 55626 4304 55632
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 1398 54904 1454 54913
rect 1398 54839 1454 54848
rect 1412 54738 1440 54839
rect 1400 54732 1452 54738
rect 1400 54674 1452 54680
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 1400 54120 1452 54126
rect 1400 54062 1452 54068
rect 1412 53961 1440 54062
rect 1398 53952 1454 53961
rect 1398 53887 1454 53896
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 1400 53032 1452 53038
rect 1398 53000 1400 53009
rect 1452 53000 1454 53009
rect 1398 52935 1454 52944
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 1398 52048 1454 52057
rect 1398 51983 1454 51992
rect 1412 51950 1440 51983
rect 1400 51944 1452 51950
rect 1400 51886 1452 51892
rect 1400 51468 1452 51474
rect 1400 51410 1452 51416
rect 1412 51241 1440 51410
rect 1398 51232 1454 51241
rect 1398 51167 1454 51176
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 1400 50380 1452 50386
rect 1400 50322 1452 50328
rect 1412 50289 1440 50322
rect 1398 50280 1454 50289
rect 1398 50215 1454 50224
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 1398 49328 1454 49337
rect 1398 49263 1400 49272
rect 1452 49263 1454 49272
rect 1400 49234 1452 49240
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 1398 48376 1454 48385
rect 1398 48311 1454 48320
rect 1412 48210 1440 48311
rect 1400 48204 1452 48210
rect 1400 48146 1452 48152
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 1400 47592 1452 47598
rect 1398 47560 1400 47569
rect 1452 47560 1454 47569
rect 1398 47495 1454 47504
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 1398 46608 1454 46617
rect 1398 46543 1454 46552
rect 1412 46510 1440 46543
rect 1400 46504 1452 46510
rect 1400 46446 1452 46452
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 1398 45656 1454 45665
rect 4220 45648 4516 45668
rect 1398 45591 1454 45600
rect 1412 45422 1440 45591
rect 1400 45416 1452 45422
rect 1400 45358 1452 45364
rect 1400 44940 1452 44946
rect 1400 44882 1452 44888
rect 1412 44713 1440 44882
rect 1398 44704 1454 44713
rect 1398 44639 1454 44648
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 1400 43852 1452 43858
rect 1400 43794 1452 43800
rect 1412 43761 1440 43794
rect 1398 43752 1454 43761
rect 1398 43687 1454 43696
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1412 42770 1440 42871
rect 1400 42764 1452 42770
rect 1400 42706 1452 42712
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 1400 42152 1452 42158
rect 1400 42094 1452 42100
rect 1412 41993 1440 42094
rect 1398 41984 1454 41993
rect 1398 41919 1454 41928
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 1400 41064 1452 41070
rect 1398 41032 1400 41041
rect 1452 41032 1454 41041
rect 1398 40967 1454 40976
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 1398 40080 1454 40089
rect 1398 40015 1454 40024
rect 1412 39982 1440 40015
rect 1400 39976 1452 39982
rect 1400 39918 1452 39924
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 1398 39128 1454 39137
rect 4220 39120 4516 39140
rect 1398 39063 1454 39072
rect 1412 38894 1440 39063
rect 1400 38888 1452 38894
rect 1400 38830 1452 38836
rect 1400 38412 1452 38418
rect 1400 38354 1452 38360
rect 1412 38321 1440 38354
rect 1398 38312 1454 38321
rect 1398 38247 1454 38256
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 1308 37732 1360 37738
rect 1308 37674 1360 37680
rect 1398 37360 1454 37369
rect 1398 37295 1400 37304
rect 1452 37295 1454 37304
rect 1400 37266 1452 37272
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 1398 36408 1454 36417
rect 1398 36343 1454 36352
rect 1412 36242 1440 36343
rect 1400 36236 1452 36242
rect 1400 36178 1452 36184
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 1400 35624 1452 35630
rect 1400 35566 1452 35572
rect 1412 35465 1440 35566
rect 1398 35456 1454 35465
rect 1398 35391 1454 35400
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 1398 34640 1454 34649
rect 1398 34575 1454 34584
rect 1412 34542 1440 34575
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 1398 33688 1454 33697
rect 4220 33680 4516 33700
rect 1398 33623 1454 33632
rect 1412 33454 1440 33623
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1412 32745 1440 32914
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1412 31793 1440 31826
rect 1398 31784 1454 31793
rect 1398 31719 1454 31728
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 1398 30832 1454 30841
rect 1398 30767 1400 30776
rect 1452 30767 1454 30776
rect 1400 30738 1452 30744
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 1400 30184 1452 30190
rect 1400 30126 1452 30132
rect 1412 30025 1440 30126
rect 1398 30016 1454 30025
rect 1398 29951 1454 29960
rect 1860 29708 1912 29714
rect 1860 29650 1912 29656
rect 1676 28552 1728 28558
rect 1676 28494 1728 28500
rect 1688 27674 1716 28494
rect 1872 28490 1900 29650
rect 1952 29504 2004 29510
rect 1952 29446 2004 29452
rect 1964 29073 1992 29446
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 2964 29096 3016 29102
rect 1950 29064 2006 29073
rect 2964 29038 3016 29044
rect 1950 28999 2006 29008
rect 2044 29028 2096 29034
rect 2044 28970 2096 28976
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 2056 28121 2084 28970
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2042 28112 2098 28121
rect 2608 28082 2636 28358
rect 2976 28218 3004 29038
rect 4712 28620 4764 28626
rect 4712 28562 4764 28568
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 2964 28212 3016 28218
rect 2964 28154 3016 28160
rect 2042 28047 2098 28056
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 4724 28014 4752 28562
rect 5078 28520 5134 28529
rect 5078 28455 5134 28464
rect 5092 28014 5120 28455
rect 2780 28008 2832 28014
rect 2780 27950 2832 27956
rect 4712 28008 4764 28014
rect 4712 27950 4764 27956
rect 5080 28008 5132 28014
rect 5080 27950 5132 27956
rect 1860 27940 1912 27946
rect 1860 27882 1912 27888
rect 1676 27668 1728 27674
rect 1676 27610 1728 27616
rect 1400 27328 1452 27334
rect 1400 27270 1452 27276
rect 1412 26217 1440 27270
rect 1872 27130 1900 27882
rect 1952 27872 2004 27878
rect 1952 27814 2004 27820
rect 1964 27169 1992 27814
rect 2792 27674 2820 27950
rect 2780 27668 2832 27674
rect 2780 27610 2832 27616
rect 2504 27532 2556 27538
rect 2504 27474 2556 27480
rect 3332 27532 3384 27538
rect 3332 27474 3384 27480
rect 1950 27160 2006 27169
rect 1860 27124 1912 27130
rect 1950 27095 2006 27104
rect 1860 27066 1912 27072
rect 2044 26784 2096 26790
rect 2044 26726 2096 26732
rect 2056 26450 2084 26726
rect 2516 26586 2544 27474
rect 3344 26994 3372 27474
rect 4724 27334 4752 27950
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 5080 27872 5132 27878
rect 5080 27814 5132 27820
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 4724 26926 4752 27270
rect 3424 26920 3476 26926
rect 3424 26862 3476 26868
rect 4528 26920 4580 26926
rect 4528 26862 4580 26868
rect 4712 26920 4764 26926
rect 4712 26862 4764 26868
rect 2504 26580 2556 26586
rect 2504 26522 2556 26528
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 1398 26208 1454 26217
rect 1398 26143 1454 26152
rect 3068 26042 3096 26386
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3056 26036 3108 26042
rect 3056 25978 3108 25984
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 1860 25356 1912 25362
rect 1860 25298 1912 25304
rect 1872 24954 1900 25298
rect 1952 25152 2004 25158
rect 1952 25094 2004 25100
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 1964 24449 1992 25094
rect 1950 24440 2006 24449
rect 1950 24375 2006 24384
rect 2688 24200 2740 24206
rect 2688 24142 2740 24148
rect 1860 24064 1912 24070
rect 1860 24006 1912 24012
rect 1952 24064 2004 24070
rect 1952 24006 2004 24012
rect 1584 23520 1636 23526
rect 1582 23488 1584 23497
rect 1636 23488 1638 23497
rect 1582 23423 1638 23432
rect 1872 23254 1900 24006
rect 1964 23662 1992 24006
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 1860 23248 1912 23254
rect 1860 23190 1912 23196
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 22545 1992 22918
rect 2136 22704 2188 22710
rect 2136 22646 2188 22652
rect 2044 22568 2096 22574
rect 1950 22536 2006 22545
rect 2044 22510 2096 22516
rect 1950 22471 2006 22480
rect 1950 21720 2006 21729
rect 1950 21655 1952 21664
rect 2004 21655 2006 21664
rect 1952 21626 2004 21632
rect 1952 20800 2004 20806
rect 1950 20768 1952 20777
rect 2004 20768 2006 20777
rect 1950 20703 2006 20712
rect 2056 20602 2084 22510
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 1858 19816 1914 19825
rect 1858 19751 1860 19760
rect 1912 19751 1914 19760
rect 1860 19722 1912 19728
rect 2044 18896 2096 18902
rect 2042 18864 2044 18873
rect 2096 18864 2098 18873
rect 2148 18834 2176 22646
rect 2608 22438 2636 23122
rect 2596 22432 2648 22438
rect 2596 22374 2648 22380
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2042 18799 2098 18808
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 1950 17912 2006 17921
rect 1950 17847 1952 17856
rect 2004 17847 2006 17856
rect 1952 17818 2004 17824
rect 2332 17814 2360 21830
rect 2608 21010 2636 22374
rect 2700 21690 2728 24142
rect 2884 23730 2912 25638
rect 3160 25401 3188 26182
rect 3146 25392 3202 25401
rect 3146 25327 3202 25336
rect 3332 25152 3384 25158
rect 3332 25094 3384 25100
rect 3344 24818 3372 25094
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 3148 24744 3200 24750
rect 3148 24686 3200 24692
rect 3056 24132 3108 24138
rect 3056 24074 3108 24080
rect 2964 23792 3016 23798
rect 2964 23734 3016 23740
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 2792 21078 2820 23462
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2884 21418 2912 22646
rect 2872 21412 2924 21418
rect 2872 21354 2924 21360
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2596 21004 2648 21010
rect 2596 20946 2648 20952
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2516 19514 2544 19926
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2608 19310 2636 20946
rect 2700 20806 2728 20946
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2700 20398 2728 20742
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2976 20058 3004 23734
rect 3068 21962 3096 24074
rect 3160 23322 3188 24686
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 3436 23186 3464 26862
rect 3884 26784 3936 26790
rect 3884 26726 3936 26732
rect 4160 26784 4212 26790
rect 4160 26726 4212 26732
rect 3896 25906 3924 26726
rect 4172 26330 4200 26726
rect 4540 26586 4568 26862
rect 4528 26580 4580 26586
rect 4528 26522 4580 26528
rect 4724 26450 4752 26862
rect 4712 26444 4764 26450
rect 4712 26386 4764 26392
rect 4080 26302 4200 26330
rect 4080 25974 4108 26302
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4068 25968 4120 25974
rect 4068 25910 4120 25916
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3620 25362 3648 25774
rect 3608 25356 3660 25362
rect 3608 25298 3660 25304
rect 3884 24608 3936 24614
rect 3884 24550 3936 24556
rect 3896 24274 3924 24550
rect 3884 24268 3936 24274
rect 3884 24210 3936 24216
rect 3988 24188 4016 25774
rect 4068 25696 4120 25702
rect 4068 25638 4120 25644
rect 4080 25362 4108 25638
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 4080 24886 4108 25298
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4068 24200 4120 24206
rect 3988 24160 4068 24188
rect 4068 24142 4120 24148
rect 4080 23186 4108 24142
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 4632 23730 4660 25094
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 24342 4844 24550
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4436 23656 4488 23662
rect 4436 23598 4488 23604
rect 3424 23180 3476 23186
rect 3424 23122 3476 23128
rect 4068 23180 4120 23186
rect 4068 23122 4120 23128
rect 3436 22098 3464 23122
rect 4448 23066 4476 23598
rect 4528 23588 4580 23594
rect 4528 23530 4580 23536
rect 4540 23474 4568 23530
rect 4804 23520 4856 23526
rect 4540 23446 4752 23474
rect 4804 23462 4856 23468
rect 4448 23038 4660 23066
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3056 21956 3108 21962
rect 3056 21898 3108 21904
rect 3436 21554 3464 22034
rect 3424 21548 3476 21554
rect 3424 21490 3476 21496
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2964 19780 3016 19786
rect 2964 19722 3016 19728
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 1768 17604 1820 17610
rect 1768 17546 1820 17552
rect 1780 6914 1808 17546
rect 2042 17096 2098 17105
rect 2042 17031 2044 17040
rect 2096 17031 2098 17040
rect 2044 17002 2096 17008
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1872 8022 1900 16730
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2042 16144 2098 16153
rect 2042 16079 2044 16088
rect 2096 16079 2098 16088
rect 2044 16050 2096 16056
rect 1950 15192 2006 15201
rect 1950 15127 1952 15136
rect 2004 15127 2006 15136
rect 1952 15098 2004 15104
rect 1952 14272 2004 14278
rect 1950 14240 1952 14249
rect 2004 14240 2006 14249
rect 1950 14175 2006 14184
rect 2042 13288 2098 13297
rect 2042 13223 2044 13232
rect 2096 13223 2098 13232
rect 2044 13194 2096 13200
rect 1950 12472 2006 12481
rect 1950 12407 1952 12416
rect 2004 12407 2006 12416
rect 1952 12378 2004 12384
rect 1952 11552 2004 11558
rect 1950 11520 1952 11529
rect 2004 11520 2006 11529
rect 1950 11455 2006 11464
rect 2042 10568 2098 10577
rect 2042 10503 2044 10512
rect 2096 10503 2098 10512
rect 2044 10474 2096 10480
rect 2044 9648 2096 9654
rect 2042 9616 2044 9625
rect 2096 9616 2098 9625
rect 2042 9551 2098 9560
rect 1952 8832 2004 8838
rect 1950 8800 1952 8809
rect 2004 8800 2006 8809
rect 1950 8735 2006 8744
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 2042 7848 2098 7857
rect 2042 7783 2044 7792
rect 2096 7783 2098 7792
rect 2044 7754 2096 7760
rect 1780 6886 1900 6914
rect 1872 5846 1900 6886
rect 2042 6896 2098 6905
rect 2042 6831 2098 6840
rect 2056 6798 2084 6831
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 1950 5944 2006 5953
rect 1950 5879 1952 5888
rect 2004 5879 2006 5888
rect 1952 5850 2004 5856
rect 1860 5840 1912 5846
rect 1860 5782 1912 5788
rect 2148 5166 2176 16662
rect 2976 9110 3004 19722
rect 3068 18970 3096 20266
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3160 18834 3188 19178
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3436 18766 3464 21354
rect 3528 21146 3556 22510
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 4080 21554 4108 21966
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4068 21412 4120 21418
rect 4068 21354 4120 21360
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3792 20936 3844 20942
rect 3792 20878 3844 20884
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3620 10606 3648 20266
rect 3804 19310 3832 20878
rect 3792 19304 3844 19310
rect 3792 19246 3844 19252
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 4080 9518 4108 21354
rect 4632 20874 4660 23038
rect 4724 21146 4752 23446
rect 4816 23254 4844 23462
rect 4804 23248 4856 23254
rect 4804 23190 4856 23196
rect 4908 22642 4936 27814
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 5000 23662 5028 24686
rect 5092 24410 5120 27814
rect 5276 26926 5304 56238
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 5460 27130 5488 27542
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5448 26988 5500 26994
rect 5448 26930 5500 26936
rect 5264 26920 5316 26926
rect 5264 26862 5316 26868
rect 5356 26852 5408 26858
rect 5356 26794 5408 26800
rect 5368 26450 5396 26794
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5172 25764 5224 25770
rect 5172 25706 5224 25712
rect 5184 25498 5212 25706
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5276 24750 5304 25298
rect 5264 24744 5316 24750
rect 5264 24686 5316 24692
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5276 24342 5304 24550
rect 5264 24336 5316 24342
rect 5264 24278 5316 24284
rect 4988 23656 5040 23662
rect 4988 23598 5040 23604
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4988 22500 5040 22506
rect 4988 22442 5040 22448
rect 4816 21690 4844 22442
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4804 21344 4856 21350
rect 4804 21286 4856 21292
rect 4816 21146 4844 21286
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4632 19258 4660 19926
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4540 19230 4660 19258
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4540 19174 4568 19230
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4724 18970 4752 19246
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 1952 5024 2004 5030
rect 1950 4992 1952 5001
rect 2004 4992 2006 5001
rect 1950 4927 2006 4936
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 2042 4176 2098 4185
rect 2042 4111 2044 4120
rect 2096 4111 2098 4120
rect 2044 4082 2096 4088
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 800 1440 2790
rect 1688 2514 1716 3130
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1964 2281 1992 3334
rect 2056 3194 2084 3334
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1950 2272 2006 2281
rect 1950 2207 2006 2216
rect 2332 800 2360 3538
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 3054 3224 3110 3233
rect 4220 3216 4516 3236
rect 3054 3159 3056 3168
rect 3108 3159 3110 3168
rect 3056 3130 3108 3136
rect 4724 3126 4752 16050
rect 4816 11694 4844 19790
rect 4908 12374 4936 21898
rect 5000 16114 5028 22442
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5092 19514 5120 20334
rect 5080 19508 5132 19514
rect 5080 19450 5132 19456
rect 5276 19242 5304 24278
rect 5460 22506 5488 26930
rect 5448 22500 5500 22506
rect 5448 22442 5500 22448
rect 5552 22098 5580 57190
rect 8220 56914 8248 59200
rect 9048 57390 9076 59200
rect 9784 57390 9812 59200
rect 9036 57384 9088 57390
rect 9036 57326 9088 57332
rect 9772 57384 9824 57390
rect 9772 57326 9824 57332
rect 8300 56976 8352 56982
rect 8300 56918 8352 56924
rect 8208 56908 8260 56914
rect 8208 56850 8260 56856
rect 8312 54806 8340 56918
rect 10612 56914 10640 59200
rect 11440 57390 11468 59200
rect 12176 57526 12204 59200
rect 11980 57520 12032 57526
rect 11980 57462 12032 57468
rect 12164 57520 12216 57526
rect 12164 57462 12216 57468
rect 11428 57384 11480 57390
rect 11428 57326 11480 57332
rect 11796 57316 11848 57322
rect 11796 57258 11848 57264
rect 11060 57248 11112 57254
rect 11060 57190 11112 57196
rect 11244 57248 11296 57254
rect 11244 57190 11296 57196
rect 10600 56908 10652 56914
rect 10600 56850 10652 56856
rect 11072 56846 11100 57190
rect 11060 56840 11112 56846
rect 11060 56782 11112 56788
rect 11256 56302 11284 57190
rect 11808 56846 11836 57258
rect 11992 56914 12020 57462
rect 12256 57384 12308 57390
rect 12256 57326 12308 57332
rect 12268 56982 12296 57326
rect 12440 57248 12492 57254
rect 12440 57190 12492 57196
rect 12256 56976 12308 56982
rect 12256 56918 12308 56924
rect 11980 56908 12032 56914
rect 11980 56850 12032 56856
rect 11796 56840 11848 56846
rect 11796 56782 11848 56788
rect 11808 56438 11836 56782
rect 11796 56432 11848 56438
rect 11796 56374 11848 56380
rect 11992 56370 12020 56850
rect 12164 56840 12216 56846
rect 12164 56782 12216 56788
rect 11980 56364 12032 56370
rect 11980 56306 12032 56312
rect 11244 56296 11296 56302
rect 11244 56238 11296 56244
rect 12072 56296 12124 56302
rect 12072 56238 12124 56244
rect 8300 54800 8352 54806
rect 8300 54742 8352 54748
rect 8312 53990 8340 54742
rect 8300 53984 8352 53990
rect 8300 53926 8352 53932
rect 8852 53984 8904 53990
rect 8852 53926 8904 53932
rect 8760 30592 8812 30598
rect 8760 30534 8812 30540
rect 6460 29708 6512 29714
rect 6460 29650 6512 29656
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 7288 29708 7340 29714
rect 7288 29650 7340 29656
rect 8208 29708 8260 29714
rect 8208 29650 8260 29656
rect 5816 28960 5868 28966
rect 5816 28902 5868 28908
rect 5828 28694 5856 28902
rect 6472 28762 6500 29650
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 7104 29504 7156 29510
rect 7104 29446 7156 29452
rect 6460 28756 6512 28762
rect 6460 28698 6512 28704
rect 5816 28688 5868 28694
rect 5816 28630 5868 28636
rect 6564 27946 6592 29446
rect 7116 29102 7144 29446
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 7104 29096 7156 29102
rect 7104 29038 7156 29044
rect 6840 28626 6868 29038
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 6828 28620 6880 28626
rect 6828 28562 6880 28568
rect 6552 27940 6604 27946
rect 6552 27882 6604 27888
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 5644 27130 5672 27406
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 6184 26444 6236 26450
rect 6184 26386 6236 26392
rect 6196 26042 6224 26386
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6184 26036 6236 26042
rect 6184 25978 6236 25984
rect 6000 25356 6052 25362
rect 6000 25298 6052 25304
rect 6184 25356 6236 25362
rect 6288 25344 6316 26182
rect 6236 25316 6316 25344
rect 6184 25298 6236 25304
rect 5632 24744 5684 24750
rect 5632 24686 5684 24692
rect 5644 24410 5672 24686
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 6012 23730 6040 25298
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 6104 24410 6132 24618
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 5908 23656 5960 23662
rect 5908 23598 5960 23604
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5736 22574 5764 22918
rect 5724 22568 5776 22574
rect 5724 22510 5776 22516
rect 5920 22438 5948 23598
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 6000 22092 6052 22098
rect 6000 22034 6052 22040
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5460 21010 5488 21626
rect 6012 21622 6040 22034
rect 6000 21616 6052 21622
rect 6000 21558 6052 21564
rect 5632 21480 5684 21486
rect 5632 21422 5684 21428
rect 5644 21078 5672 21422
rect 5632 21072 5684 21078
rect 5632 21014 5684 21020
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 5644 20330 5672 20742
rect 6012 20534 6040 21558
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5632 20324 5684 20330
rect 5632 20266 5684 20272
rect 5368 19310 5396 20266
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 5460 19446 5488 20198
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5264 19236 5316 19242
rect 5264 19178 5316 19184
rect 5552 17134 5580 20198
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5644 19174 5672 19790
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5736 18426 5764 19858
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5828 16046 5856 19654
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5920 18222 5948 18838
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6104 18426 6132 18770
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6196 18290 6224 25298
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 6380 24274 6408 24346
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 23730 6408 24210
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6288 18834 6316 22374
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6380 21010 6408 21422
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 18970 6408 19722
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 4896 12368 4948 12374
rect 4896 12310 4948 12316
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2792 1329 2820 2858
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2778 1320 2834 1329
rect 2778 1255 2834 1264
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2884 513 2912 2246
rect 3252 800 3280 2858
rect 6472 2854 6500 27406
rect 6840 26994 6868 28562
rect 6932 28218 6960 28970
rect 7208 28762 7236 29650
rect 7300 29034 7328 29650
rect 8116 29504 8168 29510
rect 8116 29446 8168 29452
rect 7288 29028 7340 29034
rect 7288 28970 7340 28976
rect 8128 28994 8156 29446
rect 8220 29306 8248 29650
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 8772 29170 8800 30534
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 7300 28626 7328 28970
rect 8128 28966 8248 28994
rect 8220 28626 8248 28966
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 6920 28212 6972 28218
rect 6920 28154 6972 28160
rect 7024 27674 7052 28562
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7012 27668 7064 27674
rect 7012 27610 7064 27616
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6748 25838 6776 26182
rect 6736 25832 6788 25838
rect 6736 25774 6788 25780
rect 6840 25684 6868 26930
rect 7116 26926 7144 28358
rect 7300 27334 7328 28562
rect 7564 28552 7616 28558
rect 8220 28529 8248 28562
rect 7564 28494 7616 28500
rect 8206 28520 8262 28529
rect 7472 28008 7524 28014
rect 7576 27996 7604 28494
rect 8206 28455 8262 28464
rect 8116 28416 8168 28422
rect 8116 28358 8168 28364
rect 8128 28082 8156 28358
rect 8116 28076 8168 28082
rect 8116 28018 8168 28024
rect 7524 27968 7604 27996
rect 7472 27950 7524 27956
rect 7576 27538 7604 27968
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 7748 27532 7800 27538
rect 7748 27474 7800 27480
rect 7288 27328 7340 27334
rect 7288 27270 7340 27276
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 7472 26784 7524 26790
rect 7472 26726 7524 26732
rect 7484 26450 7512 26726
rect 7576 26466 7604 27474
rect 7760 26586 7788 27474
rect 8128 27470 8156 28018
rect 8668 28008 8720 28014
rect 8772 27996 8800 29106
rect 8720 27968 8800 27996
rect 8668 27950 8720 27956
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 8128 27062 8156 27406
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 7012 26444 7064 26450
rect 7012 26386 7064 26392
rect 7472 26444 7524 26450
rect 7576 26438 7880 26466
rect 7472 26386 7524 26392
rect 6748 25656 6868 25684
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6564 24070 6592 25094
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6564 23866 6592 24006
rect 6552 23860 6604 23866
rect 6748 23848 6776 25656
rect 6932 25498 6960 26386
rect 6828 25492 6880 25498
rect 6828 25434 6880 25440
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6840 25158 6868 25434
rect 7024 25294 7052 26386
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 25770 7236 26250
rect 7564 26036 7616 26042
rect 7564 25978 7616 25984
rect 7196 25764 7248 25770
rect 7196 25706 7248 25712
rect 7576 25430 7604 25978
rect 7656 25764 7708 25770
rect 7656 25706 7708 25712
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 6828 25152 6880 25158
rect 6828 25094 6880 25100
rect 7024 24698 7052 25230
rect 7668 25158 7696 25706
rect 7852 25430 7880 26438
rect 7944 25838 7972 26930
rect 8116 26852 8168 26858
rect 8116 26794 8168 26800
rect 7932 25832 7984 25838
rect 7932 25774 7984 25780
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7024 24670 7236 24698
rect 7944 24682 7972 25094
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6828 23860 6880 23866
rect 6748 23820 6828 23848
rect 6552 23802 6604 23808
rect 6828 23802 6880 23808
rect 6840 23662 6868 23802
rect 6828 23656 6880 23662
rect 6828 23598 6880 23604
rect 6932 23186 6960 24006
rect 7012 23588 7064 23594
rect 7012 23530 7064 23536
rect 7024 23322 7052 23530
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6736 22160 6788 22166
rect 6736 22102 6788 22108
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6656 21554 6684 22034
rect 6748 21690 6776 22102
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6932 18970 6960 22714
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 7024 19514 7052 20266
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7116 19394 7144 24550
rect 7208 23186 7236 24670
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 7470 24304 7526 24313
rect 7470 24239 7472 24248
rect 7524 24239 7526 24248
rect 7564 24268 7616 24274
rect 7472 24210 7524 24216
rect 7564 24210 7616 24216
rect 7576 23594 7604 24210
rect 7944 24138 7972 24618
rect 8036 24614 8064 25298
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 8024 24268 8076 24274
rect 8024 24210 8076 24216
rect 7932 24132 7984 24138
rect 7932 24074 7984 24080
rect 7564 23588 7616 23594
rect 7564 23530 7616 23536
rect 7840 23520 7892 23526
rect 7840 23462 7892 23468
rect 7852 23186 7880 23462
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7288 22432 7340 22438
rect 7288 22374 7340 22380
rect 7196 21072 7248 21078
rect 7196 21014 7248 21020
rect 7208 20602 7236 21014
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7300 19854 7328 22374
rect 7484 22094 7512 22510
rect 7564 22094 7616 22098
rect 7484 22092 7616 22094
rect 7484 22066 7564 22092
rect 7564 22034 7616 22040
rect 7576 21554 7604 22034
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7944 21486 7972 23054
rect 8036 22982 8064 24210
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7024 19366 7144 19394
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7024 18834 7052 19366
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7392 14958 7420 20878
rect 7564 20324 7616 20330
rect 7564 20266 7616 20272
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7484 13462 7512 19790
rect 7576 14550 7604 20266
rect 7944 20058 7972 21286
rect 8036 20330 8064 22918
rect 8128 22438 8156 26794
rect 8220 26382 8248 27270
rect 8404 26926 8432 27474
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8404 25294 8432 26862
rect 8496 26586 8524 27882
rect 8576 26852 8628 26858
rect 8576 26794 8628 26800
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8484 25968 8536 25974
rect 8484 25910 8536 25916
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8496 24970 8524 25910
rect 8312 24942 8524 24970
rect 8312 24886 8340 24942
rect 8300 24880 8352 24886
rect 8300 24822 8352 24828
rect 8208 24744 8260 24750
rect 8484 24744 8536 24750
rect 8260 24704 8340 24732
rect 8208 24686 8260 24692
rect 8312 24614 8340 24704
rect 8484 24686 8536 24692
rect 8300 24608 8352 24614
rect 8300 24550 8352 24556
rect 8496 24410 8524 24686
rect 8588 24614 8616 26794
rect 8680 25838 8708 27950
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8116 22432 8168 22438
rect 8116 22374 8168 22380
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 18970 8064 19178
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8128 18834 8156 22374
rect 8220 22166 8248 23734
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21554 8248 21830
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8220 21010 8248 21490
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7472 13456 7524 13462
rect 7472 13398 7524 13404
rect 7852 3670 7880 18226
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 8312 3398 8340 24210
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8404 21010 8432 24006
rect 8496 23662 8524 24346
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8588 22982 8616 24550
rect 8680 24138 8708 25774
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8680 23866 8708 24074
rect 8864 23866 8892 53926
rect 11888 53236 11940 53242
rect 11888 53178 11940 53184
rect 11428 30932 11480 30938
rect 11428 30874 11480 30880
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9416 28422 9444 29650
rect 9600 29646 9628 29990
rect 9588 29640 9640 29646
rect 9588 29582 9640 29588
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 29102 9536 29446
rect 9496 29096 9548 29102
rect 9496 29038 9548 29044
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9600 28234 9628 29582
rect 9772 28960 9824 28966
rect 9772 28902 9824 28908
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 9678 28792 9734 28801
rect 9678 28727 9680 28736
rect 9732 28727 9734 28736
rect 9680 28698 9732 28704
rect 9784 28490 9812 28902
rect 10152 28626 10180 28902
rect 9956 28620 10008 28626
rect 10140 28620 10192 28626
rect 10008 28580 10088 28608
rect 9956 28562 10008 28568
rect 9772 28484 9824 28490
rect 9772 28426 9824 28432
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9600 28206 9904 28234
rect 9588 28076 9640 28082
rect 9508 28036 9588 28064
rect 9508 27606 9536 28036
rect 9588 28018 9640 28024
rect 9876 27606 9904 28206
rect 9496 27600 9548 27606
rect 9496 27542 9548 27548
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9692 27334 9720 27474
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 9508 26518 9536 27270
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9496 26512 9548 26518
rect 9496 26454 9548 26460
rect 9692 26246 9720 26522
rect 9680 26240 9732 26246
rect 9680 26182 9732 26188
rect 9784 25430 9812 27474
rect 9876 26994 9904 27542
rect 9968 27470 9996 28358
rect 10060 27946 10088 28580
rect 10140 28562 10192 28568
rect 10048 27940 10100 27946
rect 10048 27882 10100 27888
rect 10048 27532 10100 27538
rect 10048 27474 10100 27480
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 27062 9996 27406
rect 9956 27056 10008 27062
rect 9956 26998 10008 27004
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9864 26444 9916 26450
rect 9864 26386 9916 26392
rect 9876 25702 9904 26386
rect 10060 26246 10088 27474
rect 10428 27130 10456 30534
rect 10520 30394 10548 30738
rect 10508 30388 10560 30394
rect 10508 30330 10560 30336
rect 11440 30258 11468 30874
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 11428 30252 11480 30258
rect 11428 30194 11480 30200
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10138 27024 10194 27033
rect 10138 26959 10194 26968
rect 10152 26926 10180 26959
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10416 26920 10468 26926
rect 10416 26862 10468 26868
rect 10232 26852 10284 26858
rect 10232 26794 10284 26800
rect 10244 26382 10272 26794
rect 10428 26450 10456 26862
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25974 10088 26182
rect 10048 25968 10100 25974
rect 10048 25910 10100 25916
rect 10336 25770 10364 26386
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10520 25838 10548 26182
rect 10612 25838 10640 27814
rect 10704 27033 10732 28494
rect 10980 27606 11008 30126
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29850 11100 29990
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 11072 28694 11100 29650
rect 11532 29306 11560 30670
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11060 28688 11112 28694
rect 11060 28630 11112 28636
rect 11164 28014 11192 29106
rect 11532 28626 11560 29242
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11520 28620 11572 28626
rect 11520 28562 11572 28568
rect 11244 28144 11296 28150
rect 11244 28086 11296 28092
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 11152 27532 11204 27538
rect 11152 27474 11204 27480
rect 10968 27328 11020 27334
rect 11020 27276 11100 27282
rect 10968 27270 11100 27276
rect 10980 27254 11100 27270
rect 10690 27024 10746 27033
rect 10690 26959 10746 26968
rect 10968 26920 11020 26926
rect 10888 26880 10968 26908
rect 10888 26586 10916 26880
rect 10968 26862 11020 26868
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10782 26480 10838 26489
rect 10782 26415 10784 26424
rect 10836 26415 10838 26424
rect 10784 26386 10836 26392
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10324 25764 10376 25770
rect 10324 25706 10376 25712
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9772 25424 9824 25430
rect 9772 25366 9824 25372
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9600 24954 9628 25298
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9600 24177 9628 24278
rect 9586 24168 9642 24177
rect 9586 24103 9642 24112
rect 8668 23860 8720 23866
rect 8668 23802 8720 23808
rect 8852 23860 8904 23866
rect 8852 23802 8904 23808
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8484 22636 8536 22642
rect 8680 22624 8708 23802
rect 8536 22596 8708 22624
rect 8484 22578 8536 22584
rect 8496 21010 8524 22578
rect 8852 21888 8904 21894
rect 8852 21830 8904 21836
rect 8864 21486 8892 21830
rect 8576 21480 8628 21486
rect 8576 21422 8628 21428
rect 8852 21480 8904 21486
rect 8852 21422 8904 21428
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8496 19922 8524 20334
rect 8588 19922 8616 21422
rect 9140 20398 9168 23802
rect 9692 23662 9720 24550
rect 9876 23866 9904 25638
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10416 24744 10468 24750
rect 10416 24686 10468 24692
rect 10692 24744 10744 24750
rect 10692 24686 10744 24692
rect 10152 24449 10180 24686
rect 10138 24440 10194 24449
rect 10428 24410 10456 24686
rect 10138 24375 10194 24384
rect 10416 24404 10468 24410
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9692 23186 9720 23598
rect 10152 23322 10180 24375
rect 10416 24346 10468 24352
rect 10704 24070 10732 24686
rect 10796 24449 10824 26386
rect 11072 25922 11100 27254
rect 11164 27130 11192 27474
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11256 27062 11284 28086
rect 11244 27056 11296 27062
rect 11244 26998 11296 27004
rect 11256 26586 11284 26998
rect 11348 26790 11376 28562
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11440 28150 11468 28494
rect 11428 28144 11480 28150
rect 11428 28086 11480 28092
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11612 27056 11664 27062
rect 11612 26998 11664 27004
rect 11428 26852 11480 26858
rect 11428 26794 11480 26800
rect 11336 26784 11388 26790
rect 11336 26726 11388 26732
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11152 26444 11204 26450
rect 11256 26432 11284 26522
rect 11204 26404 11284 26432
rect 11152 26386 11204 26392
rect 11348 26382 11376 26726
rect 11440 26450 11468 26794
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11520 26444 11572 26450
rect 11520 26386 11572 26392
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11072 25894 11192 25922
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 11072 25158 11100 25774
rect 11164 25158 11192 25894
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10782 24440 10838 24449
rect 10782 24375 10838 24384
rect 10888 24342 10916 24550
rect 10980 24342 11008 24754
rect 10876 24336 10928 24342
rect 10876 24278 10928 24284
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 10784 24268 10836 24274
rect 10784 24210 10836 24216
rect 10692 24064 10744 24070
rect 10796 24041 10824 24210
rect 10692 24006 10744 24012
rect 10782 24032 10838 24041
rect 10782 23967 10838 23976
rect 10980 23322 11008 24278
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 9680 23180 9732 23186
rect 9680 23122 9732 23128
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 9692 22098 9720 23122
rect 10336 22574 10364 23122
rect 10508 22704 10560 22710
rect 10560 22664 10824 22692
rect 10508 22646 10560 22652
rect 10796 22574 10824 22664
rect 10980 22642 11008 23258
rect 11072 22642 11100 25094
rect 11532 24886 11560 26386
rect 11520 24880 11572 24886
rect 11520 24822 11572 24828
rect 11152 24676 11204 24682
rect 11152 24618 11204 24624
rect 11520 24676 11572 24682
rect 11520 24618 11572 24624
rect 11164 23322 11192 24618
rect 11334 24440 11390 24449
rect 11334 24375 11390 24384
rect 11348 24274 11376 24375
rect 11532 24274 11560 24618
rect 11336 24268 11388 24274
rect 11336 24210 11388 24216
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11624 24206 11652 26998
rect 11704 26240 11756 26246
rect 11704 26182 11756 26188
rect 11716 25430 11744 26182
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11808 24682 11836 27950
rect 11796 24676 11848 24682
rect 11796 24618 11848 24624
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11244 23792 11296 23798
rect 11296 23740 11376 23746
rect 11244 23734 11376 23740
rect 11256 23718 11376 23734
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11164 23186 11192 23258
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 10968 22636 11020 22642
rect 10968 22578 11020 22584
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10324 22568 10376 22574
rect 10324 22510 10376 22516
rect 10416 22568 10468 22574
rect 10416 22510 10468 22516
rect 10784 22568 10836 22574
rect 10784 22510 10836 22516
rect 10060 22098 10088 22510
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10336 22098 10364 22170
rect 10428 22166 10456 22510
rect 10980 22234 11008 22578
rect 10968 22228 11020 22234
rect 10968 22170 11020 22176
rect 11164 22166 11192 23122
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 11256 22098 11284 22918
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 10048 22094 10100 22098
rect 10048 22092 10180 22094
rect 10100 22066 10180 22092
rect 10048 22034 10100 22040
rect 10152 21486 10180 22066
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 10152 20398 10180 21422
rect 10324 21412 10376 21418
rect 10324 21354 10376 21360
rect 10336 20602 10364 21354
rect 10520 21350 10548 22034
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10336 20398 10364 20538
rect 10612 20466 10640 21558
rect 11348 21486 11376 23718
rect 11808 23186 11836 24618
rect 11900 23798 11928 53178
rect 12084 31890 12112 56238
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 12084 31482 12112 31826
rect 12176 31754 12204 56782
rect 12256 39840 12308 39846
rect 12256 39782 12308 39788
rect 12268 39574 12296 39782
rect 12256 39568 12308 39574
rect 12256 39510 12308 39516
rect 12452 31958 12480 57190
rect 13004 56982 13032 59200
rect 13740 57372 13768 59200
rect 14568 57458 14596 59200
rect 15396 57458 15424 59200
rect 14556 57452 14608 57458
rect 14556 57394 14608 57400
rect 15384 57452 15436 57458
rect 15384 57394 15436 57400
rect 13820 57384 13872 57390
rect 13740 57344 13820 57372
rect 13820 57326 13872 57332
rect 13636 57248 13688 57254
rect 13636 57190 13688 57196
rect 15108 57248 15160 57254
rect 15108 57190 15160 57196
rect 15568 57248 15620 57254
rect 15568 57190 15620 57196
rect 15660 57248 15712 57254
rect 15660 57190 15712 57196
rect 12992 56976 13044 56982
rect 12992 56918 13044 56924
rect 13176 56772 13228 56778
rect 13176 56714 13228 56720
rect 12716 56228 12768 56234
rect 12716 56170 12768 56176
rect 12624 39976 12676 39982
rect 12624 39918 12676 39924
rect 12636 39642 12664 39918
rect 12624 39636 12676 39642
rect 12624 39578 12676 39584
rect 12532 38752 12584 38758
rect 12532 38694 12584 38700
rect 12544 38486 12572 38694
rect 12532 38480 12584 38486
rect 12532 38422 12584 38428
rect 12440 31952 12492 31958
rect 12440 31894 12492 31900
rect 12176 31726 12388 31754
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 12256 31476 12308 31482
rect 12256 31418 12308 31424
rect 12268 30666 12296 31418
rect 12360 31278 12388 31726
rect 12348 31272 12400 31278
rect 12348 31214 12400 31220
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 12084 29102 12112 29446
rect 12268 29306 12296 30194
rect 12360 29782 12388 31214
rect 12452 30870 12480 31894
rect 12624 31680 12676 31686
rect 12624 31622 12676 31628
rect 12636 31414 12664 31622
rect 12624 31408 12676 31414
rect 12624 31350 12676 31356
rect 12440 30864 12492 30870
rect 12440 30806 12492 30812
rect 12452 30190 12480 30806
rect 12532 30728 12584 30734
rect 12532 30670 12584 30676
rect 12544 30326 12572 30670
rect 12532 30320 12584 30326
rect 12532 30262 12584 30268
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12348 29776 12400 29782
rect 12348 29718 12400 29724
rect 12544 29714 12572 30262
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12072 29096 12124 29102
rect 12072 29038 12124 29044
rect 12268 28762 12296 29242
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 12636 28558 12664 29514
rect 12728 28626 12756 56170
rect 13188 35034 13216 56714
rect 13360 55956 13412 55962
rect 13360 55898 13412 55904
rect 13268 39976 13320 39982
rect 13268 39918 13320 39924
rect 13280 39438 13308 39918
rect 13268 39432 13320 39438
rect 13268 39374 13320 39380
rect 13280 38894 13308 39374
rect 13268 38888 13320 38894
rect 13268 38830 13320 38836
rect 13280 38554 13308 38830
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 13188 35006 13308 35034
rect 13176 32292 13228 32298
rect 13176 32234 13228 32240
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12912 30734 12940 31758
rect 13188 31210 13216 32234
rect 13280 31890 13308 35006
rect 13372 32366 13400 55898
rect 13452 39908 13504 39914
rect 13452 39850 13504 39856
rect 13464 39642 13492 39850
rect 13452 39636 13504 39642
rect 13452 39578 13504 39584
rect 13464 38894 13492 39578
rect 13452 38888 13504 38894
rect 13452 38830 13504 38836
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 13268 31884 13320 31890
rect 13268 31826 13320 31832
rect 13280 31346 13308 31826
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13268 31340 13320 31346
rect 13268 31282 13320 31288
rect 13176 31204 13228 31210
rect 13176 31146 13228 31152
rect 12992 30796 13044 30802
rect 12992 30738 13044 30744
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12808 30592 12860 30598
rect 12808 30534 12860 30540
rect 12820 30394 12848 30534
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12820 29714 12848 30330
rect 12912 30326 12940 30670
rect 12900 30320 12952 30326
rect 12900 30262 12952 30268
rect 12808 29708 12860 29714
rect 12808 29650 12860 29656
rect 12912 29646 12940 30262
rect 12900 29640 12952 29646
rect 12900 29582 12952 29588
rect 12912 28694 12940 29582
rect 13004 29238 13032 30738
rect 13188 30190 13216 31146
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 13360 30048 13412 30054
rect 13360 29990 13412 29996
rect 12992 29232 13044 29238
rect 12992 29174 13044 29180
rect 12900 28688 12952 28694
rect 12900 28630 12952 28636
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 13004 28082 13032 29174
rect 13096 29102 13124 29990
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 13268 28416 13320 28422
rect 13268 28358 13320 28364
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 13176 28008 13228 28014
rect 13176 27950 13228 27956
rect 11978 26480 12034 26489
rect 11978 26415 11980 26424
rect 12032 26415 12034 26424
rect 11980 26386 12032 26392
rect 12084 24818 12112 27950
rect 12440 27668 12492 27674
rect 12440 27610 12492 27616
rect 12256 27328 12308 27334
rect 12254 27296 12256 27305
rect 12348 27328 12400 27334
rect 12308 27296 12310 27305
rect 12348 27270 12400 27276
rect 12254 27231 12310 27240
rect 12360 26994 12388 27270
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12452 26926 12480 27610
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12532 27396 12584 27402
rect 12532 27338 12584 27344
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12452 26586 12480 26862
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12360 26450 12388 26522
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12440 26444 12492 26450
rect 12544 26432 12572 27338
rect 12636 26994 12664 27406
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12636 26790 12664 26930
rect 12716 26920 12768 26926
rect 12714 26888 12716 26897
rect 12768 26888 12770 26897
rect 12714 26823 12770 26832
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12624 26580 12676 26586
rect 12624 26522 12676 26528
rect 12492 26404 12572 26432
rect 12440 26386 12492 26392
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12176 24886 12204 25094
rect 12164 24880 12216 24886
rect 12164 24822 12216 24828
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12440 24336 12492 24342
rect 12440 24278 12492 24284
rect 11980 24268 12032 24274
rect 11980 24210 12032 24216
rect 11992 23866 12020 24210
rect 12348 24200 12400 24206
rect 12452 24177 12480 24278
rect 12636 24274 12664 26522
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12728 25702 12756 26386
rect 12900 26240 12952 26246
rect 12900 26182 12952 26188
rect 12912 25838 12940 26182
rect 12900 25832 12952 25838
rect 12900 25774 12952 25780
rect 12716 25696 12768 25702
rect 12716 25638 12768 25644
rect 12728 25362 12756 25638
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12808 24744 12860 24750
rect 13004 24698 13032 26726
rect 13188 26382 13216 27950
rect 13280 26772 13308 28358
rect 13372 26926 13400 29990
rect 13464 28694 13492 31622
rect 13648 31278 13676 57190
rect 15120 56846 15148 57190
rect 15580 56982 15608 57190
rect 15568 56976 15620 56982
rect 15568 56918 15620 56924
rect 15672 56914 15700 57190
rect 16132 56914 16160 59200
rect 16960 57390 16988 59200
rect 16948 57384 17000 57390
rect 17696 57372 17724 59200
rect 18524 57390 18552 59200
rect 17960 57384 18012 57390
rect 17696 57344 17960 57372
rect 16948 57326 17000 57332
rect 17960 57326 18012 57332
rect 18512 57384 18564 57390
rect 19260 57372 19288 59200
rect 20088 57458 20116 59200
rect 20916 57458 20944 59200
rect 20076 57452 20128 57458
rect 20076 57394 20128 57400
rect 20904 57452 20956 57458
rect 20904 57394 20956 57400
rect 19340 57384 19392 57390
rect 19260 57344 19340 57372
rect 18512 57326 18564 57332
rect 21652 57372 21680 59200
rect 22100 57384 22152 57390
rect 21652 57344 22100 57372
rect 19340 57326 19392 57332
rect 22100 57326 22152 57332
rect 20168 57316 20220 57322
rect 20168 57258 20220 57264
rect 17960 57248 18012 57254
rect 17960 57190 18012 57196
rect 18236 57248 18288 57254
rect 18236 57190 18288 57196
rect 18880 57248 18932 57254
rect 18880 57190 18932 57196
rect 15660 56908 15712 56914
rect 15660 56850 15712 56856
rect 16120 56908 16172 56914
rect 16120 56850 16172 56856
rect 17972 56846 18000 57190
rect 18248 56982 18276 57190
rect 18236 56976 18288 56982
rect 18236 56918 18288 56924
rect 18892 56914 18920 57190
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 18880 56908 18932 56914
rect 18880 56850 18932 56856
rect 20180 56846 20208 57258
rect 20260 57248 20312 57254
rect 20260 57190 20312 57196
rect 20352 57248 20404 57254
rect 20352 57190 20404 57196
rect 21548 57248 21600 57254
rect 21548 57190 21600 57196
rect 15108 56840 15160 56846
rect 15108 56782 15160 56788
rect 17960 56840 18012 56846
rect 17960 56782 18012 56788
rect 20168 56840 20220 56846
rect 20168 56782 20220 56788
rect 20272 56778 20300 57190
rect 20364 56846 20392 57190
rect 21560 56982 21588 57190
rect 21548 56976 21600 56982
rect 21548 56918 21600 56924
rect 22480 56914 22508 59200
rect 23020 57316 23072 57322
rect 23020 57258 23072 57264
rect 22468 56908 22520 56914
rect 22468 56850 22520 56856
rect 23032 56846 23060 57258
rect 20352 56840 20404 56846
rect 20352 56782 20404 56788
rect 23020 56840 23072 56846
rect 23020 56782 23072 56788
rect 20260 56772 20312 56778
rect 20260 56714 20312 56720
rect 23112 56704 23164 56710
rect 23112 56646 23164 56652
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 22836 55344 22888 55350
rect 22836 55286 22888 55292
rect 22560 55072 22612 55078
rect 22560 55014 22612 55020
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 22572 54806 22600 55014
rect 22560 54800 22612 54806
rect 22560 54742 22612 54748
rect 22848 54738 22876 55286
rect 22928 55208 22980 55214
rect 22928 55150 22980 55156
rect 22100 54732 22152 54738
rect 22100 54674 22152 54680
rect 22836 54732 22888 54738
rect 22836 54674 22888 54680
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 22112 53718 22140 54674
rect 22940 54330 22968 55150
rect 23124 55078 23152 56646
rect 23216 56302 23244 59200
rect 24044 57594 24072 59200
rect 24032 57588 24084 57594
rect 24032 57530 24084 57536
rect 24216 57452 24268 57458
rect 24216 57394 24268 57400
rect 24124 57248 24176 57254
rect 24124 57190 24176 57196
rect 23388 56840 23440 56846
rect 23388 56782 23440 56788
rect 23400 56506 23428 56782
rect 23388 56500 23440 56506
rect 23388 56442 23440 56448
rect 24136 56302 24164 57190
rect 23204 56296 23256 56302
rect 23204 56238 23256 56244
rect 23388 56296 23440 56302
rect 23388 56238 23440 56244
rect 24124 56296 24176 56302
rect 24124 56238 24176 56244
rect 23400 55350 23428 56238
rect 24228 55826 24256 57394
rect 24308 57384 24360 57390
rect 24308 57326 24360 57332
rect 24584 57384 24636 57390
rect 24584 57326 24636 57332
rect 24320 55962 24348 57326
rect 24596 56506 24624 57326
rect 24584 56500 24636 56506
rect 24584 56442 24636 56448
rect 24308 55956 24360 55962
rect 24308 55898 24360 55904
rect 24596 55826 24624 56442
rect 24216 55820 24268 55826
rect 24216 55762 24268 55768
rect 24584 55820 24636 55826
rect 24584 55762 24636 55768
rect 23388 55344 23440 55350
rect 23388 55286 23440 55292
rect 24780 55282 24808 59200
rect 25608 57633 25636 59200
rect 26436 57798 26464 59200
rect 27172 58018 27200 59200
rect 27172 57990 27384 58018
rect 27252 57928 27304 57934
rect 27252 57870 27304 57876
rect 26424 57792 26476 57798
rect 26424 57734 26476 57740
rect 25594 57624 25650 57633
rect 25594 57559 25650 57568
rect 27068 57588 27120 57594
rect 27068 57530 27120 57536
rect 26148 57520 26200 57526
rect 26148 57462 26200 57468
rect 26700 57520 26752 57526
rect 26884 57520 26936 57526
rect 26752 57468 26832 57474
rect 26700 57462 26832 57468
rect 26884 57462 26936 57468
rect 25964 57384 26016 57390
rect 25964 57326 26016 57332
rect 25872 57248 25924 57254
rect 25872 57190 25924 57196
rect 25884 56914 25912 57190
rect 25872 56908 25924 56914
rect 25872 56850 25924 56856
rect 25596 56704 25648 56710
rect 25596 56646 25648 56652
rect 25608 56302 25636 56646
rect 25320 56296 25372 56302
rect 25320 56238 25372 56244
rect 25596 56296 25648 56302
rect 25596 56238 25648 56244
rect 25228 55820 25280 55826
rect 25228 55762 25280 55768
rect 24768 55276 24820 55282
rect 24768 55218 24820 55224
rect 23388 55208 23440 55214
rect 23388 55150 23440 55156
rect 23296 55140 23348 55146
rect 23296 55082 23348 55088
rect 23112 55072 23164 55078
rect 23112 55014 23164 55020
rect 23308 54330 23336 55082
rect 23400 54874 23428 55150
rect 23848 55140 23900 55146
rect 23848 55082 23900 55088
rect 23860 54874 23888 55082
rect 24308 55072 24360 55078
rect 24308 55014 24360 55020
rect 23388 54868 23440 54874
rect 23388 54810 23440 54816
rect 23848 54868 23900 54874
rect 23848 54810 23900 54816
rect 22928 54324 22980 54330
rect 22928 54266 22980 54272
rect 23296 54324 23348 54330
rect 23296 54266 23348 54272
rect 23400 54126 23428 54810
rect 24320 54738 24348 55014
rect 24308 54732 24360 54738
rect 24308 54674 24360 54680
rect 23940 54528 23992 54534
rect 23940 54470 23992 54476
rect 23952 54330 23980 54470
rect 23940 54324 23992 54330
rect 23940 54266 23992 54272
rect 24320 54194 24348 54674
rect 25240 54670 25268 55762
rect 25332 54738 25360 56238
rect 25884 55214 25912 56850
rect 25976 56710 26004 57326
rect 26160 57254 26188 57462
rect 26712 57446 26832 57462
rect 26332 57384 26384 57390
rect 26332 57326 26384 57332
rect 26148 57248 26200 57254
rect 26148 57190 26200 57196
rect 26344 56846 26372 57326
rect 26700 57316 26752 57322
rect 26700 57258 26752 57264
rect 26712 56914 26740 57258
rect 26700 56908 26752 56914
rect 26700 56850 26752 56856
rect 26332 56840 26384 56846
rect 26332 56782 26384 56788
rect 25964 56704 26016 56710
rect 25964 56646 26016 56652
rect 25976 55962 26004 56646
rect 26344 56506 26372 56782
rect 26804 56506 26832 57446
rect 26896 57050 26924 57462
rect 26884 57044 26936 57050
rect 26884 56986 26936 56992
rect 27080 56710 27108 57530
rect 27264 56914 27292 57870
rect 27252 56908 27304 56914
rect 27252 56850 27304 56856
rect 27068 56704 27120 56710
rect 27068 56646 27120 56652
rect 26332 56500 26384 56506
rect 26332 56442 26384 56448
rect 26792 56500 26844 56506
rect 26792 56442 26844 56448
rect 27356 56166 27384 57990
rect 28000 57866 28028 59200
rect 27988 57860 28040 57866
rect 27988 57802 28040 57808
rect 28356 57452 28408 57458
rect 28356 57394 28408 57400
rect 28264 57248 28316 57254
rect 28264 57190 28316 57196
rect 28276 56982 28304 57190
rect 28368 57089 28396 57394
rect 28354 57080 28410 57089
rect 28354 57015 28410 57024
rect 28264 56976 28316 56982
rect 28264 56918 28316 56924
rect 27988 56908 28040 56914
rect 27988 56850 28040 56856
rect 27896 56228 27948 56234
rect 27896 56170 27948 56176
rect 27344 56160 27396 56166
rect 27344 56102 27396 56108
rect 27908 55962 27936 56170
rect 25964 55956 26016 55962
rect 25964 55898 26016 55904
rect 27896 55956 27948 55962
rect 27896 55898 27948 55904
rect 28000 55826 28028 56850
rect 27896 55820 27948 55826
rect 27896 55762 27948 55768
rect 27988 55820 28040 55826
rect 27988 55762 28040 55768
rect 28264 55820 28316 55826
rect 28264 55762 28316 55768
rect 27436 55752 27488 55758
rect 27436 55694 27488 55700
rect 26516 55616 26568 55622
rect 26516 55558 26568 55564
rect 26884 55616 26936 55622
rect 26884 55558 26936 55564
rect 25872 55208 25924 55214
rect 25872 55150 25924 55156
rect 26528 54806 26556 55558
rect 26896 55214 26924 55558
rect 26884 55208 26936 55214
rect 26884 55150 26936 55156
rect 27448 55078 27476 55694
rect 27908 55146 27936 55762
rect 28276 55622 28304 55762
rect 28736 55622 28764 59200
rect 29274 57624 29330 57633
rect 29274 57559 29330 57568
rect 29288 57390 29316 57559
rect 29276 57384 29328 57390
rect 29276 57326 29328 57332
rect 29000 57316 29052 57322
rect 29184 57316 29236 57322
rect 29052 57276 29184 57304
rect 29000 57258 29052 57264
rect 29184 57258 29236 57264
rect 29274 57080 29330 57089
rect 29274 57015 29330 57024
rect 29184 56976 29236 56982
rect 29184 56918 29236 56924
rect 29196 56846 29224 56918
rect 29288 56846 29316 57015
rect 29564 56953 29592 59200
rect 30392 57866 30420 59200
rect 29828 57860 29880 57866
rect 29828 57802 29880 57808
rect 30380 57860 30432 57866
rect 30380 57802 30432 57808
rect 29840 57458 29868 57802
rect 29920 57588 29972 57594
rect 29920 57530 29972 57536
rect 29644 57452 29696 57458
rect 29644 57394 29696 57400
rect 29828 57452 29880 57458
rect 29828 57394 29880 57400
rect 29550 56944 29606 56953
rect 29550 56879 29606 56888
rect 29184 56840 29236 56846
rect 29090 56808 29146 56817
rect 29184 56782 29236 56788
rect 29276 56840 29328 56846
rect 29656 56817 29684 57394
rect 29932 56914 29960 57530
rect 31128 57089 31156 59200
rect 31668 57248 31720 57254
rect 31668 57190 31720 57196
rect 31114 57080 31170 57089
rect 31114 57015 31170 57024
rect 29920 56908 29972 56914
rect 29920 56850 29972 56856
rect 31300 56908 31352 56914
rect 31300 56850 31352 56856
rect 30748 56840 30800 56846
rect 29276 56782 29328 56788
rect 29642 56808 29698 56817
rect 29090 56743 29092 56752
rect 29144 56743 29146 56752
rect 30748 56782 30800 56788
rect 29642 56743 29698 56752
rect 29092 56714 29144 56720
rect 28908 56704 28960 56710
rect 29276 56704 29328 56710
rect 28960 56652 29276 56658
rect 28908 56646 29328 56652
rect 30288 56704 30340 56710
rect 30340 56652 30420 56658
rect 30288 56646 30420 56652
rect 28920 56630 29316 56646
rect 30300 56630 30420 56646
rect 29092 56296 29144 56302
rect 29092 56238 29144 56244
rect 29000 56160 29052 56166
rect 29000 56102 29052 56108
rect 29012 55826 29040 56102
rect 29000 55820 29052 55826
rect 29000 55762 29052 55768
rect 29104 55706 29132 56238
rect 30392 55758 30420 56630
rect 30472 56228 30524 56234
rect 30472 56170 30524 56176
rect 30484 55962 30512 56170
rect 30472 55956 30524 55962
rect 30472 55898 30524 55904
rect 29012 55678 29132 55706
rect 30380 55752 30432 55758
rect 30380 55694 30432 55700
rect 28264 55616 28316 55622
rect 28264 55558 28316 55564
rect 28724 55616 28776 55622
rect 28724 55558 28776 55564
rect 27896 55140 27948 55146
rect 27896 55082 27948 55088
rect 27436 55072 27488 55078
rect 27436 55014 27488 55020
rect 27448 54874 27476 55014
rect 27436 54868 27488 54874
rect 27436 54810 27488 54816
rect 26516 54800 26568 54806
rect 26516 54742 26568 54748
rect 27908 54738 27936 55082
rect 28276 54874 28304 55558
rect 29012 55214 29040 55678
rect 29000 55208 29052 55214
rect 29000 55150 29052 55156
rect 28264 54868 28316 54874
rect 28264 54810 28316 54816
rect 25320 54732 25372 54738
rect 25320 54674 25372 54680
rect 26148 54732 26200 54738
rect 26148 54674 26200 54680
rect 27896 54732 27948 54738
rect 27896 54674 27948 54680
rect 25228 54664 25280 54670
rect 25228 54606 25280 54612
rect 25240 54330 25268 54606
rect 25228 54324 25280 54330
rect 25228 54266 25280 54272
rect 24308 54188 24360 54194
rect 24308 54130 24360 54136
rect 22192 54120 22244 54126
rect 22192 54062 22244 54068
rect 23388 54120 23440 54126
rect 23388 54062 23440 54068
rect 24768 54120 24820 54126
rect 24768 54062 24820 54068
rect 22100 53712 22152 53718
rect 22100 53654 22152 53660
rect 21732 53644 21784 53650
rect 21732 53586 21784 53592
rect 21456 53032 21508 53038
rect 21456 52974 21508 52980
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 20904 52556 20956 52562
rect 20904 52498 20956 52504
rect 20916 51950 20944 52498
rect 21468 52494 21496 52974
rect 21744 52698 21772 53586
rect 22112 53106 22140 53654
rect 22204 53174 22232 54062
rect 24780 53650 24808 54062
rect 23572 53644 23624 53650
rect 23572 53586 23624 53592
rect 24768 53644 24820 53650
rect 24768 53586 24820 53592
rect 22560 53440 22612 53446
rect 22560 53382 22612 53388
rect 23480 53440 23532 53446
rect 23480 53382 23532 53388
rect 22192 53168 22244 53174
rect 22192 53110 22244 53116
rect 22100 53100 22152 53106
rect 22100 53042 22152 53048
rect 22204 52698 22232 53110
rect 22572 53038 22600 53382
rect 22836 53100 22888 53106
rect 22836 53042 22888 53048
rect 22560 53032 22612 53038
rect 22560 52974 22612 52980
rect 21732 52692 21784 52698
rect 21732 52634 21784 52640
rect 22192 52692 22244 52698
rect 22192 52634 22244 52640
rect 22572 52562 22600 52974
rect 22560 52556 22612 52562
rect 22560 52498 22612 52504
rect 21456 52488 21508 52494
rect 21456 52430 21508 52436
rect 22848 52018 22876 53042
rect 23492 53038 23520 53382
rect 23480 53032 23532 53038
rect 23480 52974 23532 52980
rect 23112 52896 23164 52902
rect 23112 52838 23164 52844
rect 23124 52562 23152 52838
rect 23480 52692 23532 52698
rect 23584 52680 23612 53586
rect 23940 53576 23992 53582
rect 23940 53518 23992 53524
rect 23664 53440 23716 53446
rect 23664 53382 23716 53388
rect 23676 52698 23704 53382
rect 23952 52902 23980 53518
rect 25228 53440 25280 53446
rect 25228 53382 25280 53388
rect 25240 53038 25268 53382
rect 25228 53032 25280 53038
rect 25228 52974 25280 52980
rect 25332 52970 25360 54674
rect 25412 54120 25464 54126
rect 25412 54062 25464 54068
rect 25424 53650 25452 54062
rect 25596 53984 25648 53990
rect 25596 53926 25648 53932
rect 25608 53650 25636 53926
rect 26160 53650 26188 54674
rect 28540 54528 28592 54534
rect 28540 54470 28592 54476
rect 28908 54528 28960 54534
rect 28908 54470 28960 54476
rect 27712 54188 27764 54194
rect 27712 54130 27764 54136
rect 26424 53984 26476 53990
rect 26424 53926 26476 53932
rect 26436 53718 26464 53926
rect 27724 53786 27752 54130
rect 27896 54052 27948 54058
rect 27896 53994 27948 54000
rect 27712 53780 27764 53786
rect 27712 53722 27764 53728
rect 26424 53712 26476 53718
rect 26424 53654 26476 53660
rect 25412 53644 25464 53650
rect 25412 53586 25464 53592
rect 25596 53644 25648 53650
rect 25596 53586 25648 53592
rect 26148 53644 26200 53650
rect 26148 53586 26200 53592
rect 26332 53644 26384 53650
rect 26332 53586 26384 53592
rect 25424 52970 25452 53586
rect 25608 53020 25636 53586
rect 26056 53576 26108 53582
rect 26056 53518 26108 53524
rect 26068 53174 26096 53518
rect 26056 53168 26108 53174
rect 26056 53110 26108 53116
rect 25688 53032 25740 53038
rect 25608 52992 25688 53020
rect 25688 52974 25740 52980
rect 25320 52964 25372 52970
rect 25320 52906 25372 52912
rect 25412 52964 25464 52970
rect 25412 52906 25464 52912
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 23532 52652 23612 52680
rect 23664 52692 23716 52698
rect 23480 52634 23532 52640
rect 23664 52634 23716 52640
rect 23112 52556 23164 52562
rect 23112 52498 23164 52504
rect 23756 52556 23808 52562
rect 23756 52498 23808 52504
rect 26148 52556 26200 52562
rect 26148 52498 26200 52504
rect 21364 52012 21416 52018
rect 21364 51954 21416 51960
rect 22836 52012 22888 52018
rect 22836 51954 22888 51960
rect 20904 51944 20956 51950
rect 20904 51886 20956 51892
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 20444 51400 20496 51406
rect 20444 51342 20496 51348
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 20456 50250 20484 51342
rect 20916 51066 20944 51886
rect 21088 51808 21140 51814
rect 21088 51750 21140 51756
rect 21100 51542 21128 51750
rect 21088 51536 21140 51542
rect 21088 51478 21140 51484
rect 21376 51270 21404 51954
rect 21456 51944 21508 51950
rect 21456 51886 21508 51892
rect 21364 51264 21416 51270
rect 21364 51206 21416 51212
rect 20904 51060 20956 51066
rect 20904 51002 20956 51008
rect 21376 50862 21404 51206
rect 21468 51066 21496 51886
rect 22848 51474 22876 51954
rect 23296 51944 23348 51950
rect 23296 51886 23348 51892
rect 23664 51944 23716 51950
rect 23664 51886 23716 51892
rect 22928 51808 22980 51814
rect 22928 51750 22980 51756
rect 22940 51542 22968 51750
rect 22928 51536 22980 51542
rect 22928 51478 22980 51484
rect 23308 51474 23336 51886
rect 23676 51610 23704 51886
rect 23768 51882 23796 52498
rect 25688 52352 25740 52358
rect 25688 52294 25740 52300
rect 24032 51944 24084 51950
rect 24032 51886 24084 51892
rect 23756 51876 23808 51882
rect 23756 51818 23808 51824
rect 23768 51610 23796 51818
rect 23664 51604 23716 51610
rect 23664 51546 23716 51552
rect 23756 51604 23808 51610
rect 23756 51546 23808 51552
rect 22284 51468 22336 51474
rect 22284 51410 22336 51416
rect 22836 51468 22888 51474
rect 22836 51410 22888 51416
rect 23296 51468 23348 51474
rect 23296 51410 23348 51416
rect 21456 51060 21508 51066
rect 21456 51002 21508 51008
rect 21364 50856 21416 50862
rect 21364 50798 21416 50804
rect 21640 50856 21692 50862
rect 21640 50798 21692 50804
rect 21272 50380 21324 50386
rect 21272 50322 21324 50328
rect 21456 50380 21508 50386
rect 21456 50322 21508 50328
rect 20812 50312 20864 50318
rect 20812 50254 20864 50260
rect 19432 50244 19484 50250
rect 19432 50186 19484 50192
rect 20444 50244 20496 50250
rect 20444 50186 20496 50192
rect 19444 49842 19472 50186
rect 20168 50176 20220 50182
rect 20168 50118 20220 50124
rect 20536 50176 20588 50182
rect 20536 50118 20588 50124
rect 19432 49836 19484 49842
rect 19432 49778 19484 49784
rect 20180 49774 20208 50118
rect 20548 49774 20576 50118
rect 20824 49978 20852 50254
rect 21284 49978 21312 50322
rect 20812 49972 20864 49978
rect 20812 49914 20864 49920
rect 21272 49972 21324 49978
rect 21272 49914 21324 49920
rect 20168 49768 20220 49774
rect 20168 49710 20220 49716
rect 20536 49768 20588 49774
rect 20536 49710 20588 49716
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 20548 48890 20576 49710
rect 21468 49434 21496 50322
rect 21456 49428 21508 49434
rect 21456 49370 21508 49376
rect 21652 49298 21680 50798
rect 22296 50726 22324 51410
rect 24044 50862 24072 51886
rect 25044 51876 25096 51882
rect 25044 51818 25096 51824
rect 25056 51066 25084 51818
rect 25596 51808 25648 51814
rect 25596 51750 25648 51756
rect 25608 51074 25636 51750
rect 25700 51542 25728 52294
rect 25964 52148 26016 52154
rect 25964 52090 26016 52096
rect 25872 51808 25924 51814
rect 25872 51750 25924 51756
rect 25688 51536 25740 51542
rect 25688 51478 25740 51484
rect 25044 51060 25096 51066
rect 25044 51002 25096 51008
rect 25516 51046 25636 51074
rect 25516 50862 25544 51046
rect 25884 50930 25912 51750
rect 25976 51610 26004 52090
rect 26160 51814 26188 52498
rect 26240 52488 26292 52494
rect 26240 52430 26292 52436
rect 26148 51808 26200 51814
rect 26148 51750 26200 51756
rect 25964 51604 26016 51610
rect 25964 51546 26016 51552
rect 25872 50924 25924 50930
rect 25872 50866 25924 50872
rect 24032 50856 24084 50862
rect 24032 50798 24084 50804
rect 25504 50856 25556 50862
rect 25504 50798 25556 50804
rect 22284 50720 22336 50726
rect 22284 50662 22336 50668
rect 22652 50720 22704 50726
rect 22652 50662 22704 50668
rect 22664 50250 22692 50662
rect 24044 50522 24072 50798
rect 25884 50726 25912 50866
rect 25976 50862 26004 51546
rect 26160 51474 26188 51750
rect 26148 51468 26200 51474
rect 26148 51410 26200 51416
rect 26252 51066 26280 52430
rect 26344 52154 26372 53586
rect 27908 53038 27936 53994
rect 28552 53718 28580 54470
rect 28920 54058 28948 54470
rect 28908 54052 28960 54058
rect 28908 53994 28960 54000
rect 28540 53712 28592 53718
rect 28540 53654 28592 53660
rect 27896 53032 27948 53038
rect 27896 52974 27948 52980
rect 28920 52970 28948 53994
rect 29012 53650 29040 55150
rect 29092 55140 29144 55146
rect 29092 55082 29144 55088
rect 29104 54330 29132 55082
rect 29552 55072 29604 55078
rect 29552 55014 29604 55020
rect 29368 54664 29420 54670
rect 29368 54606 29420 54612
rect 29092 54324 29144 54330
rect 29092 54266 29144 54272
rect 29380 54126 29408 54606
rect 29564 54126 29592 55014
rect 30760 54670 30788 56782
rect 31312 56506 31340 56850
rect 31300 56500 31352 56506
rect 31300 56442 31352 56448
rect 31680 56302 31708 57190
rect 31956 56506 31984 59200
rect 32312 57792 32364 57798
rect 32312 57734 32364 57740
rect 32324 57390 32352 57734
rect 32692 57390 32720 59200
rect 33520 57798 33548 59200
rect 34256 58018 34284 59200
rect 34164 57990 34284 58018
rect 33508 57792 33560 57798
rect 33508 57734 33560 57740
rect 33416 57520 33468 57526
rect 33416 57462 33468 57468
rect 32128 57384 32180 57390
rect 32128 57326 32180 57332
rect 32312 57384 32364 57390
rect 32312 57326 32364 57332
rect 32680 57384 32732 57390
rect 32680 57326 32732 57332
rect 32140 56778 32168 57326
rect 33324 56840 33376 56846
rect 33324 56782 33376 56788
rect 32128 56772 32180 56778
rect 32128 56714 32180 56720
rect 31944 56500 31996 56506
rect 31944 56442 31996 56448
rect 32140 56386 32168 56714
rect 32956 56704 33008 56710
rect 32956 56646 33008 56652
rect 33140 56704 33192 56710
rect 33140 56646 33192 56652
rect 32968 56409 32996 56646
rect 33048 56500 33100 56506
rect 33152 56488 33180 56646
rect 33100 56460 33180 56488
rect 33232 56500 33284 56506
rect 33048 56442 33100 56448
rect 33232 56442 33284 56448
rect 32048 56358 32168 56386
rect 32954 56400 33010 56409
rect 31668 56296 31720 56302
rect 31668 56238 31720 56244
rect 32048 56234 32076 56358
rect 32954 56335 33010 56344
rect 32128 56296 32180 56302
rect 32128 56238 32180 56244
rect 32588 56296 32640 56302
rect 32588 56238 32640 56244
rect 33046 56264 33102 56273
rect 31392 56228 31444 56234
rect 31392 56170 31444 56176
rect 32036 56228 32088 56234
rect 32036 56170 32088 56176
rect 30840 56160 30892 56166
rect 30840 56102 30892 56108
rect 30852 55418 30880 56102
rect 31404 55826 31432 56170
rect 31576 56160 31628 56166
rect 31576 56102 31628 56108
rect 31588 55826 31616 56102
rect 32048 55894 32076 56170
rect 32140 55962 32168 56238
rect 32128 55956 32180 55962
rect 32128 55898 32180 55904
rect 32036 55888 32088 55894
rect 31942 55856 31998 55865
rect 31392 55820 31444 55826
rect 31392 55762 31444 55768
rect 31576 55820 31628 55826
rect 32036 55830 32088 55836
rect 31942 55791 31998 55800
rect 31576 55762 31628 55768
rect 31956 55622 31984 55791
rect 31944 55616 31996 55622
rect 31944 55558 31996 55564
rect 32220 55616 32272 55622
rect 32220 55558 32272 55564
rect 30840 55412 30892 55418
rect 30840 55354 30892 55360
rect 32036 55276 32088 55282
rect 32036 55218 32088 55224
rect 32048 54874 32076 55218
rect 32232 55214 32260 55558
rect 32220 55208 32272 55214
rect 32220 55150 32272 55156
rect 32600 55146 32628 56238
rect 33046 56199 33048 56208
rect 33100 56199 33102 56208
rect 33048 56170 33100 56176
rect 33244 55962 33272 56442
rect 33140 55956 33192 55962
rect 33140 55898 33192 55904
rect 33232 55956 33284 55962
rect 33232 55898 33284 55904
rect 32864 55276 32916 55282
rect 32864 55218 32916 55224
rect 32588 55140 32640 55146
rect 32588 55082 32640 55088
rect 32036 54868 32088 54874
rect 32036 54810 32088 54816
rect 31760 54800 31812 54806
rect 31760 54742 31812 54748
rect 30748 54664 30800 54670
rect 30748 54606 30800 54612
rect 31772 54602 31800 54742
rect 32600 54738 32628 55082
rect 32876 54738 32904 55218
rect 33152 54874 33180 55898
rect 33336 55842 33364 56782
rect 33428 56370 33456 57462
rect 33784 57384 33836 57390
rect 33784 57326 33836 57332
rect 33416 56364 33468 56370
rect 33416 56306 33468 56312
rect 33416 56228 33468 56234
rect 33416 56170 33468 56176
rect 33244 55814 33364 55842
rect 33244 55758 33272 55814
rect 33232 55752 33284 55758
rect 33232 55694 33284 55700
rect 33140 54868 33192 54874
rect 33140 54810 33192 54816
rect 32588 54732 32640 54738
rect 32588 54674 32640 54680
rect 32864 54732 32916 54738
rect 33048 54732 33100 54738
rect 32864 54674 32916 54680
rect 32968 54692 33048 54720
rect 29920 54596 29972 54602
rect 29920 54538 29972 54544
rect 31760 54596 31812 54602
rect 31760 54538 31812 54544
rect 29932 54126 29960 54538
rect 29184 54120 29236 54126
rect 29184 54062 29236 54068
rect 29368 54120 29420 54126
rect 29368 54062 29420 54068
rect 29552 54120 29604 54126
rect 29552 54062 29604 54068
rect 29920 54120 29972 54126
rect 29920 54062 29972 54068
rect 31484 54120 31536 54126
rect 31484 54062 31536 54068
rect 29000 53644 29052 53650
rect 29000 53586 29052 53592
rect 29196 53242 29224 54062
rect 29380 53786 29408 54062
rect 29368 53780 29420 53786
rect 29368 53722 29420 53728
rect 29184 53236 29236 53242
rect 29184 53178 29236 53184
rect 29380 53106 29408 53722
rect 29368 53100 29420 53106
rect 29368 53042 29420 53048
rect 29564 53038 29592 54062
rect 29932 53242 29960 54062
rect 30656 53712 30708 53718
rect 30656 53654 30708 53660
rect 31300 53712 31352 53718
rect 31300 53654 31352 53660
rect 30012 53576 30064 53582
rect 30012 53518 30064 53524
rect 29920 53236 29972 53242
rect 29920 53178 29972 53184
rect 29552 53032 29604 53038
rect 29552 52974 29604 52980
rect 28908 52964 28960 52970
rect 28908 52906 28960 52912
rect 29092 52624 29144 52630
rect 29092 52566 29144 52572
rect 26332 52148 26384 52154
rect 26332 52090 26384 52096
rect 26344 51270 26372 52090
rect 28172 51944 28224 51950
rect 28172 51886 28224 51892
rect 28632 51944 28684 51950
rect 28632 51886 28684 51892
rect 27804 51808 27856 51814
rect 27804 51750 27856 51756
rect 27816 51542 27844 51750
rect 27804 51536 27856 51542
rect 27804 51478 27856 51484
rect 26332 51264 26384 51270
rect 26332 51206 26384 51212
rect 26240 51060 26292 51066
rect 26240 51002 26292 51008
rect 25964 50856 26016 50862
rect 25964 50798 26016 50804
rect 25872 50720 25924 50726
rect 25872 50662 25924 50668
rect 24032 50516 24084 50522
rect 24032 50458 24084 50464
rect 25884 50386 25912 50662
rect 23480 50380 23532 50386
rect 23480 50322 23532 50328
rect 25504 50380 25556 50386
rect 25504 50322 25556 50328
rect 25872 50380 25924 50386
rect 25872 50322 25924 50328
rect 22652 50244 22704 50250
rect 22652 50186 22704 50192
rect 22560 50176 22612 50182
rect 22560 50118 22612 50124
rect 22376 49632 22428 49638
rect 22376 49574 22428 49580
rect 22388 49298 22416 49574
rect 22572 49298 22600 50118
rect 22664 49842 22692 50186
rect 22652 49836 22704 49842
rect 22652 49778 22704 49784
rect 21640 49292 21692 49298
rect 21640 49234 21692 49240
rect 22376 49292 22428 49298
rect 22376 49234 22428 49240
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 20444 48884 20496 48890
rect 20444 48826 20496 48832
rect 20536 48884 20588 48890
rect 20536 48826 20588 48832
rect 18144 48680 18196 48686
rect 18144 48622 18196 48628
rect 16488 48272 16540 48278
rect 16488 48214 16540 48220
rect 16120 48204 16172 48210
rect 16120 48146 16172 48152
rect 15752 48136 15804 48142
rect 15752 48078 15804 48084
rect 15016 48000 15068 48006
rect 15016 47942 15068 47948
rect 15028 47598 15056 47942
rect 13912 47592 13964 47598
rect 13912 47534 13964 47540
rect 15016 47592 15068 47598
rect 15016 47534 15068 47540
rect 13924 46442 13952 47534
rect 15764 47462 15792 48078
rect 15752 47456 15804 47462
rect 15752 47398 15804 47404
rect 15764 47258 15792 47398
rect 15752 47252 15804 47258
rect 15752 47194 15804 47200
rect 15384 47116 15436 47122
rect 15384 47058 15436 47064
rect 15292 47048 15344 47054
rect 15292 46990 15344 46996
rect 14740 46912 14792 46918
rect 14740 46854 14792 46860
rect 15108 46912 15160 46918
rect 15108 46854 15160 46860
rect 14752 46510 14780 46854
rect 15120 46714 15148 46854
rect 15108 46708 15160 46714
rect 15108 46650 15160 46656
rect 15120 46510 15148 46650
rect 14740 46504 14792 46510
rect 14740 46446 14792 46452
rect 15108 46504 15160 46510
rect 15304 46492 15332 46990
rect 15396 46714 15424 47058
rect 16132 46986 16160 48146
rect 16396 48000 16448 48006
rect 16396 47942 16448 47948
rect 16408 47122 16436 47942
rect 16500 47802 16528 48214
rect 17960 48204 18012 48210
rect 17960 48146 18012 48152
rect 17408 48000 17460 48006
rect 17408 47942 17460 47948
rect 16488 47796 16540 47802
rect 16488 47738 16540 47744
rect 16500 47190 16528 47738
rect 17420 47598 17448 47942
rect 17408 47592 17460 47598
rect 17408 47534 17460 47540
rect 16488 47184 16540 47190
rect 16488 47126 16540 47132
rect 16396 47116 16448 47122
rect 16396 47058 16448 47064
rect 17040 47116 17092 47122
rect 17040 47058 17092 47064
rect 16120 46980 16172 46986
rect 16120 46922 16172 46928
rect 16408 46714 16436 47058
rect 15384 46708 15436 46714
rect 15384 46650 15436 46656
rect 16396 46708 16448 46714
rect 16396 46650 16448 46656
rect 15384 46504 15436 46510
rect 15304 46464 15384 46492
rect 15108 46446 15160 46452
rect 15384 46446 15436 46452
rect 16764 46504 16816 46510
rect 16764 46446 16816 46452
rect 13912 46436 13964 46442
rect 13912 46378 13964 46384
rect 13924 45966 13952 46378
rect 15396 46034 15424 46446
rect 15384 46028 15436 46034
rect 15384 45970 15436 45976
rect 13912 45960 13964 45966
rect 13912 45902 13964 45908
rect 13924 45554 13952 45902
rect 14832 45824 14884 45830
rect 14832 45766 14884 45772
rect 13924 45526 14044 45554
rect 14016 45490 14044 45526
rect 14004 45484 14056 45490
rect 14004 45426 14056 45432
rect 14016 39846 14044 45426
rect 14844 45422 14872 45766
rect 15396 45626 15424 45970
rect 15384 45620 15436 45626
rect 15384 45562 15436 45568
rect 14832 45416 14884 45422
rect 14832 45358 14884 45364
rect 16776 44946 16804 46446
rect 17052 46170 17080 47058
rect 17972 47054 18000 48146
rect 18156 47530 18184 48622
rect 18420 48612 18472 48618
rect 18420 48554 18472 48560
rect 20352 48612 20404 48618
rect 20352 48554 20404 48560
rect 18432 48346 18460 48554
rect 19340 48544 19392 48550
rect 19340 48486 19392 48492
rect 18420 48340 18472 48346
rect 18420 48282 18472 48288
rect 19352 48210 19380 48486
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 19340 48204 19392 48210
rect 19340 48146 19392 48152
rect 19432 48136 19484 48142
rect 19432 48078 19484 48084
rect 18788 47660 18840 47666
rect 18788 47602 18840 47608
rect 18144 47524 18196 47530
rect 18144 47466 18196 47472
rect 18800 47122 18828 47602
rect 19156 47592 19208 47598
rect 19156 47534 19208 47540
rect 19340 47592 19392 47598
rect 19340 47534 19392 47540
rect 19168 47122 19196 47534
rect 18788 47116 18840 47122
rect 18788 47058 18840 47064
rect 19156 47116 19208 47122
rect 19156 47058 19208 47064
rect 17960 47048 18012 47054
rect 17960 46990 18012 46996
rect 17776 46912 17828 46918
rect 17776 46854 17828 46860
rect 17040 46164 17092 46170
rect 17040 46106 17092 46112
rect 17052 45966 17080 46106
rect 17788 46034 17816 46854
rect 17776 46028 17828 46034
rect 17776 45970 17828 45976
rect 17040 45960 17092 45966
rect 17040 45902 17092 45908
rect 17972 45898 18000 46990
rect 18604 46912 18656 46918
rect 18604 46854 18656 46860
rect 18616 46510 18644 46854
rect 19168 46714 19196 47058
rect 19352 47054 19380 47534
rect 19444 47530 19472 48078
rect 20364 47598 20392 48554
rect 20456 48074 20484 48826
rect 21088 48680 21140 48686
rect 21088 48622 21140 48628
rect 20536 48612 20588 48618
rect 20536 48554 20588 48560
rect 20444 48068 20496 48074
rect 20444 48010 20496 48016
rect 20456 47598 20484 48010
rect 20548 48006 20576 48554
rect 20536 48000 20588 48006
rect 20536 47942 20588 47948
rect 20352 47592 20404 47598
rect 20352 47534 20404 47540
rect 20444 47592 20496 47598
rect 20444 47534 20496 47540
rect 20548 47530 20576 47942
rect 21100 47802 21128 48622
rect 21180 48544 21232 48550
rect 21180 48486 21232 48492
rect 21192 48278 21220 48486
rect 21180 48272 21232 48278
rect 21180 48214 21232 48220
rect 23492 48074 23520 50322
rect 25228 49768 25280 49774
rect 25228 49710 25280 49716
rect 24952 49632 25004 49638
rect 24952 49574 25004 49580
rect 24964 49298 24992 49574
rect 25240 49434 25268 49710
rect 25228 49428 25280 49434
rect 25228 49370 25280 49376
rect 24952 49292 25004 49298
rect 24952 49234 25004 49240
rect 25516 48890 25544 50322
rect 25780 50176 25832 50182
rect 25780 50118 25832 50124
rect 25792 49774 25820 50118
rect 26344 49774 26372 51206
rect 28184 51066 28212 51886
rect 28644 51610 28672 51886
rect 28816 51876 28868 51882
rect 28816 51818 28868 51824
rect 28632 51604 28684 51610
rect 28632 51546 28684 51552
rect 28828 51066 28856 51818
rect 29104 51610 29132 52566
rect 30024 52562 30052 53518
rect 30668 53258 30696 53654
rect 30932 53644 30984 53650
rect 30932 53586 30984 53592
rect 30668 53230 30880 53258
rect 30944 53242 30972 53586
rect 30668 53038 30696 53230
rect 30748 53100 30800 53106
rect 30748 53042 30800 53048
rect 30656 53032 30708 53038
rect 30656 52974 30708 52980
rect 30656 52896 30708 52902
rect 30656 52838 30708 52844
rect 30380 52624 30432 52630
rect 30380 52566 30432 52572
rect 30012 52556 30064 52562
rect 30012 52498 30064 52504
rect 29276 52352 29328 52358
rect 29276 52294 29328 52300
rect 29288 51882 29316 52294
rect 30024 51950 30052 52498
rect 29644 51944 29696 51950
rect 29644 51886 29696 51892
rect 30012 51944 30064 51950
rect 30012 51886 30064 51892
rect 29184 51876 29236 51882
rect 29184 51818 29236 51824
rect 29276 51876 29328 51882
rect 29276 51818 29328 51824
rect 29000 51604 29052 51610
rect 29000 51546 29052 51552
rect 29092 51604 29144 51610
rect 29092 51546 29144 51552
rect 28172 51060 28224 51066
rect 28172 51002 28224 51008
rect 28816 51060 28868 51066
rect 28816 51002 28868 51008
rect 29012 50862 29040 51546
rect 29196 51270 29224 51818
rect 29288 51490 29316 51818
rect 29552 51808 29604 51814
rect 29552 51750 29604 51756
rect 29564 51542 29592 51750
rect 29552 51536 29604 51542
rect 29288 51462 29408 51490
rect 29552 51478 29604 51484
rect 29656 51474 29684 51886
rect 29380 51406 29408 51462
rect 29644 51468 29696 51474
rect 29644 51410 29696 51416
rect 29368 51400 29420 51406
rect 29368 51342 29420 51348
rect 29184 51264 29236 51270
rect 29184 51206 29236 51212
rect 29196 51066 29224 51206
rect 29184 51060 29236 51066
rect 29184 51002 29236 51008
rect 26700 50856 26752 50862
rect 26700 50798 26752 50804
rect 28172 50856 28224 50862
rect 28172 50798 28224 50804
rect 29000 50856 29052 50862
rect 29000 50798 29052 50804
rect 26712 50386 26740 50798
rect 28184 50454 28212 50798
rect 28172 50448 28224 50454
rect 28172 50390 28224 50396
rect 30024 50386 30052 51886
rect 26700 50380 26752 50386
rect 26700 50322 26752 50328
rect 29000 50380 29052 50386
rect 29000 50322 29052 50328
rect 30012 50380 30064 50386
rect 30012 50322 30064 50328
rect 25780 49768 25832 49774
rect 25780 49710 25832 49716
rect 26332 49768 26384 49774
rect 26332 49710 26384 49716
rect 26516 49632 26568 49638
rect 26516 49574 26568 49580
rect 25688 49292 25740 49298
rect 25688 49234 25740 49240
rect 25504 48884 25556 48890
rect 25504 48826 25556 48832
rect 25700 48686 25728 49234
rect 25780 49224 25832 49230
rect 25780 49166 25832 49172
rect 25792 48686 25820 49166
rect 26528 49094 26556 49574
rect 26712 49434 26740 50322
rect 27896 50176 27948 50182
rect 27896 50118 27948 50124
rect 28356 50176 28408 50182
rect 28356 50118 28408 50124
rect 27908 49774 27936 50118
rect 27528 49768 27580 49774
rect 27528 49710 27580 49716
rect 27896 49768 27948 49774
rect 27896 49710 27948 49716
rect 26700 49428 26752 49434
rect 26700 49370 26752 49376
rect 27436 49224 27488 49230
rect 27436 49166 27488 49172
rect 26516 49088 26568 49094
rect 26516 49030 26568 49036
rect 24860 48680 24912 48686
rect 24860 48622 24912 48628
rect 25688 48680 25740 48686
rect 25688 48622 25740 48628
rect 25780 48680 25832 48686
rect 25780 48622 25832 48628
rect 24216 48204 24268 48210
rect 24216 48146 24268 48152
rect 23480 48068 23532 48074
rect 23480 48010 23532 48016
rect 21088 47796 21140 47802
rect 21088 47738 21140 47744
rect 19432 47524 19484 47530
rect 19432 47466 19484 47472
rect 20536 47524 20588 47530
rect 20536 47466 20588 47472
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19156 46708 19208 46714
rect 19156 46650 19208 46656
rect 19444 46578 19472 47466
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 23492 47122 23520 48010
rect 23572 47592 23624 47598
rect 23572 47534 23624 47540
rect 20168 47116 20220 47122
rect 20168 47058 20220 47064
rect 21456 47116 21508 47122
rect 21456 47058 21508 47064
rect 23480 47116 23532 47122
rect 23480 47058 23532 47064
rect 20076 46912 20128 46918
rect 20076 46854 20128 46860
rect 19432 46572 19484 46578
rect 19432 46514 19484 46520
rect 18604 46504 18656 46510
rect 18604 46446 18656 46452
rect 19444 46170 19472 46514
rect 20088 46510 20116 46854
rect 20180 46714 20208 47058
rect 20628 47048 20680 47054
rect 20628 46990 20680 46996
rect 20168 46708 20220 46714
rect 20168 46650 20220 46656
rect 20076 46504 20128 46510
rect 20076 46446 20128 46452
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19580 46192 19876 46212
rect 20640 46170 20668 46990
rect 20904 46504 20956 46510
rect 20904 46446 20956 46452
rect 19432 46164 19484 46170
rect 19432 46106 19484 46112
rect 20628 46164 20680 46170
rect 20628 46106 20680 46112
rect 17960 45892 18012 45898
rect 17960 45834 18012 45840
rect 18604 45824 18656 45830
rect 18604 45766 18656 45772
rect 18616 45558 18644 45766
rect 17960 45552 18012 45558
rect 17960 45494 18012 45500
rect 18604 45552 18656 45558
rect 18604 45494 18656 45500
rect 17592 45416 17644 45422
rect 17592 45358 17644 45364
rect 17408 45280 17460 45286
rect 17408 45222 17460 45228
rect 17420 45014 17448 45222
rect 17408 45008 17460 45014
rect 17408 44950 17460 44956
rect 16764 44940 16816 44946
rect 16764 44882 16816 44888
rect 15200 40588 15252 40594
rect 15200 40530 15252 40536
rect 15292 40588 15344 40594
rect 15292 40530 15344 40536
rect 13728 39840 13780 39846
rect 13728 39782 13780 39788
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 13740 39438 13768 39782
rect 13728 39432 13780 39438
rect 13728 39374 13780 39380
rect 13740 38418 13768 39374
rect 15212 39098 15240 40530
rect 15200 39092 15252 39098
rect 15200 39034 15252 39040
rect 15304 39030 15332 40530
rect 15384 40384 15436 40390
rect 15384 40326 15436 40332
rect 15396 39574 15424 40326
rect 15752 40112 15804 40118
rect 15752 40054 15804 40060
rect 15476 39840 15528 39846
rect 15476 39782 15528 39788
rect 15384 39568 15436 39574
rect 15384 39510 15436 39516
rect 15292 39024 15344 39030
rect 15292 38966 15344 38972
rect 13728 38412 13780 38418
rect 13728 38354 13780 38360
rect 13740 37806 13768 38354
rect 15108 38344 15160 38350
rect 15108 38286 15160 38292
rect 14740 38208 14792 38214
rect 14740 38150 14792 38156
rect 14752 37806 14780 38150
rect 15120 38010 15148 38286
rect 15304 38214 15332 38966
rect 15488 38758 15516 39782
rect 15568 39296 15620 39302
rect 15568 39238 15620 39244
rect 15580 38894 15608 39238
rect 15764 38894 15792 40054
rect 16776 39982 16804 44882
rect 17604 44538 17632 45358
rect 17592 44532 17644 44538
rect 17592 44474 17644 44480
rect 17972 44266 18000 45494
rect 19444 45422 19472 46106
rect 19892 46028 19944 46034
rect 19892 45970 19944 45976
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 18144 45416 18196 45422
rect 18144 45358 18196 45364
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 18156 45082 18184 45358
rect 18696 45348 18748 45354
rect 18696 45290 18748 45296
rect 18708 45082 18736 45290
rect 18144 45076 18196 45082
rect 18144 45018 18196 45024
rect 18696 45076 18748 45082
rect 18696 45018 18748 45024
rect 18156 44334 18184 45018
rect 19444 44878 19472 45358
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 19904 44810 19932 45970
rect 20076 45824 20128 45830
rect 20076 45766 20128 45772
rect 19984 45280 20036 45286
rect 19984 45222 20036 45228
rect 19996 44946 20024 45222
rect 20088 45014 20116 45766
rect 20180 45286 20208 45970
rect 20916 45422 20944 46446
rect 21468 46170 21496 47058
rect 22744 46980 22796 46986
rect 22744 46922 22796 46928
rect 23480 46980 23532 46986
rect 23584 46968 23612 47534
rect 24228 47258 24256 48146
rect 24872 48006 24900 48622
rect 26528 48618 26556 49030
rect 26700 48680 26752 48686
rect 26700 48622 26752 48628
rect 26516 48612 26568 48618
rect 26516 48554 26568 48560
rect 26608 48544 26660 48550
rect 26608 48486 26660 48492
rect 25320 48204 25372 48210
rect 25320 48146 25372 48152
rect 26332 48204 26384 48210
rect 26332 48146 26384 48152
rect 25136 48136 25188 48142
rect 25136 48078 25188 48084
rect 24860 48000 24912 48006
rect 24860 47942 24912 47948
rect 24216 47252 24268 47258
rect 24216 47194 24268 47200
rect 23532 46940 23612 46968
rect 24768 46980 24820 46986
rect 23480 46922 23532 46928
rect 24768 46922 24820 46928
rect 22560 46912 22612 46918
rect 22560 46854 22612 46860
rect 22468 46708 22520 46714
rect 22468 46650 22520 46656
rect 22100 46368 22152 46374
rect 22100 46310 22152 46316
rect 22112 46170 22140 46310
rect 21456 46164 21508 46170
rect 21456 46106 21508 46112
rect 22100 46164 22152 46170
rect 22100 46106 22152 46112
rect 22112 45898 22140 46106
rect 22100 45892 22152 45898
rect 22100 45834 22152 45840
rect 22480 45830 22508 46650
rect 22572 46442 22600 46854
rect 22560 46436 22612 46442
rect 22560 46378 22612 46384
rect 22572 46050 22600 46378
rect 22756 46102 22784 46922
rect 23388 46504 23440 46510
rect 23388 46446 23440 46452
rect 22836 46436 22888 46442
rect 22836 46378 22888 46384
rect 22744 46096 22796 46102
rect 22572 46034 22692 46050
rect 22744 46038 22796 46044
rect 22560 46028 22692 46034
rect 22612 46022 22692 46028
rect 22560 45970 22612 45976
rect 22572 45939 22600 45970
rect 22560 45892 22612 45898
rect 22560 45834 22612 45840
rect 22468 45824 22520 45830
rect 22468 45766 22520 45772
rect 22480 45422 22508 45766
rect 20904 45416 20956 45422
rect 20904 45358 20956 45364
rect 20996 45416 21048 45422
rect 20996 45358 21048 45364
rect 21640 45416 21692 45422
rect 21640 45358 21692 45364
rect 22468 45416 22520 45422
rect 22468 45358 22520 45364
rect 20168 45280 20220 45286
rect 20168 45222 20220 45228
rect 20720 45280 20772 45286
rect 20720 45222 20772 45228
rect 20732 45014 20760 45222
rect 20076 45008 20128 45014
rect 20076 44950 20128 44956
rect 20352 45008 20404 45014
rect 20352 44950 20404 44956
rect 20720 45008 20772 45014
rect 20720 44950 20772 44956
rect 19984 44940 20036 44946
rect 19984 44882 20036 44888
rect 19340 44804 19392 44810
rect 19340 44746 19392 44752
rect 19892 44804 19944 44810
rect 19892 44746 19944 44752
rect 19352 44538 19380 44746
rect 19340 44532 19392 44538
rect 19340 44474 19392 44480
rect 20364 44334 20392 44950
rect 20916 44538 20944 45358
rect 20904 44532 20956 44538
rect 20904 44474 20956 44480
rect 21008 44334 21036 45358
rect 21652 45082 21680 45358
rect 21640 45076 21692 45082
rect 21640 45018 21692 45024
rect 21652 44334 21680 45018
rect 22572 44334 22600 45834
rect 22664 45354 22692 46022
rect 22848 45422 22876 46378
rect 22928 46368 22980 46374
rect 22928 46310 22980 46316
rect 23020 46368 23072 46374
rect 23020 46310 23072 46316
rect 22940 45422 22968 46310
rect 23032 46102 23060 46310
rect 23020 46096 23072 46102
rect 23020 46038 23072 46044
rect 23400 45626 23428 46446
rect 23492 46034 23520 46922
rect 24676 46572 24728 46578
rect 24676 46514 24728 46520
rect 24584 46368 24636 46374
rect 24584 46310 24636 46316
rect 24596 46102 24624 46310
rect 24584 46096 24636 46102
rect 24584 46038 24636 46044
rect 23480 46028 23532 46034
rect 23480 45970 23532 45976
rect 24688 45966 24716 46514
rect 24780 46510 24808 46922
rect 24768 46504 24820 46510
rect 24768 46446 24820 46452
rect 24952 46504 25004 46510
rect 24952 46446 25004 46452
rect 25044 46504 25096 46510
rect 25044 46446 25096 46452
rect 24676 45960 24728 45966
rect 24676 45902 24728 45908
rect 23388 45620 23440 45626
rect 23388 45562 23440 45568
rect 24308 45484 24360 45490
rect 24308 45426 24360 45432
rect 22836 45416 22888 45422
rect 22836 45358 22888 45364
rect 22928 45416 22980 45422
rect 22928 45358 22980 45364
rect 23940 45416 23992 45422
rect 23940 45358 23992 45364
rect 24216 45416 24268 45422
rect 24216 45358 24268 45364
rect 22652 45348 22704 45354
rect 22652 45290 22704 45296
rect 22940 44878 22968 45358
rect 23388 45280 23440 45286
rect 23388 45222 23440 45228
rect 23400 44946 23428 45222
rect 23388 44940 23440 44946
rect 23388 44882 23440 44888
rect 22928 44872 22980 44878
rect 22928 44814 22980 44820
rect 22652 44736 22704 44742
rect 22652 44678 22704 44684
rect 22664 44334 22692 44678
rect 18144 44328 18196 44334
rect 18144 44270 18196 44276
rect 20352 44328 20404 44334
rect 20352 44270 20404 44276
rect 20996 44328 21048 44334
rect 20996 44270 21048 44276
rect 21640 44328 21692 44334
rect 21640 44270 21692 44276
rect 22560 44328 22612 44334
rect 22560 44270 22612 44276
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 17960 44260 18012 44266
rect 17960 44202 18012 44208
rect 22572 44180 22600 44270
rect 22572 44152 22692 44180
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 21088 43920 21140 43926
rect 21088 43862 21140 43868
rect 21180 43920 21232 43926
rect 21180 43862 21232 43868
rect 20904 43784 20956 43790
rect 20904 43726 20956 43732
rect 20444 43648 20496 43654
rect 20444 43590 20496 43596
rect 20456 43246 20484 43590
rect 20168 43240 20220 43246
rect 20168 43182 20220 43188
rect 20444 43240 20496 43246
rect 20444 43182 20496 43188
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 20180 42090 20208 43182
rect 20260 42560 20312 42566
rect 20260 42502 20312 42508
rect 20272 42158 20300 42502
rect 20916 42362 20944 43726
rect 21100 42770 21128 43862
rect 21192 42906 21220 43862
rect 21364 43648 21416 43654
rect 21364 43590 21416 43596
rect 21376 43110 21404 43590
rect 22664 43178 22692 44152
rect 23400 43858 23428 44882
rect 23952 44878 23980 45358
rect 23940 44872 23992 44878
rect 23940 44814 23992 44820
rect 23848 44736 23900 44742
rect 23848 44678 23900 44684
rect 23860 44402 23888 44678
rect 23952 44538 23980 44814
rect 24228 44742 24256 45358
rect 24320 44878 24348 45426
rect 24492 45280 24544 45286
rect 24492 45222 24544 45228
rect 24504 44946 24532 45222
rect 24688 44946 24716 45902
rect 24780 45830 24808 46446
rect 24964 46034 24992 46446
rect 25056 46170 25084 46446
rect 25044 46164 25096 46170
rect 25044 46106 25096 46112
rect 24952 46028 25004 46034
rect 24952 45970 25004 45976
rect 24768 45824 24820 45830
rect 24768 45766 24820 45772
rect 24964 45626 24992 45970
rect 24952 45620 25004 45626
rect 24952 45562 25004 45568
rect 25148 45082 25176 48078
rect 25332 47802 25360 48146
rect 25412 48000 25464 48006
rect 25412 47942 25464 47948
rect 25320 47796 25372 47802
rect 25320 47738 25372 47744
rect 25228 47524 25280 47530
rect 25228 47466 25280 47472
rect 25240 47258 25268 47466
rect 25228 47252 25280 47258
rect 25228 47194 25280 47200
rect 25332 47190 25360 47738
rect 25320 47184 25372 47190
rect 25320 47126 25372 47132
rect 25424 47122 25452 47942
rect 26344 47802 26372 48146
rect 26332 47796 26384 47802
rect 26332 47738 26384 47744
rect 26620 47598 26648 48486
rect 26712 47802 26740 48622
rect 26700 47796 26752 47802
rect 26700 47738 26752 47744
rect 26608 47592 26660 47598
rect 26608 47534 26660 47540
rect 26712 47122 26740 47738
rect 25412 47116 25464 47122
rect 25412 47058 25464 47064
rect 26700 47116 26752 47122
rect 26700 47058 26752 47064
rect 26608 46912 26660 46918
rect 26608 46854 26660 46860
rect 26620 46510 26648 46854
rect 26608 46504 26660 46510
rect 26608 46446 26660 46452
rect 27448 46034 27476 49166
rect 27540 48754 27568 49710
rect 28368 49434 28396 50118
rect 29012 49978 29040 50322
rect 29000 49972 29052 49978
rect 29000 49914 29052 49920
rect 28356 49428 28408 49434
rect 28356 49370 28408 49376
rect 27528 48748 27580 48754
rect 27528 48690 27580 48696
rect 27540 48278 27568 48690
rect 27804 48680 27856 48686
rect 27804 48622 27856 48628
rect 27712 48544 27764 48550
rect 27712 48486 27764 48492
rect 27528 48272 27580 48278
rect 27528 48214 27580 48220
rect 27724 48142 27752 48486
rect 27712 48136 27764 48142
rect 27712 48078 27764 48084
rect 27724 47598 27752 48078
rect 27816 48074 27844 48622
rect 27804 48068 27856 48074
rect 27804 48010 27856 48016
rect 27816 47734 27844 48010
rect 28080 48000 28132 48006
rect 28080 47942 28132 47948
rect 28264 48000 28316 48006
rect 28264 47942 28316 47948
rect 28092 47802 28120 47942
rect 28080 47796 28132 47802
rect 28080 47738 28132 47744
rect 27804 47728 27856 47734
rect 27804 47670 27856 47676
rect 27712 47592 27764 47598
rect 27712 47534 27764 47540
rect 27896 47592 27948 47598
rect 27896 47534 27948 47540
rect 27908 47122 27936 47534
rect 27988 47524 28040 47530
rect 27988 47466 28040 47472
rect 27896 47116 27948 47122
rect 27896 47058 27948 47064
rect 27620 47048 27672 47054
rect 27620 46990 27672 46996
rect 27632 46374 27660 46990
rect 27804 46980 27856 46986
rect 27804 46922 27856 46928
rect 27816 46714 27844 46922
rect 27804 46708 27856 46714
rect 27724 46668 27804 46696
rect 27620 46368 27672 46374
rect 27620 46310 27672 46316
rect 27436 46028 27488 46034
rect 27436 45970 27488 45976
rect 26240 45416 26292 45422
rect 26240 45358 26292 45364
rect 25136 45076 25188 45082
rect 25136 45018 25188 45024
rect 24492 44940 24544 44946
rect 24492 44882 24544 44888
rect 24676 44940 24728 44946
rect 24676 44882 24728 44888
rect 24308 44872 24360 44878
rect 24308 44814 24360 44820
rect 24216 44736 24268 44742
rect 24216 44678 24268 44684
rect 23940 44532 23992 44538
rect 23940 44474 23992 44480
rect 23848 44396 23900 44402
rect 23848 44338 23900 44344
rect 24228 43994 24256 44678
rect 24320 44538 24348 44814
rect 24308 44532 24360 44538
rect 24308 44474 24360 44480
rect 25148 43994 25176 45018
rect 25228 44260 25280 44266
rect 25228 44202 25280 44208
rect 24216 43988 24268 43994
rect 24216 43930 24268 43936
rect 25136 43988 25188 43994
rect 25136 43930 25188 43936
rect 23388 43852 23440 43858
rect 23388 43794 23440 43800
rect 22744 43716 22796 43722
rect 22744 43658 22796 43664
rect 22756 43382 22784 43658
rect 22744 43376 22796 43382
rect 22744 43318 22796 43324
rect 23664 43376 23716 43382
rect 23664 43318 23716 43324
rect 22652 43172 22704 43178
rect 22652 43114 22704 43120
rect 21364 43104 21416 43110
rect 21364 43046 21416 43052
rect 22560 43104 22612 43110
rect 22560 43046 22612 43052
rect 21180 42900 21232 42906
rect 21180 42842 21232 42848
rect 21088 42764 21140 42770
rect 21088 42706 21140 42712
rect 20904 42356 20956 42362
rect 20904 42298 20956 42304
rect 20260 42152 20312 42158
rect 20260 42094 20312 42100
rect 20168 42084 20220 42090
rect 20168 42026 20220 42032
rect 20720 42084 20772 42090
rect 20720 42026 20772 42032
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 20732 41614 20760 42026
rect 21100 42022 21128 42706
rect 21192 42702 21220 42842
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 21192 42226 21220 42638
rect 21180 42220 21232 42226
rect 21180 42162 21232 42168
rect 21088 42016 21140 42022
rect 21088 41958 21140 41964
rect 21192 41818 21220 42162
rect 21376 42158 21404 43046
rect 22572 42838 22600 43046
rect 22560 42832 22612 42838
rect 22560 42774 22612 42780
rect 22664 42770 22692 43114
rect 22756 43110 22784 43318
rect 23388 43240 23440 43246
rect 23388 43182 23440 43188
rect 22744 43104 22796 43110
rect 22744 43046 22796 43052
rect 23400 42838 23428 43182
rect 23676 42906 23704 43318
rect 24308 43172 24360 43178
rect 24308 43114 24360 43120
rect 23664 42900 23716 42906
rect 23664 42842 23716 42848
rect 23848 42900 23900 42906
rect 23848 42842 23900 42848
rect 23388 42832 23440 42838
rect 23388 42774 23440 42780
rect 22652 42764 22704 42770
rect 22652 42706 22704 42712
rect 21364 42152 21416 42158
rect 21364 42094 21416 42100
rect 21180 41812 21232 41818
rect 21180 41754 21232 41760
rect 20812 41676 20864 41682
rect 20812 41618 20864 41624
rect 21180 41676 21232 41682
rect 21180 41618 21232 41624
rect 20720 41608 20772 41614
rect 20720 41550 20772 41556
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 20076 40656 20128 40662
rect 20076 40598 20128 40604
rect 19984 40588 20036 40594
rect 19984 40530 20036 40536
rect 19708 40520 19760 40526
rect 19708 40462 19760 40468
rect 18604 40384 18656 40390
rect 18604 40326 18656 40332
rect 18616 39982 18644 40326
rect 19720 40186 19748 40462
rect 19708 40180 19760 40186
rect 19708 40122 19760 40128
rect 16764 39976 16816 39982
rect 16764 39918 16816 39924
rect 17684 39976 17736 39982
rect 17684 39918 17736 39924
rect 18604 39976 18656 39982
rect 18604 39918 18656 39924
rect 16776 39642 16804 39918
rect 16764 39636 16816 39642
rect 16764 39578 16816 39584
rect 15568 38888 15620 38894
rect 15568 38830 15620 38836
rect 15752 38888 15804 38894
rect 15752 38830 15804 38836
rect 15476 38752 15528 38758
rect 15476 38694 15528 38700
rect 16776 38486 16804 39578
rect 17696 38962 17724 39918
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 18052 39500 18104 39506
rect 18052 39442 18104 39448
rect 17684 38956 17736 38962
rect 17684 38898 17736 38904
rect 17696 38842 17724 38898
rect 17604 38814 17724 38842
rect 16764 38480 16816 38486
rect 16764 38422 16816 38428
rect 15660 38412 15712 38418
rect 15660 38354 15712 38360
rect 17316 38412 17368 38418
rect 17316 38354 17368 38360
rect 15292 38208 15344 38214
rect 15292 38150 15344 38156
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 15304 37806 15332 38150
rect 15672 38010 15700 38354
rect 17328 38010 17356 38354
rect 15660 38004 15712 38010
rect 15660 37946 15712 37952
rect 17316 38004 17368 38010
rect 17316 37946 17368 37952
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 14740 37800 14792 37806
rect 14740 37742 14792 37748
rect 15292 37800 15344 37806
rect 15292 37742 15344 37748
rect 13740 36718 13768 37742
rect 15672 37330 15700 37946
rect 16396 37800 16448 37806
rect 16396 37742 16448 37748
rect 16212 37664 16264 37670
rect 16212 37606 16264 37612
rect 15752 37392 15804 37398
rect 15752 37334 15804 37340
rect 15660 37324 15712 37330
rect 15660 37266 15712 37272
rect 15200 37256 15252 37262
rect 15200 37198 15252 37204
rect 14740 37120 14792 37126
rect 14740 37062 14792 37068
rect 14752 36718 14780 37062
rect 15212 36922 15240 37198
rect 15200 36916 15252 36922
rect 15200 36858 15252 36864
rect 15764 36718 15792 37334
rect 15844 37188 15896 37194
rect 15844 37130 15896 37136
rect 15856 36922 15884 37130
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 13728 36712 13780 36718
rect 13728 36654 13780 36660
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 15752 36712 15804 36718
rect 15752 36654 15804 36660
rect 16224 36650 16252 37606
rect 16408 37466 16436 37742
rect 16396 37460 16448 37466
rect 16396 37402 16448 37408
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 17132 37324 17184 37330
rect 17132 37266 17184 37272
rect 16212 36644 16264 36650
rect 16212 36586 16264 36592
rect 16224 36310 16252 36586
rect 16212 36304 16264 36310
rect 16212 36246 16264 36252
rect 16960 36174 16988 37266
rect 17144 36378 17172 37266
rect 17604 36786 17632 38814
rect 17960 38480 18012 38486
rect 17960 38422 18012 38428
rect 17972 37874 18000 38422
rect 17960 37868 18012 37874
rect 17960 37810 18012 37816
rect 18064 37754 18092 39442
rect 19996 39098 20024 40530
rect 20088 39506 20116 40598
rect 20444 40384 20496 40390
rect 20444 40326 20496 40332
rect 20456 39982 20484 40326
rect 20444 39976 20496 39982
rect 20444 39918 20496 39924
rect 20732 39914 20760 41550
rect 20824 41070 20852 41618
rect 21192 41274 21220 41618
rect 22376 41472 22428 41478
rect 22376 41414 22428 41420
rect 21180 41268 21232 41274
rect 21180 41210 21232 41216
rect 22388 41070 22416 41414
rect 22664 41138 22692 42706
rect 23400 42158 23428 42774
rect 23572 42560 23624 42566
rect 23572 42502 23624 42508
rect 23388 42152 23440 42158
rect 23388 42094 23440 42100
rect 23584 42090 23612 42502
rect 23860 42158 23888 42842
rect 24320 42362 24348 43114
rect 25136 43104 25188 43110
rect 25136 43046 25188 43052
rect 25148 42634 25176 43046
rect 25240 42770 25268 44202
rect 26252 43994 26280 45358
rect 26424 45348 26476 45354
rect 26424 45290 26476 45296
rect 26436 45014 26464 45290
rect 26424 45008 26476 45014
rect 26424 44950 26476 44956
rect 27632 44946 27660 46310
rect 27724 45422 27752 46668
rect 27804 46650 27856 46656
rect 27804 46028 27856 46034
rect 27804 45970 27856 45976
rect 27816 45626 27844 45970
rect 27804 45620 27856 45626
rect 27804 45562 27856 45568
rect 27712 45416 27764 45422
rect 27712 45358 27764 45364
rect 27908 45082 27936 47058
rect 28000 46986 28028 47466
rect 28276 47122 28304 47942
rect 28368 47258 28396 49370
rect 29276 49292 29328 49298
rect 29276 49234 29328 49240
rect 28448 49088 28500 49094
rect 28448 49030 28500 49036
rect 28460 48686 28488 49030
rect 28448 48680 28500 48686
rect 28448 48622 28500 48628
rect 28540 48544 28592 48550
rect 28540 48486 28592 48492
rect 28552 48278 28580 48486
rect 28540 48272 28592 48278
rect 28540 48214 28592 48220
rect 29288 48074 29316 49234
rect 29276 48068 29328 48074
rect 29276 48010 29328 48016
rect 29920 48000 29972 48006
rect 29920 47942 29972 47948
rect 29932 47802 29960 47942
rect 29920 47796 29972 47802
rect 29920 47738 29972 47744
rect 29736 47592 29788 47598
rect 29736 47534 29788 47540
rect 28448 47456 28500 47462
rect 28448 47398 28500 47404
rect 29552 47456 29604 47462
rect 29552 47398 29604 47404
rect 28356 47252 28408 47258
rect 28356 47194 28408 47200
rect 28460 47122 28488 47398
rect 28264 47116 28316 47122
rect 28264 47058 28316 47064
rect 28448 47116 28500 47122
rect 28448 47058 28500 47064
rect 27988 46980 28040 46986
rect 27988 46922 28040 46928
rect 28000 46510 28028 46922
rect 27988 46504 28040 46510
rect 27988 46446 28040 46452
rect 28000 45354 28028 46446
rect 28460 46442 28488 47058
rect 29564 46442 29592 47398
rect 29748 47258 29776 47534
rect 29736 47252 29788 47258
rect 29736 47194 29788 47200
rect 29932 47190 29960 47738
rect 30288 47592 30340 47598
rect 30288 47534 30340 47540
rect 29920 47184 29972 47190
rect 29920 47126 29972 47132
rect 30300 47122 30328 47534
rect 30288 47116 30340 47122
rect 30288 47058 30340 47064
rect 30300 46714 30328 47058
rect 30288 46708 30340 46714
rect 30288 46650 30340 46656
rect 28448 46436 28500 46442
rect 28448 46378 28500 46384
rect 29552 46436 29604 46442
rect 29552 46378 29604 46384
rect 28460 45422 28488 46378
rect 29276 46096 29328 46102
rect 29276 46038 29328 46044
rect 29092 45824 29144 45830
rect 29092 45766 29144 45772
rect 29104 45422 29132 45766
rect 29288 45490 29316 46038
rect 29276 45484 29328 45490
rect 29276 45426 29328 45432
rect 28448 45416 28500 45422
rect 28448 45358 28500 45364
rect 29092 45416 29144 45422
rect 29092 45358 29144 45364
rect 27988 45348 28040 45354
rect 27988 45290 28040 45296
rect 27896 45076 27948 45082
rect 27896 45018 27948 45024
rect 27620 44940 27672 44946
rect 27620 44882 27672 44888
rect 27252 44736 27304 44742
rect 27252 44678 27304 44684
rect 27264 44334 27292 44678
rect 28460 44538 28488 45358
rect 28908 44940 28960 44946
rect 28908 44882 28960 44888
rect 28448 44532 28500 44538
rect 28448 44474 28500 44480
rect 28264 44464 28316 44470
rect 28264 44406 28316 44412
rect 26332 44328 26384 44334
rect 26332 44270 26384 44276
rect 27252 44328 27304 44334
rect 27252 44270 27304 44276
rect 26240 43988 26292 43994
rect 26240 43930 26292 43936
rect 26344 43858 26372 44270
rect 26700 44260 26752 44266
rect 26700 44202 26752 44208
rect 28080 44260 28132 44266
rect 28080 44202 28132 44208
rect 25320 43852 25372 43858
rect 25320 43794 25372 43800
rect 26332 43852 26384 43858
rect 26332 43794 26384 43800
rect 25228 42764 25280 42770
rect 25228 42706 25280 42712
rect 25136 42628 25188 42634
rect 25136 42570 25188 42576
rect 24492 42560 24544 42566
rect 24492 42502 24544 42508
rect 24308 42356 24360 42362
rect 24308 42298 24360 42304
rect 24504 42158 24532 42502
rect 25240 42362 25268 42706
rect 24952 42356 25004 42362
rect 24952 42298 25004 42304
rect 25228 42356 25280 42362
rect 25228 42298 25280 42304
rect 23848 42152 23900 42158
rect 23848 42094 23900 42100
rect 24492 42152 24544 42158
rect 24492 42094 24544 42100
rect 24584 42152 24636 42158
rect 24584 42094 24636 42100
rect 23572 42084 23624 42090
rect 23572 42026 23624 42032
rect 24216 41744 24268 41750
rect 24216 41686 24268 41692
rect 24032 41676 24084 41682
rect 24032 41618 24084 41624
rect 23664 41472 23716 41478
rect 23664 41414 23716 41420
rect 22652 41132 22704 41138
rect 22652 41074 22704 41080
rect 23676 41070 23704 41414
rect 20812 41064 20864 41070
rect 20812 41006 20864 41012
rect 21548 41064 21600 41070
rect 21548 41006 21600 41012
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 21560 40730 21588 41006
rect 21732 40996 21784 41002
rect 21732 40938 21784 40944
rect 21744 40730 21772 40938
rect 21548 40724 21600 40730
rect 21548 40666 21600 40672
rect 21732 40724 21784 40730
rect 21732 40666 21784 40672
rect 22388 40594 22416 41006
rect 24044 40594 24072 41618
rect 24124 41608 24176 41614
rect 24124 41550 24176 41556
rect 24136 41274 24164 41550
rect 24124 41268 24176 41274
rect 24124 41210 24176 41216
rect 24136 40594 24164 41210
rect 24228 40730 24256 41686
rect 24504 41682 24532 42094
rect 24596 41750 24624 42094
rect 24584 41744 24636 41750
rect 24584 41686 24636 41692
rect 24492 41676 24544 41682
rect 24492 41618 24544 41624
rect 24964 41070 24992 42298
rect 25228 41472 25280 41478
rect 25228 41414 25280 41420
rect 25240 41070 25268 41414
rect 24952 41064 25004 41070
rect 24952 41006 25004 41012
rect 25228 41064 25280 41070
rect 25228 41006 25280 41012
rect 24216 40724 24268 40730
rect 24216 40666 24268 40672
rect 20904 40588 20956 40594
rect 20904 40530 20956 40536
rect 22376 40588 22428 40594
rect 22376 40530 22428 40536
rect 24032 40588 24084 40594
rect 24032 40530 24084 40536
rect 24124 40588 24176 40594
rect 24124 40530 24176 40536
rect 20812 40384 20864 40390
rect 20812 40326 20864 40332
rect 20720 39908 20772 39914
rect 20720 39850 20772 39856
rect 20076 39500 20128 39506
rect 20076 39442 20128 39448
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 20732 38894 20760 39850
rect 20824 39506 20852 40326
rect 20916 39642 20944 40530
rect 21088 40520 21140 40526
rect 21088 40462 21140 40468
rect 21100 40186 21128 40462
rect 21088 40180 21140 40186
rect 21088 40122 21140 40128
rect 20904 39636 20956 39642
rect 20904 39578 20956 39584
rect 21100 39506 21128 40122
rect 20812 39500 20864 39506
rect 20812 39442 20864 39448
rect 21088 39500 21140 39506
rect 21088 39442 21140 39448
rect 19892 38888 19944 38894
rect 19892 38830 19944 38836
rect 19984 38888 20036 38894
rect 19984 38830 20036 38836
rect 20444 38888 20496 38894
rect 20444 38830 20496 38836
rect 20720 38888 20772 38894
rect 20720 38830 20772 38836
rect 18972 38820 19024 38826
rect 18972 38762 19024 38768
rect 18236 38752 18288 38758
rect 18236 38694 18288 38700
rect 18248 38214 18276 38694
rect 18984 38554 19012 38762
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 18972 38548 19024 38554
rect 18972 38490 19024 38496
rect 18696 38480 18748 38486
rect 18696 38422 18748 38428
rect 18236 38208 18288 38214
rect 18236 38150 18288 38156
rect 18248 37806 18276 38150
rect 18708 37806 18736 38422
rect 19904 38418 19932 38830
rect 19996 38554 20024 38830
rect 20168 38752 20220 38758
rect 20168 38694 20220 38700
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 18880 38412 18932 38418
rect 18880 38354 18932 38360
rect 19892 38412 19944 38418
rect 19892 38354 19944 38360
rect 18892 38010 18920 38354
rect 18880 38004 18932 38010
rect 18880 37946 18932 37952
rect 17972 37726 18092 37754
rect 18236 37800 18288 37806
rect 18236 37742 18288 37748
rect 18696 37800 18748 37806
rect 18696 37742 18748 37748
rect 17972 37466 18000 37726
rect 18708 37670 18736 37742
rect 18696 37664 18748 37670
rect 18696 37606 18748 37612
rect 18708 37466 18736 37606
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 17960 37460 18012 37466
rect 17960 37402 18012 37408
rect 18696 37460 18748 37466
rect 18696 37402 18748 37408
rect 17684 37120 17736 37126
rect 17684 37062 17736 37068
rect 17592 36780 17644 36786
rect 17592 36722 17644 36728
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17696 36242 17724 37062
rect 17684 36236 17736 36242
rect 17684 36178 17736 36184
rect 16948 36168 17000 36174
rect 16948 36110 17000 36116
rect 17696 35630 17724 36178
rect 17972 35766 18000 37402
rect 18604 37392 18656 37398
rect 18604 37334 18656 37340
rect 18052 37324 18104 37330
rect 18052 37266 18104 37272
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 18064 35834 18092 37266
rect 18248 36922 18276 37266
rect 18236 36916 18288 36922
rect 18236 36858 18288 36864
rect 18420 36644 18472 36650
rect 18420 36586 18472 36592
rect 18432 36378 18460 36586
rect 18420 36372 18472 36378
rect 18420 36314 18472 36320
rect 18616 36242 18644 37334
rect 19904 37330 19932 38354
rect 19996 37346 20024 38490
rect 20180 38486 20208 38694
rect 20168 38480 20220 38486
rect 20168 38422 20220 38428
rect 20456 37466 20484 38830
rect 20732 38418 20760 38830
rect 20720 38412 20772 38418
rect 20720 38354 20772 38360
rect 20732 37466 20760 38354
rect 25332 37874 25360 43794
rect 26712 43790 26740 44202
rect 28092 43858 28120 44202
rect 28276 43858 28304 44406
rect 27896 43852 27948 43858
rect 27896 43794 27948 43800
rect 28080 43852 28132 43858
rect 28080 43794 28132 43800
rect 28264 43852 28316 43858
rect 28264 43794 28316 43800
rect 26700 43784 26752 43790
rect 26700 43726 26752 43732
rect 27528 43784 27580 43790
rect 27528 43726 27580 43732
rect 26332 43716 26384 43722
rect 26332 43658 26384 43664
rect 26344 43450 26372 43658
rect 26332 43444 26384 43450
rect 26332 43386 26384 43392
rect 26240 43240 26292 43246
rect 26240 43182 26292 43188
rect 25872 43104 25924 43110
rect 25872 43046 25924 43052
rect 25884 42838 25912 43046
rect 25872 42832 25924 42838
rect 25872 42774 25924 42780
rect 26252 42362 26280 43182
rect 26148 42356 26200 42362
rect 26148 42298 26200 42304
rect 26240 42356 26292 42362
rect 26240 42298 26292 42304
rect 25688 42016 25740 42022
rect 25688 41958 25740 41964
rect 25700 41682 25728 41958
rect 26160 41682 26188 42298
rect 26344 42158 26372 43386
rect 26712 43246 26740 43726
rect 26700 43240 26752 43246
rect 26700 43182 26752 43188
rect 27160 43240 27212 43246
rect 27160 43182 27212 43188
rect 26608 43172 26660 43178
rect 26608 43114 26660 43120
rect 26620 42906 26648 43114
rect 27172 42906 27200 43182
rect 26608 42900 26660 42906
rect 26608 42842 26660 42848
rect 27160 42900 27212 42906
rect 27160 42842 27212 42848
rect 27540 42770 27568 43726
rect 27804 43240 27856 43246
rect 27804 43182 27856 43188
rect 27528 42764 27580 42770
rect 27528 42706 27580 42712
rect 27816 42294 27844 43182
rect 27908 43110 27936 43794
rect 28092 43722 28120 43794
rect 28920 43722 28948 44882
rect 29000 44872 29052 44878
rect 29000 44814 29052 44820
rect 29012 44402 29040 44814
rect 29092 44736 29144 44742
rect 29092 44678 29144 44684
rect 29000 44396 29052 44402
rect 29000 44338 29052 44344
rect 29012 43926 29040 44338
rect 29000 43920 29052 43926
rect 29000 43862 29052 43868
rect 29104 43858 29132 44678
rect 29368 44260 29420 44266
rect 29368 44202 29420 44208
rect 29092 43852 29144 43858
rect 29092 43794 29144 43800
rect 28080 43716 28132 43722
rect 28080 43658 28132 43664
rect 28908 43716 28960 43722
rect 28908 43658 28960 43664
rect 27988 43172 28040 43178
rect 27988 43114 28040 43120
rect 27896 43104 27948 43110
rect 27896 43046 27948 43052
rect 27908 42702 27936 43046
rect 28000 42906 28028 43114
rect 27988 42900 28040 42906
rect 27988 42842 28040 42848
rect 27896 42696 27948 42702
rect 27896 42638 27948 42644
rect 27804 42288 27856 42294
rect 27804 42230 27856 42236
rect 26332 42152 26384 42158
rect 26332 42094 26384 42100
rect 27816 41818 27844 42230
rect 28092 42158 28120 43658
rect 28920 43246 28948 43658
rect 28908 43240 28960 43246
rect 28908 43182 28960 43188
rect 29104 42770 29132 43794
rect 29380 43722 29408 44202
rect 29368 43716 29420 43722
rect 29368 43658 29420 43664
rect 29736 43172 29788 43178
rect 29736 43114 29788 43120
rect 29092 42764 29144 42770
rect 29092 42706 29144 42712
rect 29552 42764 29604 42770
rect 29552 42706 29604 42712
rect 28448 42560 28500 42566
rect 28448 42502 28500 42508
rect 28460 42362 28488 42502
rect 28448 42356 28500 42362
rect 28448 42298 28500 42304
rect 28172 42288 28224 42294
rect 28172 42230 28224 42236
rect 28080 42152 28132 42158
rect 28080 42094 28132 42100
rect 27896 42084 27948 42090
rect 27896 42026 27948 42032
rect 27804 41812 27856 41818
rect 27804 41754 27856 41760
rect 27908 41682 27936 42026
rect 25504 41676 25556 41682
rect 25504 41618 25556 41624
rect 25688 41676 25740 41682
rect 25688 41618 25740 41624
rect 26148 41676 26200 41682
rect 26148 41618 26200 41624
rect 27804 41676 27856 41682
rect 27804 41618 27856 41624
rect 27896 41676 27948 41682
rect 27896 41618 27948 41624
rect 28080 41676 28132 41682
rect 28080 41618 28132 41624
rect 25412 40996 25464 41002
rect 25412 40938 25464 40944
rect 25424 40338 25452 40938
rect 25516 40458 25544 41618
rect 25700 40594 25728 41618
rect 25872 41608 25924 41614
rect 25872 41550 25924 41556
rect 25884 41274 25912 41550
rect 27816 41274 27844 41618
rect 25872 41268 25924 41274
rect 25872 41210 25924 41216
rect 27804 41268 27856 41274
rect 27804 41210 27856 41216
rect 25884 40594 25912 41210
rect 28092 41070 28120 41618
rect 28184 41546 28212 42230
rect 28448 42220 28500 42226
rect 28448 42162 28500 42168
rect 28460 41682 28488 42162
rect 28816 42152 28868 42158
rect 28816 42094 28868 42100
rect 28828 41818 28856 42094
rect 28816 41812 28868 41818
rect 28816 41754 28868 41760
rect 28448 41676 28500 41682
rect 28448 41618 28500 41624
rect 28172 41540 28224 41546
rect 28172 41482 28224 41488
rect 27620 41064 27672 41070
rect 27620 41006 27672 41012
rect 28080 41064 28132 41070
rect 28080 41006 28132 41012
rect 25688 40588 25740 40594
rect 25688 40530 25740 40536
rect 25872 40588 25924 40594
rect 25872 40530 25924 40536
rect 27632 40526 27660 41006
rect 27804 40996 27856 41002
rect 27804 40938 27856 40944
rect 27988 40996 28040 41002
rect 27988 40938 28040 40944
rect 27620 40520 27672 40526
rect 27620 40462 27672 40468
rect 27816 40458 27844 40938
rect 28000 40662 28028 40938
rect 27988 40656 28040 40662
rect 27988 40598 28040 40604
rect 27988 40520 28040 40526
rect 27988 40462 28040 40468
rect 25504 40452 25556 40458
rect 25504 40394 25556 40400
rect 27804 40452 27856 40458
rect 27804 40394 27856 40400
rect 27712 40384 27764 40390
rect 25424 40310 25544 40338
rect 27712 40326 27764 40332
rect 25516 39438 25544 40310
rect 25964 39976 26016 39982
rect 25964 39918 26016 39924
rect 25976 39642 26004 39918
rect 27724 39914 27752 40326
rect 27712 39908 27764 39914
rect 27712 39850 27764 39856
rect 26056 39840 26108 39846
rect 26056 39782 26108 39788
rect 27896 39840 27948 39846
rect 28000 39794 28028 40462
rect 27948 39788 28028 39794
rect 27896 39782 28028 39788
rect 25964 39636 26016 39642
rect 25964 39578 26016 39584
rect 25504 39432 25556 39438
rect 25504 39374 25556 39380
rect 25516 38350 25544 39374
rect 25872 39024 25924 39030
rect 25872 38966 25924 38972
rect 25884 38418 25912 38966
rect 25976 38962 26004 39578
rect 26068 39574 26096 39782
rect 27908 39766 28028 39782
rect 26056 39568 26108 39574
rect 26056 39510 26108 39516
rect 28000 39506 28028 39766
rect 28184 39642 28212 41482
rect 28460 41002 28488 41618
rect 28828 41138 28856 41754
rect 28908 41608 28960 41614
rect 28908 41550 28960 41556
rect 28816 41132 28868 41138
rect 28816 41074 28868 41080
rect 28920 41070 28948 41550
rect 28908 41064 28960 41070
rect 28908 41006 28960 41012
rect 28448 40996 28500 41002
rect 28448 40938 28500 40944
rect 28920 40594 28948 41006
rect 29564 41002 29592 42706
rect 29748 42158 29776 43114
rect 29736 42152 29788 42158
rect 29736 42094 29788 42100
rect 29828 41132 29880 41138
rect 29828 41074 29880 41080
rect 29000 40996 29052 41002
rect 29000 40938 29052 40944
rect 29552 40996 29604 41002
rect 29552 40938 29604 40944
rect 29012 40730 29040 40938
rect 29000 40724 29052 40730
rect 29000 40666 29052 40672
rect 29564 40594 29592 40938
rect 28908 40588 28960 40594
rect 28908 40530 28960 40536
rect 29276 40588 29328 40594
rect 29276 40530 29328 40536
rect 29552 40588 29604 40594
rect 29552 40530 29604 40536
rect 29288 40186 29316 40530
rect 29840 40458 29868 41074
rect 30196 40928 30248 40934
rect 30196 40870 30248 40876
rect 30208 40662 30236 40870
rect 30196 40656 30248 40662
rect 30196 40598 30248 40604
rect 29828 40452 29880 40458
rect 29828 40394 29880 40400
rect 29276 40180 29328 40186
rect 29276 40122 29328 40128
rect 29840 39982 29868 40394
rect 29828 39976 29880 39982
rect 29828 39918 29880 39924
rect 28172 39636 28224 39642
rect 28172 39578 28224 39584
rect 27344 39500 27396 39506
rect 27344 39442 27396 39448
rect 27988 39500 28040 39506
rect 27988 39442 28040 39448
rect 25964 38956 26016 38962
rect 25964 38898 26016 38904
rect 25976 38418 26004 38898
rect 27356 38894 27384 39442
rect 28540 39296 28592 39302
rect 28540 39238 28592 39244
rect 26516 38888 26568 38894
rect 26516 38830 26568 38836
rect 27344 38888 27396 38894
rect 27344 38830 27396 38836
rect 26528 38554 26556 38830
rect 26516 38548 26568 38554
rect 26516 38490 26568 38496
rect 28448 38480 28500 38486
rect 28448 38422 28500 38428
rect 25872 38412 25924 38418
rect 25872 38354 25924 38360
rect 25964 38412 26016 38418
rect 25964 38354 26016 38360
rect 27804 38412 27856 38418
rect 27804 38354 27856 38360
rect 25504 38344 25556 38350
rect 25504 38286 25556 38292
rect 27816 38010 27844 38354
rect 27804 38004 27856 38010
rect 27804 37946 27856 37952
rect 28460 37874 28488 38422
rect 28552 38350 28580 39238
rect 28816 38820 28868 38826
rect 28816 38762 28868 38768
rect 28540 38344 28592 38350
rect 28540 38286 28592 38292
rect 28552 38214 28580 38286
rect 28540 38208 28592 38214
rect 28540 38150 28592 38156
rect 28724 38208 28776 38214
rect 28724 38150 28776 38156
rect 28552 38010 28580 38150
rect 28540 38004 28592 38010
rect 28540 37946 28592 37952
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 28448 37868 28500 37874
rect 28448 37810 28500 37816
rect 21008 37670 21036 37810
rect 28552 37670 28580 37946
rect 28736 37874 28764 38150
rect 28828 38010 28856 38762
rect 29184 38752 29236 38758
rect 29184 38694 29236 38700
rect 29196 38486 29224 38694
rect 29184 38480 29236 38486
rect 29184 38422 29236 38428
rect 28908 38208 28960 38214
rect 28908 38150 28960 38156
rect 28816 38004 28868 38010
rect 28816 37946 28868 37952
rect 28724 37868 28776 37874
rect 28724 37810 28776 37816
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 28540 37664 28592 37670
rect 28540 37606 28592 37612
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 19996 37330 20116 37346
rect 19892 37324 19944 37330
rect 19996 37324 20128 37330
rect 19996 37318 20076 37324
rect 19892 37266 19944 37272
rect 20076 37266 20128 37272
rect 20720 37324 20772 37330
rect 20720 37266 20772 37272
rect 18880 36916 18932 36922
rect 18880 36858 18932 36864
rect 18892 36242 18920 36858
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 18880 36236 18932 36242
rect 18880 36178 18932 36184
rect 18788 36032 18840 36038
rect 18788 35974 18840 35980
rect 18800 35834 18828 35974
rect 18052 35828 18104 35834
rect 18052 35770 18104 35776
rect 18788 35828 18840 35834
rect 18788 35770 18840 35776
rect 17960 35760 18012 35766
rect 17960 35702 18012 35708
rect 17684 35624 17736 35630
rect 17684 35566 17736 35572
rect 18328 35624 18380 35630
rect 18328 35566 18380 35572
rect 18340 35154 18368 35566
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 18340 34746 18368 35090
rect 20732 34950 20760 37266
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 20732 34542 20760 34886
rect 17868 34536 17920 34542
rect 17868 34478 17920 34484
rect 20720 34536 20772 34542
rect 20720 34478 20772 34484
rect 13728 33040 13780 33046
rect 13728 32982 13780 32988
rect 13740 32434 13768 32982
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13636 31272 13688 31278
rect 13636 31214 13688 31220
rect 13648 30394 13676 31214
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13636 30388 13688 30394
rect 13636 30330 13688 30336
rect 13544 29504 13596 29510
rect 13596 29464 13676 29492
rect 13544 29446 13596 29452
rect 13452 28688 13504 28694
rect 13452 28630 13504 28636
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13464 26790 13492 28630
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13556 26926 13584 27270
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13452 26784 13504 26790
rect 13280 26744 13400 26772
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 12860 24692 13032 24698
rect 12808 24686 13032 24692
rect 12820 24682 13032 24686
rect 12820 24676 13044 24682
rect 12820 24670 12992 24676
rect 12992 24618 13044 24624
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12348 24142 12400 24148
rect 12438 24168 12494 24177
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11978 23760 12034 23769
rect 11978 23695 11980 23704
rect 12032 23695 12034 23704
rect 11980 23666 12032 23672
rect 12360 23662 12388 24142
rect 12438 24103 12494 24112
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12084 23254 12112 23598
rect 12072 23248 12124 23254
rect 12072 23190 12124 23196
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11440 22166 11468 22510
rect 11532 22438 11560 23122
rect 11704 23112 11756 23118
rect 11704 23054 11756 23060
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11428 22160 11480 22166
rect 11428 22102 11480 22108
rect 11532 21962 11560 22374
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 10876 21480 10928 21486
rect 10796 21440 10876 21468
rect 10796 20806 10824 21440
rect 10876 21422 10928 21428
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11152 21344 11204 21350
rect 11152 21286 11204 21292
rect 11164 21078 11192 21286
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 8852 20392 8904 20398
rect 8852 20334 8904 20340
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8864 18902 8892 20334
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9692 19378 9720 20198
rect 10704 19718 10732 20334
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8496 18154 8524 18566
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8956 3058 8984 19178
rect 9692 18834 9720 19314
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10060 18970 10088 19110
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18290 9720 18770
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 10152 18086 10180 19110
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10324 18080 10376 18086
rect 10324 18022 10376 18028
rect 10336 17202 10364 18022
rect 10520 17678 10548 19110
rect 10704 18222 10732 19654
rect 10796 19310 10824 20742
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10888 19990 10916 20198
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10980 18222 11008 20742
rect 11348 19922 11376 21422
rect 11624 21010 11652 22578
rect 11716 22506 11744 23054
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12176 22574 12204 22918
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 11704 22500 11756 22506
rect 11704 22442 11756 22448
rect 11980 22160 12032 22166
rect 11980 22102 12032 22108
rect 11992 21894 12020 22102
rect 12360 22098 12388 23122
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 11980 21888 12032 21894
rect 11980 21830 12032 21836
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11624 19310 11652 20946
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11808 19922 11836 20538
rect 12084 20398 12112 22034
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12992 21956 13044 21962
rect 12992 21898 13044 21904
rect 12452 21622 12480 21898
rect 12440 21616 12492 21622
rect 12440 21558 12492 21564
rect 12452 21486 12480 21558
rect 12256 21480 12308 21486
rect 12256 21422 12308 21428
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12268 20602 12296 21422
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 12348 20324 12400 20330
rect 12348 20266 12400 20272
rect 12360 20058 12388 20266
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12268 19922 12296 19994
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11164 18766 11192 19246
rect 12084 19242 12112 19858
rect 12452 19854 12480 21422
rect 12636 20806 12664 21422
rect 13004 21418 13032 21898
rect 13266 21856 13322 21865
rect 13266 21791 13322 21800
rect 13280 21486 13308 21791
rect 13372 21486 13400 26744
rect 13452 26726 13504 26732
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 13464 25378 13492 26318
rect 13556 26314 13584 26862
rect 13544 26308 13596 26314
rect 13544 26250 13596 26256
rect 13648 25922 13676 29464
rect 13740 28014 13768 30534
rect 13832 30394 13860 32302
rect 13912 32292 13964 32298
rect 13912 32234 13964 32240
rect 13924 30938 13952 32234
rect 14740 32224 14792 32230
rect 14740 32166 14792 32172
rect 14556 31952 14608 31958
rect 14556 31894 14608 31900
rect 14004 31748 14056 31754
rect 14004 31690 14056 31696
rect 13912 30932 13964 30938
rect 13912 30874 13964 30880
rect 13820 30388 13872 30394
rect 13820 30330 13872 30336
rect 13832 29034 13860 30330
rect 14016 29646 14044 31690
rect 14568 31142 14596 31894
rect 14556 31136 14608 31142
rect 14556 31078 14608 31084
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14384 29646 14412 30670
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14372 29640 14424 29646
rect 14372 29582 14424 29588
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13740 27674 13768 27950
rect 13912 27940 13964 27946
rect 13912 27882 13964 27888
rect 13728 27668 13780 27674
rect 13728 27610 13780 27616
rect 13728 27464 13780 27470
rect 13728 27406 13780 27412
rect 13740 26976 13768 27406
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13832 27305 13860 27338
rect 13818 27296 13874 27305
rect 13818 27231 13874 27240
rect 13820 26988 13872 26994
rect 13740 26948 13820 26976
rect 13820 26930 13872 26936
rect 13832 26382 13860 26930
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13648 25894 13768 25922
rect 13636 25764 13688 25770
rect 13636 25706 13688 25712
rect 13648 25430 13676 25706
rect 13636 25424 13688 25430
rect 13464 25350 13584 25378
rect 13636 25366 13688 25372
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13464 24954 13492 25094
rect 13452 24948 13504 24954
rect 13452 24890 13504 24896
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13464 24070 13492 24550
rect 13556 24070 13584 25350
rect 13648 24954 13676 25366
rect 13636 24948 13688 24954
rect 13636 24890 13688 24896
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13544 24064 13596 24070
rect 13544 24006 13596 24012
rect 13556 22094 13584 24006
rect 13556 22066 13676 22094
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12820 21078 12848 21286
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 13268 20596 13320 20602
rect 13372 20584 13400 21422
rect 13320 20556 13400 20584
rect 13268 20538 13320 20544
rect 13556 20466 13584 21422
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12900 19848 12952 19854
rect 13176 19848 13228 19854
rect 12952 19808 13176 19836
rect 12900 19790 12952 19796
rect 13176 19790 13228 19796
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19310 12480 19654
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9784 16658 9812 17070
rect 10428 16726 10456 17138
rect 10612 16794 10640 17750
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 11256 3670 11284 18022
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12084 16658 12112 17682
rect 12176 17610 12204 19246
rect 12992 19236 13044 19242
rect 12992 19178 13044 19184
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12254 18728 12310 18737
rect 12254 18663 12310 18672
rect 12268 18358 12296 18663
rect 12452 18578 12480 18906
rect 12544 18698 12572 18906
rect 13004 18834 13032 19178
rect 13372 18970 13400 19858
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13464 18850 13492 18906
rect 13556 18902 13584 19654
rect 12992 18828 13044 18834
rect 12992 18770 13044 18776
rect 13372 18822 13492 18850
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13648 18834 13676 22066
rect 13740 21554 13768 25894
rect 13924 22658 13952 27882
rect 14016 27878 14044 29582
rect 14384 28558 14412 29582
rect 14464 29028 14516 29034
rect 14464 28970 14516 28976
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 14016 26081 14044 27814
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14108 26858 14136 27066
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 14096 26852 14148 26858
rect 14096 26794 14148 26800
rect 14200 26761 14228 26862
rect 14186 26752 14242 26761
rect 14186 26687 14242 26696
rect 14384 26382 14412 28494
rect 14476 28014 14504 28970
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 14476 27849 14504 27950
rect 14462 27840 14518 27849
rect 14462 27775 14518 27784
rect 14568 27334 14596 31078
rect 14752 29782 14780 32166
rect 14936 31890 14964 32370
rect 15384 32360 15436 32366
rect 15384 32302 15436 32308
rect 15568 32360 15620 32366
rect 15568 32302 15620 32308
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 15016 31816 15068 31822
rect 14936 31764 15016 31770
rect 14936 31758 15068 31764
rect 14936 31726 15056 31758
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 14740 29776 14792 29782
rect 14740 29718 14792 29724
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14660 26994 14688 27474
rect 14648 26988 14700 26994
rect 14648 26930 14700 26936
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14002 26072 14058 26081
rect 14002 26007 14058 26016
rect 14280 25764 14332 25770
rect 14280 25706 14332 25712
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14016 23866 14044 24550
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14016 22982 14044 23802
rect 14200 23730 14228 24142
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14200 23610 14228 23666
rect 14292 23662 14320 25706
rect 14384 24750 14412 26318
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14476 24410 14504 24754
rect 14464 24404 14516 24410
rect 14464 24346 14516 24352
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14108 23582 14228 23610
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14476 23594 14504 24210
rect 14464 23588 14516 23594
rect 14108 23118 14136 23582
rect 14464 23530 14516 23536
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14096 23112 14148 23118
rect 14096 23054 14148 23060
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14016 22710 14044 22918
rect 13832 22630 13952 22658
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 14108 22642 14136 23054
rect 14200 22778 14228 23462
rect 14568 23254 14596 24890
rect 14660 24614 14688 25298
rect 14752 24682 14780 29446
rect 14936 28694 14964 31622
rect 14924 28688 14976 28694
rect 14924 28630 14976 28636
rect 15028 26518 15056 31726
rect 15108 31680 15160 31686
rect 15108 31622 15160 31628
rect 15120 30734 15148 31622
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 15120 29782 15148 30126
rect 15108 29776 15160 29782
rect 15108 29718 15160 29724
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15120 28422 15148 29038
rect 15108 28416 15160 28422
rect 15108 28358 15160 28364
rect 15120 28014 15148 28358
rect 15212 28014 15240 31214
rect 15396 30938 15424 32302
rect 15476 31952 15528 31958
rect 15476 31894 15528 31900
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15292 29232 15344 29238
rect 15292 29174 15344 29180
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15304 27470 15332 29174
rect 15488 28994 15516 31894
rect 15580 31890 15608 32302
rect 16028 32224 16080 32230
rect 16028 32166 16080 32172
rect 15568 31884 15620 31890
rect 15568 31826 15620 31832
rect 15580 29714 15608 31826
rect 15660 31272 15712 31278
rect 15660 31214 15712 31220
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15396 28966 15516 28994
rect 15396 27538 15424 28966
rect 15672 28150 15700 31214
rect 15844 30320 15896 30326
rect 15844 30262 15896 30268
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15764 29646 15792 29990
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15856 28801 15884 30262
rect 15936 29844 15988 29850
rect 15936 29786 15988 29792
rect 15948 29306 15976 29786
rect 15936 29300 15988 29306
rect 15936 29242 15988 29248
rect 15842 28792 15898 28801
rect 15842 28727 15898 28736
rect 15752 28484 15804 28490
rect 15752 28426 15804 28432
rect 15764 28218 15792 28426
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15660 28144 15712 28150
rect 15660 28086 15712 28092
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15488 27606 15516 27882
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15476 27600 15528 27606
rect 15476 27542 15528 27548
rect 15580 27538 15608 27814
rect 15384 27532 15436 27538
rect 15384 27474 15436 27480
rect 15568 27532 15620 27538
rect 15568 27474 15620 27480
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15016 26512 15068 26518
rect 15016 26454 15068 26460
rect 15108 25832 15160 25838
rect 15106 25800 15108 25809
rect 15160 25800 15162 25809
rect 15106 25735 15162 25744
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14740 24676 14792 24682
rect 14740 24618 14792 24624
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14844 24274 14872 25298
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 14844 23866 14872 24210
rect 14832 23860 14884 23866
rect 14832 23802 14884 23808
rect 14936 23662 14964 24210
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14096 22636 14148 22642
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13832 21486 13860 22630
rect 14096 22578 14148 22584
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 22234 13952 22510
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 14200 22030 14228 22374
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 14292 21962 14320 22374
rect 14280 21956 14332 21962
rect 14280 21898 14332 21904
rect 13820 21480 13872 21486
rect 13820 21422 13872 21428
rect 13728 21412 13780 21418
rect 13728 21354 13780 21360
rect 13740 20942 13768 21354
rect 14568 20942 14596 23190
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15028 21486 15056 22034
rect 15016 21480 15068 21486
rect 15016 21422 15068 21428
rect 14832 21004 14884 21010
rect 14832 20946 14884 20952
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14844 20602 14872 20946
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14832 20596 14884 20602
rect 14832 20538 14884 20544
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 20392 13872 20398
rect 13924 20380 13952 20470
rect 13872 20352 13952 20380
rect 13820 20334 13872 20340
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13636 18828 13688 18834
rect 13372 18698 13400 18822
rect 13636 18770 13688 18776
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 12452 18550 12572 18578
rect 12544 18426 12572 18550
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12452 18306 12480 18362
rect 12624 18352 12676 18358
rect 12452 18300 12624 18306
rect 12452 18294 12676 18300
rect 12452 18278 12664 18294
rect 12912 18222 12940 18634
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12900 18216 12952 18222
rect 12438 18184 12494 18193
rect 12900 18158 12952 18164
rect 12438 18119 12440 18128
rect 12492 18119 12494 18128
rect 12440 18090 12492 18096
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 17066 12296 17478
rect 13004 17202 13032 18566
rect 13648 18358 13676 18770
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13832 18290 13860 18566
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13832 17066 13860 17478
rect 12256 17060 12308 17066
rect 12256 17002 12308 17008
rect 13176 17060 13228 17066
rect 13176 17002 13228 17008
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 13188 4010 13216 17002
rect 13924 16794 13952 18090
rect 14016 17882 14044 19450
rect 14108 19446 14136 20538
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 19990 14228 20198
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14200 19514 14228 19722
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14096 19440 14148 19446
rect 14096 19382 14148 19388
rect 14292 19378 14320 20402
rect 15028 20398 15056 21422
rect 15120 21146 15148 25735
rect 15396 25702 15424 27474
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15488 27062 15516 27338
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15488 26450 15516 26998
rect 15856 26926 15884 28018
rect 15948 28014 15976 28086
rect 15936 28008 15988 28014
rect 15936 27950 15988 27956
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15476 26444 15528 26450
rect 15476 26386 15528 26392
rect 15488 26246 15516 26386
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15384 25696 15436 25702
rect 15580 25673 15608 25774
rect 15384 25638 15436 25644
rect 15566 25664 15622 25673
rect 15566 25599 15622 25608
rect 15660 25288 15712 25294
rect 15660 25230 15712 25236
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15212 21894 15240 23666
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15304 21962 15332 23122
rect 15396 22098 15424 23462
rect 15580 22137 15608 25162
rect 15672 24954 15700 25230
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15856 24206 15884 24686
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 22778 15700 23598
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15566 22128 15622 22137
rect 15384 22092 15436 22098
rect 15566 22063 15622 22072
rect 15384 22034 15436 22040
rect 15292 21956 15344 21962
rect 15292 21898 15344 21904
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21554 15424 21830
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15212 21146 15240 21490
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15016 20392 15068 20398
rect 15016 20334 15068 20340
rect 15028 19922 15056 20334
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14844 18902 14872 19654
rect 14936 19514 14964 19858
rect 15016 19712 15068 19718
rect 15016 19654 15068 19660
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 15028 19310 15056 19654
rect 15016 19304 15068 19310
rect 15120 19281 15148 21082
rect 15304 20466 15332 21422
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15396 19446 15424 21490
rect 15580 21486 15608 22063
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15488 21010 15516 21422
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 19786 15516 20742
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15292 19304 15344 19310
rect 15016 19246 15068 19252
rect 15106 19272 15162 19281
rect 15292 19246 15344 19252
rect 15106 19207 15162 19216
rect 14832 18896 14884 18902
rect 14832 18838 14884 18844
rect 15200 18896 15252 18902
rect 15200 18838 15252 18844
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14936 18290 14964 18566
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 14016 17338 14044 17682
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14200 17202 14228 18022
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14660 6866 14688 18090
rect 14936 17746 14964 18226
rect 15212 17882 15240 18838
rect 15304 18834 15332 19246
rect 15488 18902 15516 19722
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15580 18358 15608 20198
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15672 17814 15700 22714
rect 15844 22092 15896 22098
rect 16040 22094 16068 32166
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16304 31816 16356 31822
rect 16304 31758 16356 31764
rect 16212 27872 16264 27878
rect 16212 27814 16264 27820
rect 16224 27674 16252 27814
rect 16212 27668 16264 27674
rect 16212 27610 16264 27616
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 16132 27033 16160 27270
rect 16118 27024 16174 27033
rect 16118 26959 16174 26968
rect 16132 25158 16160 26959
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16224 26586 16252 26862
rect 16212 26580 16264 26586
rect 16212 26522 16264 26528
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 16224 25838 16252 26318
rect 16212 25832 16264 25838
rect 16212 25774 16264 25780
rect 16316 25430 16344 31758
rect 16868 31754 16896 31962
rect 17052 31890 17080 32438
rect 17880 32026 17908 34478
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 20628 34060 20680 34066
rect 20628 34002 20680 34008
rect 19892 33992 19944 33998
rect 19892 33934 19944 33940
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19904 32910 19932 33934
rect 20640 33658 20668 34002
rect 20628 33652 20680 33658
rect 20628 33594 20680 33600
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 19892 32904 19944 32910
rect 19892 32846 19944 32852
rect 18880 32360 18932 32366
rect 18880 32302 18932 32308
rect 19432 32360 19484 32366
rect 19432 32302 19484 32308
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 17972 31958 18000 32166
rect 17684 31952 17736 31958
rect 17684 31894 17736 31900
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 17040 31884 17092 31890
rect 17040 31826 17092 31832
rect 16776 31726 16896 31754
rect 16396 30932 16448 30938
rect 16396 30874 16448 30880
rect 16408 30190 16436 30874
rect 16776 30802 16804 31726
rect 17500 31204 17552 31210
rect 17500 31146 17552 31152
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 17512 30598 17540 31146
rect 17592 31136 17644 31142
rect 17592 31078 17644 31084
rect 17604 30870 17632 31078
rect 17592 30864 17644 30870
rect 17592 30806 17644 30812
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 16396 30184 16448 30190
rect 16396 30126 16448 30132
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 29714 16620 30126
rect 16684 29714 16712 30534
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 16856 29776 16908 29782
rect 16856 29718 16908 29724
rect 16396 29708 16448 29714
rect 16396 29650 16448 29656
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16672 29708 16724 29714
rect 16672 29650 16724 29656
rect 16408 27282 16436 29650
rect 16488 28960 16540 28966
rect 16488 28902 16540 28908
rect 16500 28626 16528 28902
rect 16488 28620 16540 28626
rect 16488 28562 16540 28568
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16488 27940 16540 27946
rect 16488 27882 16540 27888
rect 16500 27402 16528 27882
rect 16488 27396 16540 27402
rect 16488 27338 16540 27344
rect 16408 27254 16528 27282
rect 16500 26489 16528 27254
rect 16592 27033 16620 28358
rect 16578 27024 16634 27033
rect 16578 26959 16634 26968
rect 16486 26480 16542 26489
rect 16486 26415 16542 26424
rect 16304 25424 16356 25430
rect 16304 25366 16356 25372
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16224 25242 16252 25298
rect 16592 25242 16620 26959
rect 16670 26072 16726 26081
rect 16670 26007 16726 26016
rect 16684 25362 16712 26007
rect 16868 25362 16896 29718
rect 17144 29034 17172 30194
rect 17512 30190 17540 30534
rect 17500 30184 17552 30190
rect 17500 30126 17552 30132
rect 17696 29714 17724 31894
rect 18052 31680 18104 31686
rect 18052 31622 18104 31628
rect 18064 31278 18092 31622
rect 18892 31346 18920 32302
rect 19340 32224 19392 32230
rect 19340 32166 19392 32172
rect 19352 31482 19380 32166
rect 19444 32026 19472 32302
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 18432 30938 18460 31214
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18524 30818 18552 31282
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 18144 30796 18196 30802
rect 18144 30738 18196 30744
rect 18328 30796 18380 30802
rect 18328 30738 18380 30744
rect 18432 30790 18552 30818
rect 18604 30864 18656 30870
rect 18604 30806 18656 30812
rect 17972 30598 18000 30738
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 18156 30326 18184 30738
rect 18340 30394 18368 30738
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 30122 17908 30194
rect 17868 30116 17920 30122
rect 17868 30058 17920 30064
rect 17880 29850 17908 30058
rect 17868 29844 17920 29850
rect 17868 29786 17920 29792
rect 17224 29708 17276 29714
rect 17224 29650 17276 29656
rect 17684 29708 17736 29714
rect 17684 29650 17736 29656
rect 17236 29102 17264 29650
rect 17316 29504 17368 29510
rect 17316 29446 17368 29452
rect 18432 29458 18460 30790
rect 18512 30184 18564 30190
rect 18512 30126 18564 30132
rect 18524 29578 18552 30126
rect 18616 29714 18644 30806
rect 18892 30190 18920 31282
rect 19156 31136 19208 31142
rect 19156 31078 19208 31084
rect 18972 30252 19024 30258
rect 18972 30194 19024 30200
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 18880 30184 18932 30190
rect 18880 30126 18932 30132
rect 18708 29714 18736 30126
rect 18892 30054 18920 30126
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18696 29708 18748 29714
rect 18696 29650 18748 29656
rect 18512 29572 18564 29578
rect 18512 29514 18564 29520
rect 18604 29504 18656 29510
rect 18432 29452 18604 29458
rect 18432 29446 18656 29452
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17132 29028 17184 29034
rect 17132 28970 17184 28976
rect 17236 28626 17264 29038
rect 17224 28620 17276 28626
rect 17224 28562 17276 28568
rect 17328 28014 17356 29446
rect 18432 29430 18644 29446
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18052 29028 18104 29034
rect 18052 28970 18104 28976
rect 17866 28656 17922 28665
rect 17776 28620 17828 28626
rect 17866 28591 17922 28600
rect 17776 28562 17828 28568
rect 17684 28212 17736 28218
rect 17684 28154 17736 28160
rect 17316 28008 17368 28014
rect 17316 27950 17368 27956
rect 17592 28008 17644 28014
rect 17592 27950 17644 27956
rect 17052 27538 17264 27554
rect 17604 27538 17632 27950
rect 17040 27532 17264 27538
rect 17092 27526 17264 27532
rect 17040 27474 17092 27480
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 17052 27169 17080 27270
rect 17038 27160 17094 27169
rect 17038 27095 17094 27104
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 16946 26888 17002 26897
rect 16946 26823 17002 26832
rect 16960 26586 16988 26823
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 17052 26518 17080 26930
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16960 25702 16988 26386
rect 17144 26246 17172 27406
rect 17236 26994 17264 27526
rect 17408 27532 17460 27538
rect 17328 27492 17408 27520
rect 17328 27130 17356 27492
rect 17592 27532 17644 27538
rect 17408 27474 17460 27480
rect 17512 27492 17592 27520
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 17224 26988 17276 26994
rect 17224 26930 17276 26936
rect 17328 26314 17356 27066
rect 17512 26926 17540 27492
rect 17592 27474 17644 27480
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17604 26926 17632 27338
rect 17696 26994 17724 28154
rect 17788 27062 17816 28562
rect 17880 28558 17908 28591
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 17960 28552 18012 28558
rect 18064 28529 18092 28970
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 17960 28494 18012 28500
rect 18050 28520 18106 28529
rect 17972 28150 18000 28494
rect 18050 28455 18106 28464
rect 18236 28416 18288 28422
rect 18236 28358 18288 28364
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 18248 28014 18276 28358
rect 17960 28008 18012 28014
rect 17958 27976 17960 27985
rect 18052 28008 18104 28014
rect 18012 27976 18014 27985
rect 18052 27950 18104 27956
rect 18236 28008 18288 28014
rect 18236 27950 18288 27956
rect 17958 27911 18014 27920
rect 18064 27538 18092 27950
rect 18142 27840 18198 27849
rect 18142 27775 18198 27784
rect 18052 27532 18104 27538
rect 18052 27474 18104 27480
rect 17868 27464 17920 27470
rect 17868 27406 17920 27412
rect 17880 27130 17908 27406
rect 18156 27334 18184 27775
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18144 27328 18196 27334
rect 18144 27270 18196 27276
rect 17868 27124 17920 27130
rect 17868 27066 17920 27072
rect 17960 27124 18012 27130
rect 17960 27066 18012 27072
rect 17776 27056 17828 27062
rect 17776 26998 17828 27004
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17500 26920 17552 26926
rect 17592 26920 17644 26926
rect 17500 26862 17552 26868
rect 17590 26888 17592 26897
rect 17868 26920 17920 26926
rect 17644 26888 17646 26897
rect 17868 26862 17920 26868
rect 17590 26823 17646 26832
rect 17880 26772 17908 26862
rect 17512 26744 17908 26772
rect 17972 26761 18000 27066
rect 17958 26752 18014 26761
rect 17512 26450 17540 26744
rect 17958 26687 18014 26696
rect 17866 26480 17922 26489
rect 17500 26444 17552 26450
rect 17500 26386 17552 26392
rect 17592 26444 17644 26450
rect 17866 26415 17922 26424
rect 17592 26386 17644 26392
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 17604 26058 17632 26386
rect 17880 26382 17908 26415
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17420 26030 17632 26058
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 17316 25696 17368 25702
rect 17316 25638 17368 25644
rect 17328 25362 17356 25638
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 16224 25214 16620 25242
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 16684 24818 16712 25298
rect 16868 25242 16896 25298
rect 16776 25214 16896 25242
rect 16776 24954 16804 25214
rect 17420 25158 17448 26030
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17972 25498 18000 25774
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17500 25288 17552 25294
rect 17500 25230 17552 25236
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17512 25158 17540 25230
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16868 24750 16896 25094
rect 17420 24954 17448 25094
rect 17408 24948 17460 24954
rect 17408 24890 17460 24896
rect 17604 24886 17632 25230
rect 18064 24970 18092 27270
rect 18340 26738 18368 28562
rect 18524 27470 18552 29242
rect 18616 28626 18644 29430
rect 18708 29238 18736 29650
rect 18984 29306 19012 30194
rect 19168 29714 19196 31078
rect 19352 30122 19380 31418
rect 19444 31278 19472 31962
rect 19904 31822 19932 32846
rect 20640 32366 20668 33390
rect 20720 32564 20772 32570
rect 20720 32506 20772 32512
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20444 32224 20496 32230
rect 20444 32166 20496 32172
rect 20456 31890 20484 32166
rect 20732 31958 20760 32506
rect 21008 32502 21036 37606
rect 28080 37392 28132 37398
rect 28080 37334 28132 37340
rect 28092 36718 28120 37334
rect 28632 37324 28684 37330
rect 28632 37266 28684 37272
rect 28264 37256 28316 37262
rect 28264 37198 28316 37204
rect 28276 36922 28304 37198
rect 28264 36916 28316 36922
rect 28264 36858 28316 36864
rect 28644 36718 28672 37266
rect 28736 37262 28764 37810
rect 28920 37806 28948 38150
rect 28908 37800 28960 37806
rect 28908 37742 28960 37748
rect 28724 37256 28776 37262
rect 28724 37198 28776 37204
rect 28080 36712 28132 36718
rect 28080 36654 28132 36660
rect 28632 36712 28684 36718
rect 28632 36654 28684 36660
rect 27896 36576 27948 36582
rect 27896 36518 27948 36524
rect 27908 36310 27936 36518
rect 28644 36378 28672 36654
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 27252 36168 27304 36174
rect 27252 36110 27304 36116
rect 27264 35086 27292 36110
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27264 34746 27292 35022
rect 27252 34740 27304 34746
rect 27252 34682 27304 34688
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 25688 34060 25740 34066
rect 25688 34002 25740 34008
rect 22192 33652 22244 33658
rect 22192 33594 22244 33600
rect 22100 33448 22152 33454
rect 22100 33390 22152 33396
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 32978 21404 33254
rect 22112 33114 22140 33390
rect 22100 33108 22152 33114
rect 22100 33050 22152 33056
rect 21088 32972 21140 32978
rect 21088 32914 21140 32920
rect 21364 32972 21416 32978
rect 21364 32914 21416 32920
rect 20996 32496 21048 32502
rect 20996 32438 21048 32444
rect 20996 32360 21048 32366
rect 20996 32302 21048 32308
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 19984 31884 20036 31890
rect 19984 31826 20036 31832
rect 20444 31884 20496 31890
rect 20444 31826 20496 31832
rect 19892 31816 19944 31822
rect 19892 31758 19944 31764
rect 19996 31754 20024 31826
rect 20536 31816 20588 31822
rect 20536 31758 20588 31764
rect 19984 31748 20036 31754
rect 19984 31690 20036 31696
rect 19996 31414 20024 31690
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 20076 31272 20128 31278
rect 20076 31214 20128 31220
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19444 30666 19472 31078
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 20088 30938 20116 31214
rect 20076 30932 20128 30938
rect 19904 30892 20076 30920
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 19536 30122 19564 30262
rect 19904 30258 19932 30892
rect 20076 30874 20128 30880
rect 20548 30870 20576 31758
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20536 30864 20588 30870
rect 20536 30806 20588 30812
rect 20076 30796 20128 30802
rect 20076 30738 20128 30744
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19616 30184 19668 30190
rect 19614 30152 19616 30161
rect 19668 30152 19670 30161
rect 19340 30116 19392 30122
rect 19340 30058 19392 30064
rect 19524 30116 19576 30122
rect 19614 30087 19670 30096
rect 19524 30058 19576 30064
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19156 29708 19208 29714
rect 19156 29650 19208 29656
rect 18972 29300 19024 29306
rect 18972 29242 19024 29248
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 19168 29102 19196 29650
rect 20088 29646 20116 30738
rect 20272 30394 20300 30738
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20536 29708 20588 29714
rect 20536 29650 20588 29656
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19444 29102 19472 29514
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 19156 29096 19208 29102
rect 19432 29096 19484 29102
rect 19156 29038 19208 29044
rect 19430 29064 19432 29073
rect 19484 29064 19486 29073
rect 19430 28999 19486 29008
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 20456 28694 20484 29242
rect 20548 29170 20576 29650
rect 20536 29164 20588 29170
rect 20536 29106 20588 29112
rect 20536 29028 20588 29034
rect 20536 28970 20588 28976
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 18604 28620 18656 28626
rect 18604 28562 18656 28568
rect 18880 28620 18932 28626
rect 18880 28562 18932 28568
rect 19064 28620 19116 28626
rect 19064 28562 19116 28568
rect 19156 28620 19208 28626
rect 19156 28562 19208 28568
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18694 27976 18750 27985
rect 18616 27674 18644 27950
rect 18694 27911 18750 27920
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18616 27538 18644 27610
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18512 27464 18564 27470
rect 18512 27406 18564 27412
rect 18708 26926 18736 27911
rect 18892 27674 18920 28562
rect 19076 28218 19104 28562
rect 19064 28212 19116 28218
rect 19064 28154 19116 28160
rect 19168 27985 19196 28562
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19352 28150 19380 28494
rect 20548 28150 20576 28970
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20640 28014 20668 31078
rect 20720 30592 20772 30598
rect 20720 30534 20772 30540
rect 20732 30326 20760 30534
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20824 29084 20852 31622
rect 20916 29782 20944 32166
rect 21008 30326 21036 32302
rect 21100 32026 21128 32914
rect 21640 32768 21692 32774
rect 21640 32710 21692 32716
rect 21456 32360 21508 32366
rect 21456 32302 21508 32308
rect 21180 32224 21232 32230
rect 21180 32166 21232 32172
rect 21088 32020 21140 32026
rect 21088 31962 21140 31968
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 20996 30320 21048 30326
rect 20996 30262 21048 30268
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 20904 29232 20956 29238
rect 21008 29220 21036 30126
rect 21100 29510 21128 31826
rect 21192 31278 21220 32166
rect 21468 31278 21496 32302
rect 21652 31346 21680 32710
rect 22112 31958 22140 33050
rect 22204 32978 22232 33594
rect 22664 33454 22692 34002
rect 23112 33992 23164 33998
rect 23112 33934 23164 33940
rect 22928 33924 22980 33930
rect 22928 33866 22980 33872
rect 22652 33448 22704 33454
rect 22652 33390 22704 33396
rect 22192 32972 22244 32978
rect 22192 32914 22244 32920
rect 22100 31952 22152 31958
rect 22100 31894 22152 31900
rect 21824 31884 21876 31890
rect 21824 31826 21876 31832
rect 21836 31482 21864 31826
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 22100 31340 22152 31346
rect 22100 31282 22152 31288
rect 21180 31272 21232 31278
rect 21180 31214 21232 31220
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21652 30802 21680 31282
rect 21640 30796 21692 30802
rect 21640 30738 21692 30744
rect 22008 30320 22060 30326
rect 22008 30262 22060 30268
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 21100 29306 21128 29446
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 20956 29192 21036 29220
rect 20904 29174 20956 29180
rect 20904 29096 20956 29102
rect 20824 29056 20904 29084
rect 20904 29038 20956 29044
rect 20812 28960 20864 28966
rect 20812 28902 20864 28908
rect 20628 28008 20680 28014
rect 19154 27976 19210 27985
rect 19154 27911 19210 27920
rect 20548 27968 20628 27996
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 20168 27532 20220 27538
rect 20168 27474 20220 27480
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 18786 27160 18842 27169
rect 18786 27095 18842 27104
rect 18696 26920 18748 26926
rect 18418 26888 18474 26897
rect 18696 26862 18748 26868
rect 18418 26823 18420 26832
rect 18472 26823 18474 26832
rect 18420 26794 18472 26800
rect 18340 26710 18460 26738
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 18340 25906 18368 26318
rect 18432 25945 18460 26710
rect 18510 26072 18566 26081
rect 18510 26007 18566 26016
rect 18418 25936 18474 25945
rect 18328 25900 18380 25906
rect 18418 25871 18474 25880
rect 18328 25842 18380 25848
rect 18236 25696 18288 25702
rect 18142 25664 18198 25673
rect 18236 25638 18288 25644
rect 18142 25599 18198 25608
rect 18156 25498 18184 25599
rect 18144 25492 18196 25498
rect 18144 25434 18196 25440
rect 17880 24942 18092 24970
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 17500 24744 17552 24750
rect 17880 24698 17908 24942
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17552 24692 17908 24698
rect 17500 24686 17908 24692
rect 16764 24336 16816 24342
rect 16764 24278 16816 24284
rect 16212 23656 16264 23662
rect 16212 23598 16264 23604
rect 16396 23656 16448 23662
rect 16396 23598 16448 23604
rect 16224 23254 16252 23598
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16132 22574 16160 22918
rect 16120 22568 16172 22574
rect 16120 22510 16172 22516
rect 16408 22506 16436 23598
rect 16396 22500 16448 22506
rect 16396 22442 16448 22448
rect 16486 22128 16542 22137
rect 16040 22066 16344 22094
rect 15844 22034 15896 22040
rect 15856 21690 15884 22034
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15844 21480 15896 21486
rect 15844 21422 15896 21428
rect 15856 20262 15884 21422
rect 15948 20806 15976 21966
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21690 16160 21830
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15764 19514 15792 19858
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 16040 18222 16068 20402
rect 16132 20398 16160 20742
rect 16120 20392 16172 20398
rect 16120 20334 16172 20340
rect 16224 19922 16252 20742
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16120 19304 16172 19310
rect 16118 19272 16120 19281
rect 16172 19272 16174 19281
rect 16118 19207 16174 19216
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16132 18086 16160 19207
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15660 17808 15712 17814
rect 15660 17750 15712 17756
rect 16316 17746 16344 22066
rect 16486 22063 16542 22072
rect 16500 19310 16528 22063
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16408 18902 16436 19246
rect 16500 19174 16528 19246
rect 16672 19236 16724 19242
rect 16672 19178 16724 19184
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16684 18970 16712 19178
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16396 18896 16448 18902
rect 16396 18838 16448 18844
rect 16776 18426 16804 24278
rect 16868 18766 16896 24686
rect 17132 24676 17184 24682
rect 17512 24670 17908 24686
rect 17132 24618 17184 24624
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 17052 23186 17080 23802
rect 17040 23180 17092 23186
rect 17040 23122 17092 23128
rect 17040 22976 17092 22982
rect 17040 22918 17092 22924
rect 17052 21350 17080 22918
rect 17040 21344 17092 21350
rect 17040 21286 17092 21292
rect 17052 21010 17080 21286
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 16856 18760 16908 18766
rect 17144 18737 17172 24618
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17592 24132 17644 24138
rect 17788 24120 17816 24550
rect 17972 24274 18000 24822
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 17960 24268 18012 24274
rect 18156 24256 18184 24754
rect 18248 24596 18276 25638
rect 18432 25362 18460 25871
rect 18524 25770 18552 26007
rect 18512 25764 18564 25770
rect 18512 25706 18564 25712
rect 18604 25696 18656 25702
rect 18604 25638 18656 25644
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 18328 24880 18380 24886
rect 18524 24868 18552 25366
rect 18380 24840 18552 24868
rect 18328 24822 18380 24828
rect 18616 24750 18644 25638
rect 18708 25514 18736 26862
rect 18800 25702 18828 27095
rect 19432 26852 19484 26858
rect 19432 26794 19484 26800
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19352 26450 19380 26726
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19064 26376 19116 26382
rect 19064 26318 19116 26324
rect 19076 25974 19104 26318
rect 19064 25968 19116 25974
rect 19064 25910 19116 25916
rect 19248 25900 19300 25906
rect 19352 25888 19380 26386
rect 19444 25974 19472 26794
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19892 26444 19944 26450
rect 19892 26386 19944 26392
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 19300 25860 19380 25888
rect 19248 25842 19300 25848
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 19062 25800 19118 25809
rect 18788 25696 18840 25702
rect 18788 25638 18840 25644
rect 18708 25486 18828 25514
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18696 24676 18748 24682
rect 18696 24618 18748 24624
rect 18248 24568 18644 24596
rect 18616 24274 18644 24568
rect 18236 24268 18288 24274
rect 18156 24228 18236 24256
rect 17960 24210 18012 24216
rect 18236 24210 18288 24216
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 18052 24200 18104 24206
rect 18052 24142 18104 24148
rect 17644 24092 17816 24120
rect 17592 24074 17644 24080
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 16856 18702 16908 18708
rect 17130 18728 17186 18737
rect 17130 18663 17186 18672
rect 16764 18420 16816 18426
rect 16764 18362 16816 18368
rect 17328 18222 17356 24006
rect 17788 23186 17816 24092
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17972 24041 18000 24074
rect 17958 24032 18014 24041
rect 17958 23967 18014 23976
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17408 22568 17460 22574
rect 17408 22510 17460 22516
rect 17420 20806 17448 22510
rect 17684 22432 17736 22438
rect 17684 22374 17736 22380
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17512 20398 17540 21830
rect 17604 21146 17632 21830
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17696 21078 17724 22374
rect 17788 21486 17816 23122
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17684 21072 17736 21078
rect 17682 21040 17684 21049
rect 17736 21040 17738 21049
rect 17682 20975 17738 20984
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17684 20392 17736 20398
rect 17788 20380 17816 21422
rect 17880 21146 17908 23598
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17972 21690 18000 22442
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17972 21010 18000 21626
rect 17960 21004 18012 21010
rect 17960 20946 18012 20952
rect 17736 20352 17816 20380
rect 17684 20334 17736 20340
rect 17684 19372 17736 19378
rect 17684 19314 17736 19320
rect 17696 19174 17724 19314
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17788 18834 17816 20352
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 18290 17816 18770
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17880 18154 17908 19246
rect 17972 18222 18000 20946
rect 17960 18216 18012 18222
rect 18064 18193 18092 24142
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18524 23254 18552 23462
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 18616 22506 18644 24210
rect 18708 23769 18736 24618
rect 18800 24614 18828 25486
rect 18892 25362 18920 25774
rect 18972 25764 19024 25770
rect 19062 25735 19118 25744
rect 18972 25706 19024 25712
rect 18984 25673 19012 25706
rect 18970 25664 19026 25673
rect 18970 25599 19026 25608
rect 18880 25356 18932 25362
rect 18880 25298 18932 25304
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 19076 24342 19104 25735
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19904 25226 19932 26386
rect 20180 25838 20208 27474
rect 20456 27334 20484 27474
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 20168 25832 20220 25838
rect 20168 25774 20220 25780
rect 19892 25220 19944 25226
rect 19892 25162 19944 25168
rect 20180 24886 20208 25774
rect 20168 24880 20220 24886
rect 20168 24822 20220 24828
rect 20548 24818 20576 27968
rect 20628 27950 20680 27956
rect 20720 28008 20772 28014
rect 20720 27950 20772 27956
rect 20628 27328 20680 27334
rect 20628 27270 20680 27276
rect 20640 25430 20668 27270
rect 20732 26790 20760 27950
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20824 26568 20852 28902
rect 20916 27826 20944 29038
rect 21008 28966 21036 29192
rect 21088 29096 21140 29102
rect 21088 29038 21140 29044
rect 20996 28960 21048 28966
rect 20996 28902 21048 28908
rect 21008 28762 21036 28902
rect 20996 28756 21048 28762
rect 20996 28698 21048 28704
rect 21100 28218 21128 29038
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21180 28620 21232 28626
rect 21180 28562 21232 28568
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 20916 27798 21036 27826
rect 21008 27674 21036 27798
rect 21192 27674 21220 28562
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 21180 27668 21232 27674
rect 21180 27610 21232 27616
rect 20732 26540 20852 26568
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 18694 23760 18750 23769
rect 18694 23695 18750 23704
rect 20088 23662 20116 24550
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20076 23656 20128 23662
rect 20076 23598 20128 23604
rect 19432 23588 19484 23594
rect 19432 23530 19484 23536
rect 18788 23044 18840 23050
rect 18788 22986 18840 22992
rect 18800 22930 18828 22986
rect 18708 22902 18828 22930
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 18708 22710 18736 22902
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18788 22704 18840 22710
rect 18788 22646 18840 22652
rect 18604 22500 18656 22506
rect 18604 22442 18656 22448
rect 18800 22438 18828 22646
rect 19076 22642 19104 22918
rect 19064 22636 19116 22642
rect 19064 22578 19116 22584
rect 18972 22568 19024 22574
rect 18972 22510 19024 22516
rect 18984 22438 19012 22510
rect 18788 22432 18840 22438
rect 18788 22374 18840 22380
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18234 22128 18290 22137
rect 18234 22063 18236 22072
rect 18288 22063 18290 22072
rect 18512 22092 18564 22098
rect 18236 22034 18288 22040
rect 18512 22034 18564 22040
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18144 21888 18196 21894
rect 18142 21856 18144 21865
rect 18196 21856 18198 21865
rect 18142 21791 18198 21800
rect 18340 21486 18368 21966
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18524 20398 18552 22034
rect 18800 21690 18828 22374
rect 18788 21684 18840 21690
rect 18788 21626 18840 21632
rect 19168 20942 19196 22918
rect 19340 22704 19392 22710
rect 19338 22672 19340 22681
rect 19392 22672 19394 22681
rect 19338 22607 19394 22616
rect 19340 22568 19392 22574
rect 19340 22510 19392 22516
rect 19352 22137 19380 22510
rect 19338 22128 19394 22137
rect 19338 22063 19394 22072
rect 19352 21690 19380 22063
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19246 21040 19302 21049
rect 19246 20975 19248 20984
rect 19300 20975 19302 20984
rect 19248 20946 19300 20952
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18892 19922 18920 20402
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 18222 18276 19654
rect 18892 19310 18920 19858
rect 18972 19712 19024 19718
rect 18972 19654 19024 19660
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18432 18358 18460 19246
rect 18984 19174 19012 19654
rect 19076 19514 19104 19654
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 19352 19394 19380 21490
rect 19260 19366 19380 19394
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 18972 18828 19024 18834
rect 18972 18770 19024 18776
rect 18984 18426 19012 18770
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 19168 18222 19196 19110
rect 19260 18902 19288 19366
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 18970 19380 19246
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 18236 18216 18288 18222
rect 17960 18158 18012 18164
rect 18050 18184 18106 18193
rect 17868 18148 17920 18154
rect 18236 18158 18288 18164
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 18050 18119 18106 18128
rect 17868 18090 17920 18096
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16046 14780 17002
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 15028 5574 15056 15914
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 14752 3602 14780 5510
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 11072 2582 11100 3470
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 4172 2394 4200 2450
rect 4080 2366 4200 2394
rect 4080 1986 4108 2366
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4080 1958 4200 1986
rect 4172 800 4200 1958
rect 5092 800 5120 2450
rect 6012 800 6040 2450
rect 6932 800 6960 2450
rect 7852 800 7880 2450
rect 8772 800 8800 2450
rect 9692 800 9720 2450
rect 10612 800 10640 2450
rect 11532 800 11560 2450
rect 12452 800 12480 2450
rect 13372 800 13400 2450
rect 14292 800 14320 2450
rect 15212 800 15240 2450
rect 16132 800 16160 2450
rect 17052 800 17080 2450
rect 17972 800 18000 2450
rect 18892 800 18920 2450
rect 19444 2310 19472 23530
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 20180 23186 20208 24006
rect 20364 23866 20392 24142
rect 20548 24070 20576 24754
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20536 24064 20588 24070
rect 20536 24006 20588 24012
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19996 22778 20024 23054
rect 20088 22953 20116 23122
rect 20074 22944 20130 22953
rect 20074 22879 20130 22888
rect 20364 22778 20392 23530
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 19524 22704 19576 22710
rect 19524 22646 19576 22652
rect 19536 22574 19564 22646
rect 19524 22568 19576 22574
rect 19812 22545 19840 22714
rect 20076 22568 20128 22574
rect 19524 22510 19576 22516
rect 19798 22536 19854 22545
rect 20076 22510 20128 22516
rect 19798 22471 19854 22480
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 20088 22098 20116 22510
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19720 21554 19748 21966
rect 20180 21894 20208 22714
rect 20456 22658 20484 23054
rect 20364 22630 20484 22658
rect 20364 22506 20392 22630
rect 20444 22568 20496 22574
rect 20444 22510 20496 22516
rect 20352 22500 20404 22506
rect 20352 22442 20404 22448
rect 20456 22030 20484 22510
rect 20444 22024 20496 22030
rect 20444 21966 20496 21972
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20180 21570 20208 21830
rect 19708 21548 19760 21554
rect 19708 21490 19760 21496
rect 20088 21542 20208 21570
rect 19984 21480 20036 21486
rect 19904 21440 19984 21468
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19798 20904 19854 20913
rect 19720 20806 19748 20878
rect 19798 20839 19800 20848
rect 19852 20839 19854 20848
rect 19800 20810 19852 20816
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19614 20496 19670 20505
rect 19536 20398 19564 20470
rect 19614 20431 19670 20440
rect 19628 20398 19656 20431
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19904 19718 19932 21440
rect 19984 21422 20036 21428
rect 20088 21350 20116 21542
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19984 21344 20036 21350
rect 20076 21344 20128 21350
rect 19984 21286 20036 21292
rect 20074 21312 20076 21321
rect 20128 21312 20130 21321
rect 19996 20466 20024 21286
rect 20074 21247 20130 21256
rect 20076 21140 20128 21146
rect 20180 21128 20208 21422
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20272 21146 20300 21354
rect 20128 21100 20208 21128
rect 20076 21082 20128 21088
rect 20076 20868 20128 20874
rect 20076 20810 20128 20816
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20088 20346 20116 20810
rect 20180 20398 20208 21100
rect 20260 21140 20312 21146
rect 20260 21082 20312 21088
rect 20258 21040 20314 21049
rect 20258 20975 20314 20984
rect 19996 20318 20116 20346
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19996 19786 20024 20318
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19310 19932 19654
rect 19892 19304 19944 19310
rect 19522 19272 19578 19281
rect 19892 19246 19944 19252
rect 19522 19207 19524 19216
rect 19576 19207 19578 19216
rect 19524 19178 19576 19184
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19996 18442 20024 19722
rect 20088 19514 20116 20198
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20088 18970 20116 19450
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 20088 18698 20116 18906
rect 20272 18714 20300 20975
rect 20364 20942 20392 21830
rect 20456 21690 20484 21966
rect 20444 21684 20496 21690
rect 20444 21626 20496 21632
rect 20640 21570 20668 24210
rect 20732 23882 20760 26540
rect 20812 26444 20864 26450
rect 20812 26386 20864 26392
rect 20824 24750 20852 26386
rect 21008 26058 21036 27610
rect 21192 27538 21220 27610
rect 21180 27532 21232 27538
rect 21180 27474 21232 27480
rect 21284 27470 21312 28970
rect 21836 28762 21864 29242
rect 21824 28756 21876 28762
rect 21824 28698 21876 28704
rect 21836 27946 21864 28698
rect 22020 28626 22048 30262
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 21364 27940 21416 27946
rect 21364 27882 21416 27888
rect 21824 27940 21876 27946
rect 21824 27882 21876 27888
rect 21376 27538 21404 27882
rect 21364 27532 21416 27538
rect 21364 27474 21416 27480
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21180 27396 21232 27402
rect 21180 27338 21232 27344
rect 21456 27396 21508 27402
rect 21456 27338 21508 27344
rect 21086 27024 21142 27033
rect 21086 26959 21088 26968
rect 21140 26959 21142 26968
rect 21088 26930 21140 26936
rect 21088 26444 21140 26450
rect 21088 26386 21140 26392
rect 21100 26246 21128 26386
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 20916 26030 21036 26058
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20916 24070 20944 26030
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 21008 24682 21036 25774
rect 21088 24948 21140 24954
rect 21088 24890 21140 24896
rect 20996 24676 21048 24682
rect 20996 24618 21048 24624
rect 21100 24562 21128 24890
rect 21008 24534 21128 24562
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20732 23854 20852 23882
rect 20718 23216 20774 23225
rect 20718 23151 20720 23160
rect 20772 23151 20774 23160
rect 20720 23122 20772 23128
rect 20720 22432 20772 22438
rect 20824 22409 20852 23854
rect 20720 22374 20772 22380
rect 20810 22400 20866 22409
rect 20732 22030 20760 22374
rect 20810 22335 20866 22344
rect 20916 22094 20944 24006
rect 21008 22574 21036 24534
rect 21192 24342 21220 27338
rect 21468 27130 21496 27338
rect 21456 27124 21508 27130
rect 21456 27066 21508 27072
rect 21822 27024 21878 27033
rect 21822 26959 21878 26968
rect 21364 26920 21416 26926
rect 21362 26888 21364 26897
rect 21416 26888 21418 26897
rect 21362 26823 21418 26832
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21376 26586 21404 26726
rect 21836 26586 21864 26959
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 21456 26444 21508 26450
rect 21824 26444 21876 26450
rect 21456 26386 21508 26392
rect 21744 26404 21824 26432
rect 21272 26240 21324 26246
rect 21272 26182 21324 26188
rect 21284 26081 21312 26182
rect 21270 26072 21326 26081
rect 21270 26007 21326 26016
rect 21364 25968 21416 25974
rect 21362 25936 21364 25945
rect 21416 25936 21418 25945
rect 21362 25871 21418 25880
rect 21468 25838 21496 26386
rect 21640 26240 21692 26246
rect 21640 26182 21692 26188
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21456 25832 21508 25838
rect 21456 25774 21508 25780
rect 21376 25498 21404 25774
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21652 25430 21680 26182
rect 21640 25424 21692 25430
rect 21640 25366 21692 25372
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21180 24336 21232 24342
rect 21180 24278 21232 24284
rect 21468 23594 21496 24686
rect 21560 23798 21588 25230
rect 21744 24750 21772 26404
rect 21824 26386 21876 26392
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21836 24818 21864 26250
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21548 23792 21600 23798
rect 21548 23734 21600 23740
rect 21456 23588 21508 23594
rect 21456 23530 21508 23536
rect 21560 23118 21588 23734
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 20916 22066 21036 22094
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20548 21542 20668 21570
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20444 20936 20496 20942
rect 20444 20878 20496 20884
rect 20456 19446 20484 20878
rect 20548 20641 20576 21542
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20534 20632 20590 20641
rect 20534 20567 20590 20576
rect 20548 20466 20576 20567
rect 20640 20466 20668 21422
rect 20732 20874 20760 21966
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20824 21146 20852 21422
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20916 20505 20944 21830
rect 21008 20534 21036 22066
rect 20996 20528 21048 20534
rect 20902 20496 20958 20505
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20628 20460 20680 20466
rect 20996 20470 21048 20476
rect 20902 20431 20958 20440
rect 20628 20402 20680 20408
rect 20534 20360 20590 20369
rect 20640 20346 20668 20402
rect 20904 20392 20956 20398
rect 20640 20318 20760 20346
rect 20904 20334 20956 20340
rect 20534 20295 20590 20304
rect 20548 19922 20576 20295
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20640 19854 20668 20198
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20732 19786 20760 20318
rect 20916 20262 20944 20334
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 21100 20074 21128 22510
rect 21376 22506 21404 22918
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21376 21486 21404 22442
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21468 21162 21496 22510
rect 21376 21134 21496 21162
rect 21270 20632 21326 20641
rect 21270 20567 21326 20576
rect 21284 20534 21312 20567
rect 21272 20528 21324 20534
rect 21272 20470 21324 20476
rect 21180 20324 21232 20330
rect 21180 20266 21232 20272
rect 20916 20046 21128 20074
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20732 19514 20760 19722
rect 20824 19514 20852 19858
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20916 19310 20944 20046
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 21008 18970 21036 19858
rect 21192 19174 21220 20266
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21284 19786 21312 20198
rect 21272 19780 21324 19786
rect 21272 19722 21324 19728
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 21192 18834 21220 19110
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 20996 18760 21048 18766
rect 20076 18692 20128 18698
rect 20272 18686 20392 18714
rect 20996 18702 21048 18708
rect 20076 18634 20128 18640
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 19996 18414 20116 18442
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19996 17746 20024 18226
rect 20088 17882 20116 18414
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20180 17814 20208 18022
rect 20168 17808 20220 17814
rect 20168 17750 20220 17756
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 20364 17202 20392 18686
rect 21008 18154 21036 18702
rect 21376 18426 21404 21134
rect 21560 21078 21588 23054
rect 21652 22574 21680 23462
rect 21744 23338 21772 24686
rect 21928 24342 21956 27406
rect 22020 26897 22048 27474
rect 22006 26888 22062 26897
rect 22006 26823 22062 26832
rect 22020 26382 22048 26823
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 22112 25158 22140 31282
rect 22204 27033 22232 32914
rect 22664 32910 22692 33390
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 22652 32904 22704 32910
rect 22652 32846 22704 32852
rect 22664 32774 22692 32846
rect 22848 32774 22876 32914
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22836 32768 22888 32774
rect 22836 32710 22888 32716
rect 22836 32360 22888 32366
rect 22836 32302 22888 32308
rect 22560 32292 22612 32298
rect 22560 32234 22612 32240
rect 22572 31890 22600 32234
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22560 31884 22612 31890
rect 22560 31826 22612 31832
rect 22480 31210 22508 31826
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22468 31204 22520 31210
rect 22468 31146 22520 31152
rect 22480 30938 22508 31146
rect 22468 30932 22520 30938
rect 22468 30874 22520 30880
rect 22376 30796 22428 30802
rect 22376 30738 22428 30744
rect 22284 30184 22336 30190
rect 22284 30126 22336 30132
rect 22296 29578 22324 30126
rect 22388 30054 22416 30738
rect 22468 30660 22520 30666
rect 22468 30602 22520 30608
rect 22480 30161 22508 30602
rect 22466 30152 22522 30161
rect 22664 30122 22692 31758
rect 22756 31754 22784 31894
rect 22744 31748 22796 31754
rect 22744 31690 22796 31696
rect 22756 31278 22784 31690
rect 22848 31414 22876 32302
rect 22836 31408 22888 31414
rect 22836 31350 22888 31356
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 22466 30087 22522 30096
rect 22652 30116 22704 30122
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22284 29572 22336 29578
rect 22284 29514 22336 29520
rect 22296 28558 22324 29514
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22296 28014 22324 28494
rect 22284 28008 22336 28014
rect 22284 27950 22336 27956
rect 22284 27600 22336 27606
rect 22284 27542 22336 27548
rect 22190 27024 22246 27033
rect 22190 26959 22246 26968
rect 22296 26790 22324 27542
rect 22284 26784 22336 26790
rect 22284 26726 22336 26732
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22204 25702 22232 26386
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 22204 25498 22232 25638
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21836 23526 21864 24278
rect 21914 24168 21970 24177
rect 22020 24138 22048 24618
rect 21914 24103 21916 24112
rect 21968 24103 21970 24112
rect 22008 24132 22060 24138
rect 21916 24074 21968 24080
rect 22008 24074 22060 24080
rect 22296 23662 22324 25774
rect 22388 25430 22416 29990
rect 22480 25809 22508 30087
rect 22652 30058 22704 30064
rect 22664 29714 22692 30058
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22652 29572 22704 29578
rect 22652 29514 22704 29520
rect 22560 29300 22612 29306
rect 22664 29288 22692 29514
rect 22612 29260 22692 29288
rect 22560 29242 22612 29248
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22664 29034 22692 29106
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22560 28960 22612 28966
rect 22560 28902 22612 28908
rect 22572 28626 22600 28902
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 22572 27946 22600 28562
rect 22756 28490 22784 29990
rect 22940 29646 22968 33866
rect 23124 32978 23152 33934
rect 23400 33114 23428 34002
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33318 23704 33798
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 23940 33380 23992 33386
rect 23940 33322 23992 33328
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23112 32972 23164 32978
rect 23112 32914 23164 32920
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23308 32502 23336 32710
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23480 32360 23532 32366
rect 23110 32328 23166 32337
rect 23480 32302 23532 32308
rect 23110 32263 23112 32272
rect 23164 32263 23166 32272
rect 23112 32234 23164 32240
rect 23020 31680 23072 31686
rect 23020 31622 23072 31628
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22848 28694 22876 29446
rect 22928 29028 22980 29034
rect 22928 28970 22980 28976
rect 22940 28762 22968 28970
rect 22928 28756 22980 28762
rect 22928 28698 22980 28704
rect 22836 28688 22888 28694
rect 22836 28630 22888 28636
rect 22744 28484 22796 28490
rect 22744 28426 22796 28432
rect 22560 27940 22612 27946
rect 22560 27882 22612 27888
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 22664 25838 22692 26862
rect 23032 26858 23060 31622
rect 23124 31278 23152 32234
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23308 30802 23336 31078
rect 23296 30796 23348 30802
rect 23296 30738 23348 30744
rect 23204 30184 23256 30190
rect 23204 30126 23256 30132
rect 23216 29170 23244 30126
rect 23400 29730 23428 31826
rect 23492 31754 23520 32302
rect 23584 32298 23612 32982
rect 23572 32292 23624 32298
rect 23572 32234 23624 32240
rect 23480 31748 23532 31754
rect 23480 31690 23532 31696
rect 23492 31346 23520 31690
rect 23676 31482 23704 33254
rect 23952 33114 23980 33322
rect 24860 33312 24912 33318
rect 24860 33254 24912 33260
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23848 32972 23900 32978
rect 23848 32914 23900 32920
rect 24032 32972 24084 32978
rect 24032 32914 24084 32920
rect 23860 31822 23888 32914
rect 23940 32360 23992 32366
rect 24044 32337 24072 32914
rect 24872 32774 24900 33254
rect 24964 32978 24992 33390
rect 24952 32972 25004 32978
rect 24952 32914 25004 32920
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24964 32366 24992 32914
rect 25700 32434 25728 34002
rect 26148 33312 26200 33318
rect 26148 33254 26200 33260
rect 25780 32972 25832 32978
rect 25780 32914 25832 32920
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 24952 32360 25004 32366
rect 23940 32302 23992 32308
rect 24030 32328 24086 32337
rect 23848 31816 23900 31822
rect 23848 31758 23900 31764
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 23480 31340 23532 31346
rect 23480 31282 23532 31288
rect 23480 31204 23532 31210
rect 23480 31146 23532 31152
rect 23308 29702 23428 29730
rect 23492 29714 23520 31146
rect 23676 30954 23704 31418
rect 23860 31278 23888 31758
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23584 30926 23704 30954
rect 23584 30190 23612 30926
rect 23664 30796 23716 30802
rect 23664 30738 23716 30744
rect 23676 30394 23704 30738
rect 23952 30734 23980 32302
rect 24952 32302 25004 32308
rect 25412 32360 25464 32366
rect 25412 32302 25464 32308
rect 24030 32263 24032 32272
rect 24084 32263 24086 32272
rect 24032 32234 24084 32240
rect 24964 32026 24992 32302
rect 24952 32020 25004 32026
rect 24952 31962 25004 31968
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 24492 30728 24544 30734
rect 24492 30670 24544 30676
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23664 30388 23716 30394
rect 23664 30330 23716 30336
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 23480 29708 23532 29714
rect 23308 29220 23336 29702
rect 23480 29650 23532 29656
rect 23308 29192 23612 29220
rect 23112 29164 23164 29170
rect 23112 29106 23164 29112
rect 23204 29164 23256 29170
rect 23204 29106 23256 29112
rect 23124 28218 23152 29106
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 23478 29064 23534 29073
rect 23308 28966 23336 29038
rect 23478 28999 23480 29008
rect 23532 28999 23534 29008
rect 23480 28970 23532 28976
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 23204 28416 23256 28422
rect 23204 28358 23256 28364
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23216 28014 23244 28358
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23204 28008 23256 28014
rect 23204 27950 23256 27956
rect 23216 27470 23244 27950
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23020 26852 23072 26858
rect 23020 26794 23072 26800
rect 23400 26586 23428 28018
rect 23492 27946 23520 28562
rect 23480 27940 23532 27946
rect 23480 27882 23532 27888
rect 23492 27538 23520 27882
rect 23584 27606 23612 29192
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 22652 25832 22704 25838
rect 22466 25800 22522 25809
rect 22652 25774 22704 25780
rect 23296 25832 23348 25838
rect 23296 25774 23348 25780
rect 22466 25735 22522 25744
rect 22376 25424 22428 25430
rect 22376 25366 22428 25372
rect 22480 24818 22508 25735
rect 22836 25492 22888 25498
rect 22836 25434 22888 25440
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22848 24274 22876 25434
rect 23308 24721 23336 25774
rect 23294 24712 23350 24721
rect 23400 24682 23428 26386
rect 23492 25498 23520 27474
rect 23676 26518 23704 30330
rect 23768 30190 23796 30534
rect 24504 30326 24532 30670
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 23756 30184 23808 30190
rect 23756 30126 23808 30132
rect 24492 30116 24544 30122
rect 24492 30058 24544 30064
rect 23940 29640 23992 29646
rect 23940 29582 23992 29588
rect 23756 29028 23808 29034
rect 23756 28970 23808 28976
rect 23768 28694 23796 28970
rect 23848 28960 23900 28966
rect 23848 28902 23900 28908
rect 23756 28688 23808 28694
rect 23756 28630 23808 28636
rect 23860 28014 23888 28902
rect 23952 28626 23980 29582
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 24044 28694 24072 29446
rect 24504 29102 24532 30058
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24492 29096 24544 29102
rect 24492 29038 24544 29044
rect 24596 29034 24624 29242
rect 24584 29028 24636 29034
rect 24584 28970 24636 28976
rect 24032 28688 24084 28694
rect 24032 28630 24084 28636
rect 23940 28620 23992 28626
rect 23940 28562 23992 28568
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23848 28008 23900 28014
rect 23848 27950 23900 27956
rect 23664 26512 23716 26518
rect 23664 26454 23716 26460
rect 23676 26353 23704 26454
rect 23662 26344 23718 26353
rect 23662 26279 23718 26288
rect 23664 26240 23716 26246
rect 23664 26182 23716 26188
rect 23480 25492 23532 25498
rect 23480 25434 23532 25440
rect 23572 25356 23624 25362
rect 23572 25298 23624 25304
rect 23294 24647 23350 24656
rect 23388 24676 23440 24682
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22192 23656 22244 23662
rect 22192 23598 22244 23604
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 21824 23520 21876 23526
rect 22204 23497 22232 23598
rect 22664 23594 22692 24210
rect 23112 24064 23164 24070
rect 23112 24006 23164 24012
rect 22836 23656 22888 23662
rect 22836 23598 22888 23604
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 21824 23462 21876 23468
rect 22190 23488 22246 23497
rect 22190 23423 22246 23432
rect 21744 23310 21864 23338
rect 21836 23225 21864 23310
rect 21822 23216 21878 23225
rect 21732 23180 21784 23186
rect 21822 23151 21878 23160
rect 21732 23122 21784 23128
rect 21744 22778 21772 23122
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22664 22574 22692 23530
rect 22848 23186 22876 23598
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 21640 22568 21692 22574
rect 21640 22510 21692 22516
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 21638 22400 21694 22409
rect 21638 22335 21694 22344
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21548 20460 21600 20466
rect 21548 20402 21600 20408
rect 21456 19984 21508 19990
rect 21456 19926 21508 19932
rect 21468 19786 21496 19926
rect 21456 19780 21508 19786
rect 21456 19722 21508 19728
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21468 18358 21496 19246
rect 21560 18698 21588 20402
rect 21652 18766 21680 22335
rect 22192 22160 22244 22166
rect 21822 22128 21878 22137
rect 22192 22102 22244 22108
rect 22926 22128 22982 22137
rect 21822 22063 21824 22072
rect 21876 22063 21878 22072
rect 21824 22034 21876 22040
rect 22204 20262 22232 22102
rect 22560 22092 22612 22098
rect 22926 22063 22982 22072
rect 22560 22034 22612 22040
rect 22572 21622 22600 22034
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22192 20256 22244 20262
rect 22192 20198 22244 20204
rect 22204 19990 22232 20198
rect 22192 19984 22244 19990
rect 22192 19926 22244 19932
rect 21732 19916 21784 19922
rect 21732 19858 21784 19864
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21744 19514 21772 19858
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21928 19310 21956 19858
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 22664 18902 22692 19654
rect 22848 19310 22876 21966
rect 22940 21486 22968 22063
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23124 21842 23152 24006
rect 23308 23798 23336 24647
rect 23388 24618 23440 24624
rect 23584 24070 23612 25298
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23866 23612 24006
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 23308 23662 23336 23734
rect 23296 23656 23348 23662
rect 23400 23633 23428 23802
rect 23676 23746 23704 26182
rect 23492 23718 23704 23746
rect 23296 23598 23348 23604
rect 23386 23624 23442 23633
rect 23386 23559 23442 23568
rect 23032 21706 23060 21830
rect 23124 21814 23244 21842
rect 23032 21678 23152 21706
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 23032 20602 23060 21490
rect 23124 21486 23152 21678
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 23124 21146 23152 21422
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23020 20596 23072 20602
rect 23020 20538 23072 20544
rect 22940 19961 22968 20538
rect 22926 19952 22982 19961
rect 23216 19922 23244 21814
rect 23492 21486 23520 23718
rect 23846 23216 23902 23225
rect 23846 23151 23848 23160
rect 23900 23151 23902 23160
rect 23848 23122 23900 23128
rect 23952 23066 23980 28426
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24136 27130 24164 27474
rect 24688 27130 24716 31214
rect 24780 27606 24808 31758
rect 25424 30054 25452 32302
rect 25792 32230 25820 32914
rect 26160 32366 26188 33254
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25780 31952 25832 31958
rect 25780 31894 25832 31900
rect 25504 30660 25556 30666
rect 25504 30602 25556 30608
rect 25516 30394 25544 30602
rect 25504 30388 25556 30394
rect 25504 30330 25556 30336
rect 25792 30190 25820 31894
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 27804 31884 27856 31890
rect 27804 31826 27856 31832
rect 25964 31204 26016 31210
rect 25964 31146 26016 31152
rect 25976 30938 26004 31146
rect 25964 30932 26016 30938
rect 25964 30874 26016 30880
rect 26344 30326 26372 31826
rect 27068 31816 27120 31822
rect 27068 31758 27120 31764
rect 27080 31482 27108 31758
rect 27816 31482 27844 31826
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 27068 31476 27120 31482
rect 27068 31418 27120 31424
rect 27252 31476 27304 31482
rect 27252 31418 27304 31424
rect 27804 31476 27856 31482
rect 27804 31418 27856 31424
rect 26516 31136 26568 31142
rect 26516 31078 26568 31084
rect 26528 30802 26556 31078
rect 26516 30796 26568 30802
rect 26516 30738 26568 30744
rect 26976 30796 27028 30802
rect 26976 30738 27028 30744
rect 26332 30320 26384 30326
rect 26332 30262 26384 30268
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 26056 30184 26108 30190
rect 26056 30126 26108 30132
rect 25412 30048 25464 30054
rect 25412 29990 25464 29996
rect 25044 29708 25096 29714
rect 25044 29650 25096 29656
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 24872 29170 24900 29446
rect 24964 29238 24992 29582
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 24872 28762 24900 29106
rect 25056 29102 25084 29650
rect 25320 29504 25372 29510
rect 25320 29446 25372 29452
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25044 29096 25096 29102
rect 25044 29038 25096 29044
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 25240 26858 25268 28018
rect 25332 27878 25360 29446
rect 25780 29232 25832 29238
rect 25780 29174 25832 29180
rect 25688 28620 25740 28626
rect 25688 28562 25740 28568
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25608 26994 25636 28358
rect 25700 28014 25728 28562
rect 25688 28008 25740 28014
rect 25688 27950 25740 27956
rect 25700 27402 25728 27950
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 24584 26852 24636 26858
rect 24584 26794 24636 26800
rect 25228 26852 25280 26858
rect 25228 26794 25280 26800
rect 24596 25702 24624 26794
rect 25240 26042 25268 26794
rect 25608 26586 25636 26930
rect 25792 26926 25820 29174
rect 25884 29102 25912 29446
rect 25872 29096 25924 29102
rect 25872 29038 25924 29044
rect 26068 28558 26096 30126
rect 26240 29708 26292 29714
rect 26240 29650 26292 29656
rect 26148 29096 26200 29102
rect 26148 29038 26200 29044
rect 26252 29050 26280 29650
rect 26344 29238 26372 30262
rect 26528 30190 26556 30738
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26792 30592 26844 30598
rect 26792 30534 26844 30540
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 26516 30184 26568 30190
rect 26516 30126 26568 30132
rect 26620 29714 26648 30262
rect 26712 30190 26740 30534
rect 26700 30184 26752 30190
rect 26700 30126 26752 30132
rect 26804 30002 26832 30534
rect 26988 30326 27016 30738
rect 27264 30734 27292 31418
rect 28172 31272 28224 31278
rect 28172 31214 28224 31220
rect 27252 30728 27304 30734
rect 27252 30670 27304 30676
rect 26976 30320 27028 30326
rect 26976 30262 27028 30268
rect 26712 29974 26832 30002
rect 26712 29714 26740 29974
rect 26424 29708 26476 29714
rect 26424 29650 26476 29656
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26700 29708 26752 29714
rect 26700 29650 26752 29656
rect 26332 29232 26384 29238
rect 26332 29174 26384 29180
rect 26436 29102 26464 29650
rect 26712 29102 26740 29650
rect 26332 29096 26384 29102
rect 26252 29044 26332 29050
rect 26252 29038 26384 29044
rect 26424 29096 26476 29102
rect 26424 29038 26476 29044
rect 26700 29096 26752 29102
rect 26700 29038 26752 29044
rect 26056 28552 26108 28558
rect 26056 28494 26108 28500
rect 25872 28416 25924 28422
rect 25872 28358 25924 28364
rect 25884 28218 25912 28358
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 26068 28082 26096 28494
rect 26160 28218 26188 29038
rect 26252 29022 26372 29038
rect 26344 28778 26372 29022
rect 26344 28750 26464 28778
rect 26148 28212 26200 28218
rect 26148 28154 26200 28160
rect 26240 28144 26292 28150
rect 26240 28086 26292 28092
rect 26332 28144 26384 28150
rect 26332 28086 26384 28092
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26056 27940 26108 27946
rect 26056 27882 26108 27888
rect 25872 27396 25924 27402
rect 25872 27338 25924 27344
rect 25884 27130 25912 27338
rect 25964 27328 26016 27334
rect 25964 27270 26016 27276
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25780 26920 25832 26926
rect 25780 26862 25832 26868
rect 25596 26580 25648 26586
rect 25596 26522 25648 26528
rect 25792 26382 25820 26862
rect 25976 26518 26004 27270
rect 26068 27130 26096 27882
rect 26160 27878 26188 27950
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26148 27532 26200 27538
rect 26148 27474 26200 27480
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 25964 26512 26016 26518
rect 25964 26454 26016 26460
rect 25780 26376 25832 26382
rect 25780 26318 25832 26324
rect 25504 26240 25556 26246
rect 25504 26182 25556 26188
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 24584 25696 24636 25702
rect 24584 25638 24636 25644
rect 24596 24954 24624 25638
rect 25516 25362 25544 26182
rect 25792 26042 25820 26318
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25780 26036 25832 26042
rect 25780 25978 25832 25984
rect 25504 25356 25556 25362
rect 25504 25298 25556 25304
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 24584 24948 24636 24954
rect 24584 24890 24636 24896
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24400 24608 24452 24614
rect 24400 24550 24452 24556
rect 24412 24410 24440 24550
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24216 23656 24268 23662
rect 24216 23598 24268 23604
rect 24228 23497 24256 23598
rect 24214 23488 24270 23497
rect 24214 23423 24270 23432
rect 24216 23180 24268 23186
rect 24216 23122 24268 23128
rect 24308 23180 24360 23186
rect 24308 23122 24360 23128
rect 23860 23038 23980 23066
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 23860 22438 23888 23038
rect 24044 22778 24072 23054
rect 24228 22982 24256 23122
rect 24320 23089 24348 23122
rect 24306 23080 24362 23089
rect 24306 23015 24362 23024
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 24032 22772 24084 22778
rect 24032 22714 24084 22720
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 24030 22536 24086 22545
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23952 22166 23980 22510
rect 24030 22471 24086 22480
rect 23940 22160 23992 22166
rect 23940 22102 23992 22108
rect 23572 21956 23624 21962
rect 23572 21898 23624 21904
rect 23584 21865 23612 21898
rect 23570 21856 23626 21865
rect 23570 21791 23626 21800
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23492 20602 23520 21422
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21078 23704 21286
rect 23860 21146 23888 21490
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23296 20392 23348 20398
rect 23572 20392 23624 20398
rect 23296 20334 23348 20340
rect 23570 20360 23572 20369
rect 23624 20360 23626 20369
rect 22926 19887 22982 19896
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22652 18896 22704 18902
rect 22652 18838 22704 18844
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21376 17882 21404 18226
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 21376 17134 21404 17818
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 21560 16726 21588 18634
rect 21652 18154 21680 18702
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21836 18290 21864 18566
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21640 18148 21692 18154
rect 21640 18090 21692 18096
rect 21652 17338 21680 18090
rect 21836 17746 21864 18226
rect 21928 18086 21956 18770
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 22020 18358 22048 18702
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 22848 18222 22876 19246
rect 23032 18630 23060 19858
rect 23308 19514 23336 20334
rect 23570 20295 23626 20304
rect 23664 20324 23716 20330
rect 23584 19922 23612 20295
rect 23664 20266 23716 20272
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23492 19310 23520 19654
rect 23480 19304 23532 19310
rect 23480 19246 23532 19252
rect 23492 18834 23520 19246
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 22836 18216 22888 18222
rect 22836 18158 22888 18164
rect 21916 18080 21968 18086
rect 21916 18022 21968 18028
rect 21928 17882 21956 18022
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22848 17746 22876 18158
rect 23400 17814 23428 18226
rect 23492 17882 23520 18770
rect 23676 18426 23704 20266
rect 23860 19310 23888 21082
rect 23952 20602 23980 22102
rect 24044 21690 24072 22471
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24228 21486 24256 22918
rect 24412 22574 24440 24346
rect 24504 22778 24532 24822
rect 25792 24750 25820 25094
rect 25504 24744 25556 24750
rect 25502 24712 25504 24721
rect 25780 24744 25832 24750
rect 25556 24712 25558 24721
rect 24584 24676 24636 24682
rect 24636 24636 24900 24664
rect 25558 24670 25636 24698
rect 25780 24686 25832 24692
rect 25502 24647 25558 24656
rect 24584 24618 24636 24624
rect 24872 23254 24900 24636
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 25042 23624 25098 23633
rect 25042 23559 25098 23568
rect 25056 23526 25084 23559
rect 25044 23520 25096 23526
rect 25044 23462 25096 23468
rect 24860 23248 24912 23254
rect 24860 23190 24912 23196
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21690 24440 21830
rect 24400 21684 24452 21690
rect 24400 21626 24452 21632
rect 24412 21554 24440 21626
rect 24400 21548 24452 21554
rect 24400 21490 24452 21496
rect 24216 21480 24268 21486
rect 24216 21422 24268 21428
rect 24400 21344 24452 21350
rect 24398 21312 24400 21321
rect 24452 21312 24454 21321
rect 24398 21247 24454 21256
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24044 19922 24072 20470
rect 24504 19990 24532 22714
rect 24584 22568 24636 22574
rect 24584 22510 24636 22516
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24596 20262 24624 22510
rect 24688 21321 24716 22510
rect 24860 22500 24912 22506
rect 24860 22442 24912 22448
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 24872 21418 24900 22442
rect 24860 21412 24912 21418
rect 24860 21354 24912 21360
rect 24674 21312 24730 21321
rect 24674 21247 24730 21256
rect 24964 21010 24992 22442
rect 25148 22438 25176 24006
rect 25320 23588 25372 23594
rect 25320 23530 25372 23536
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 22166 25176 22374
rect 25332 22166 25360 23530
rect 25424 22545 25452 24210
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25410 22536 25466 22545
rect 25410 22471 25466 22480
rect 25136 22160 25188 22166
rect 25136 22102 25188 22108
rect 25320 22160 25372 22166
rect 25320 22102 25372 22108
rect 25148 21486 25176 22102
rect 25516 22098 25544 23598
rect 25608 23118 25636 24670
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 25596 23112 25648 23118
rect 25596 23054 25648 23060
rect 25228 22092 25280 22098
rect 25228 22034 25280 22040
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25240 21622 25268 22034
rect 25608 22030 25636 23054
rect 25700 22982 25728 24210
rect 25884 23254 25912 26250
rect 26160 25974 26188 27474
rect 26148 25968 26200 25974
rect 26148 25910 26200 25916
rect 26252 25838 26280 28086
rect 26344 28014 26372 28086
rect 26332 28008 26384 28014
rect 26332 27950 26384 27956
rect 26436 27402 26464 28750
rect 26608 28144 26660 28150
rect 26608 28086 26660 28092
rect 26620 27538 26648 28086
rect 26608 27532 26660 27538
rect 26608 27474 26660 27480
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26424 27124 26476 27130
rect 26424 27066 26476 27072
rect 25964 25832 26016 25838
rect 26148 25832 26200 25838
rect 26016 25792 26096 25820
rect 25964 25774 26016 25780
rect 26068 25158 26096 25792
rect 26148 25774 26200 25780
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 26160 24954 26188 25774
rect 26436 25208 26464 27066
rect 26620 27062 26648 27474
rect 26608 27056 26660 27062
rect 26608 26998 26660 27004
rect 26516 26988 26568 26994
rect 26516 26930 26568 26936
rect 26528 26432 26556 26930
rect 26608 26444 26660 26450
rect 26528 26404 26608 26432
rect 26608 26386 26660 26392
rect 26514 26344 26570 26353
rect 26514 26279 26570 26288
rect 26528 25838 26556 26279
rect 26516 25832 26568 25838
rect 26516 25774 26568 25780
rect 26528 25430 26556 25774
rect 26516 25424 26568 25430
rect 26516 25366 26568 25372
rect 26516 25220 26568 25226
rect 26436 25180 26516 25208
rect 26516 25162 26568 25168
rect 26148 24948 26200 24954
rect 26148 24890 26200 24896
rect 26528 24721 26556 25162
rect 26514 24712 26570 24721
rect 26148 24676 26200 24682
rect 26514 24647 26570 24656
rect 26148 24618 26200 24624
rect 26160 23866 26188 24618
rect 26516 24200 26568 24206
rect 26516 24142 26568 24148
rect 26148 23860 26200 23866
rect 26148 23802 26200 23808
rect 25964 23520 26016 23526
rect 25964 23462 26016 23468
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25884 22574 25912 22714
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25700 22166 25728 22374
rect 25688 22160 25740 22166
rect 25688 22102 25740 22108
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25412 21412 25464 21418
rect 25412 21354 25464 21360
rect 25424 21146 25452 21354
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 25318 21040 25374 21049
rect 24952 21004 25004 21010
rect 25318 20975 25320 20984
rect 24952 20946 25004 20952
rect 25372 20975 25374 20984
rect 25320 20946 25372 20952
rect 25516 20618 25544 21286
rect 25424 20602 25544 20618
rect 25412 20596 25544 20602
rect 25464 20590 25544 20596
rect 25412 20538 25464 20544
rect 25516 20398 25544 20590
rect 25596 20460 25648 20466
rect 25596 20402 25648 20408
rect 25504 20392 25556 20398
rect 25504 20334 25556 20340
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24124 19984 24176 19990
rect 24124 19926 24176 19932
rect 24492 19984 24544 19990
rect 24492 19926 24544 19932
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23848 19304 23900 19310
rect 23848 19246 23900 19252
rect 23756 19236 23808 19242
rect 23756 19178 23808 19184
rect 23768 18902 23796 19178
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23860 18834 23888 19246
rect 24136 18834 24164 19926
rect 24596 19922 24624 20198
rect 24216 19916 24268 19922
rect 24216 19858 24268 19864
rect 24584 19916 24636 19922
rect 24584 19858 24636 19864
rect 25320 19916 25372 19922
rect 25320 19858 25372 19864
rect 25504 19916 25556 19922
rect 25608 19904 25636 20402
rect 25792 20074 25820 22510
rect 25872 21004 25924 21010
rect 25872 20946 25924 20952
rect 25884 20602 25912 20946
rect 25872 20596 25924 20602
rect 25872 20538 25924 20544
rect 25976 20448 26004 23462
rect 26160 22574 26188 23802
rect 26528 23798 26556 24142
rect 26516 23792 26568 23798
rect 26516 23734 26568 23740
rect 26332 23248 26384 23254
rect 26332 23190 26384 23196
rect 26148 22568 26200 22574
rect 25556 19876 25636 19904
rect 25700 20046 25820 20074
rect 25884 20420 26004 20448
rect 26068 22528 26148 22556
rect 25504 19858 25556 19864
rect 24228 19378 24256 19858
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24688 19514 24716 19654
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 24228 18630 24256 19314
rect 24676 19236 24728 19242
rect 24676 19178 24728 19184
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23388 17808 23440 17814
rect 23388 17750 23440 17756
rect 24044 17746 24072 18022
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 24032 17740 24084 17746
rect 24032 17682 24084 17688
rect 21640 17332 21692 17338
rect 21640 17274 21692 17280
rect 22848 17134 22876 17682
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 22836 17128 22888 17134
rect 22836 17070 22888 17076
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 22848 16658 22876 17070
rect 22836 16652 22888 16658
rect 22836 16594 22888 16600
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 23400 13258 23428 17138
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24136 16794 24164 17070
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24228 16658 24256 18566
rect 24688 18086 24716 19178
rect 24768 18148 24820 18154
rect 24768 18090 24820 18096
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24780 17338 24808 18090
rect 25148 17746 25176 19790
rect 25332 17882 25360 19858
rect 25516 19514 25544 19858
rect 25700 19786 25728 20046
rect 25778 19952 25834 19961
rect 25778 19887 25834 19896
rect 25792 19854 25820 19887
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25884 19666 25912 20420
rect 25792 19638 25912 19666
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25504 18624 25556 18630
rect 25504 18566 25556 18572
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25516 17814 25544 18566
rect 25792 18154 25820 19638
rect 26068 19334 26096 22528
rect 26148 22510 26200 22516
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 25976 19306 26096 19334
rect 25976 18834 26004 19306
rect 26160 18834 26188 19654
rect 25964 18828 26016 18834
rect 25964 18770 26016 18776
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 26148 18692 26200 18698
rect 26148 18634 26200 18640
rect 26160 18290 26188 18634
rect 26344 18426 26372 23190
rect 26528 23186 26556 23734
rect 26620 23730 26648 26386
rect 26712 24177 26740 29038
rect 26884 28620 26936 28626
rect 26884 28562 26936 28568
rect 26896 27674 26924 28562
rect 26884 27668 26936 27674
rect 26884 27610 26936 27616
rect 27160 27464 27212 27470
rect 27264 27452 27292 30670
rect 27988 30252 28040 30258
rect 27988 30194 28040 30200
rect 27436 30116 27488 30122
rect 27436 30058 27488 30064
rect 27344 29504 27396 29510
rect 27344 29446 27396 29452
rect 27356 28558 27384 29446
rect 27344 28552 27396 28558
rect 27344 28494 27396 28500
rect 27356 28014 27384 28494
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27448 27538 27476 30058
rect 28000 30054 28028 30194
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 27804 29708 27856 29714
rect 27804 29650 27856 29656
rect 27528 29232 27580 29238
rect 27528 29174 27580 29180
rect 27540 28218 27568 29174
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27632 28626 27660 28902
rect 27620 28620 27672 28626
rect 27620 28562 27672 28568
rect 27528 28212 27580 28218
rect 27528 28154 27580 28160
rect 27436 27532 27488 27538
rect 27436 27474 27488 27480
rect 27212 27424 27292 27452
rect 27160 27406 27212 27412
rect 27172 27130 27200 27406
rect 27724 27130 27752 28970
rect 27816 28694 27844 29650
rect 27896 29300 27948 29306
rect 27896 29242 27948 29248
rect 27804 28688 27856 28694
rect 27804 28630 27856 28636
rect 27908 28626 27936 29242
rect 28000 29102 28028 29990
rect 28184 29714 28212 31214
rect 28460 30190 28488 31622
rect 29828 30728 29880 30734
rect 29828 30670 29880 30676
rect 29840 30326 29868 30670
rect 30104 30592 30156 30598
rect 30104 30534 30156 30540
rect 28724 30320 28776 30326
rect 28724 30262 28776 30268
rect 29828 30320 29880 30326
rect 29828 30262 29880 30268
rect 28448 30184 28500 30190
rect 28448 30126 28500 30132
rect 28632 30184 28684 30190
rect 28632 30126 28684 30132
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 28264 30048 28316 30054
rect 28264 29990 28316 29996
rect 28276 29714 28304 29990
rect 28172 29708 28224 29714
rect 28172 29650 28224 29656
rect 28264 29708 28316 29714
rect 28264 29650 28316 29656
rect 28184 29594 28212 29650
rect 28184 29578 28304 29594
rect 28184 29572 28316 29578
rect 28184 29566 28264 29572
rect 28264 29514 28316 29520
rect 28080 29504 28132 29510
rect 28080 29446 28132 29452
rect 27988 29096 28040 29102
rect 27988 29038 28040 29044
rect 27896 28620 27948 28626
rect 27896 28562 27948 28568
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27160 27124 27212 27130
rect 27712 27124 27764 27130
rect 27212 27084 27292 27112
rect 27160 27066 27212 27072
rect 26792 26920 26844 26926
rect 26792 26862 26844 26868
rect 26804 26450 26832 26862
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 26884 26444 26936 26450
rect 26884 26386 26936 26392
rect 26792 25288 26844 25294
rect 26896 25242 26924 26386
rect 27264 26382 27292 27084
rect 27712 27066 27764 27072
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 26844 25236 26924 25242
rect 26792 25230 26924 25236
rect 26804 25214 26924 25230
rect 26896 24954 26924 25214
rect 26884 24948 26936 24954
rect 26884 24890 26936 24896
rect 26698 24168 26754 24177
rect 26698 24103 26754 24112
rect 26608 23724 26660 23730
rect 26608 23666 26660 23672
rect 26896 23662 26924 24890
rect 26884 23656 26936 23662
rect 26884 23598 26936 23604
rect 27172 23526 27200 26318
rect 27816 26314 27844 28426
rect 28092 28150 28120 29446
rect 28368 28966 28396 30058
rect 28460 29646 28488 30126
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28644 29306 28672 30126
rect 28736 30054 28764 30262
rect 29828 30184 29880 30190
rect 29826 30152 29828 30161
rect 30012 30184 30064 30190
rect 29880 30152 29882 30161
rect 30012 30126 30064 30132
rect 29826 30087 29882 30096
rect 30024 30054 30052 30126
rect 30116 30054 30144 30534
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 30012 30048 30064 30054
rect 30012 29990 30064 29996
rect 30104 30048 30156 30054
rect 30104 29990 30156 29996
rect 28632 29300 28684 29306
rect 28632 29242 28684 29248
rect 28736 29102 28764 29990
rect 28816 29708 28868 29714
rect 28816 29650 28868 29656
rect 28828 29306 28856 29650
rect 30392 29646 30420 52566
rect 30668 52562 30696 52838
rect 30656 52556 30708 52562
rect 30656 52498 30708 52504
rect 30564 51468 30616 51474
rect 30564 51410 30616 51416
rect 30576 51066 30604 51410
rect 30656 51400 30708 51406
rect 30656 51342 30708 51348
rect 30564 51060 30616 51066
rect 30564 51002 30616 51008
rect 30668 50862 30696 51342
rect 30656 50856 30708 50862
rect 30656 50798 30708 50804
rect 30472 49768 30524 49774
rect 30472 49710 30524 49716
rect 30484 48890 30512 49710
rect 30656 49224 30708 49230
rect 30656 49166 30708 49172
rect 30472 48884 30524 48890
rect 30472 48826 30524 48832
rect 30668 48822 30696 49166
rect 30656 48816 30708 48822
rect 30656 48758 30708 48764
rect 30668 47598 30696 48758
rect 30472 47592 30524 47598
rect 30472 47534 30524 47540
rect 30656 47592 30708 47598
rect 30656 47534 30708 47540
rect 30484 47190 30512 47534
rect 30472 47184 30524 47190
rect 30472 47126 30524 47132
rect 30484 46034 30512 47126
rect 30472 46028 30524 46034
rect 30472 45970 30524 45976
rect 30656 46028 30708 46034
rect 30656 45970 30708 45976
rect 30472 45348 30524 45354
rect 30472 45290 30524 45296
rect 30484 45082 30512 45290
rect 30472 45076 30524 45082
rect 30472 45018 30524 45024
rect 30668 44810 30696 45970
rect 30656 44804 30708 44810
rect 30656 44746 30708 44752
rect 30564 44328 30616 44334
rect 30564 44270 30616 44276
rect 30472 44192 30524 44198
rect 30472 44134 30524 44140
rect 30484 43858 30512 44134
rect 30472 43852 30524 43858
rect 30472 43794 30524 43800
rect 30576 43790 30604 44270
rect 30564 43784 30616 43790
rect 30564 43726 30616 43732
rect 30576 43382 30604 43726
rect 30564 43376 30616 43382
rect 30564 43318 30616 43324
rect 30564 43240 30616 43246
rect 30564 43182 30616 43188
rect 30472 42764 30524 42770
rect 30472 42706 30524 42712
rect 30484 42362 30512 42706
rect 30472 42356 30524 42362
rect 30472 42298 30524 42304
rect 30576 41274 30604 43182
rect 30668 42770 30696 44746
rect 30656 42764 30708 42770
rect 30656 42706 30708 42712
rect 30564 41268 30616 41274
rect 30564 41210 30616 41216
rect 30472 37324 30524 37330
rect 30472 37266 30524 37272
rect 30656 37324 30708 37330
rect 30656 37266 30708 37272
rect 30484 36922 30512 37266
rect 30564 37120 30616 37126
rect 30564 37062 30616 37068
rect 30472 36916 30524 36922
rect 30472 36858 30524 36864
rect 30576 36718 30604 37062
rect 30668 36854 30696 37266
rect 30656 36848 30708 36854
rect 30656 36790 30708 36796
rect 30564 36712 30616 36718
rect 30564 36654 30616 36660
rect 30576 36242 30604 36654
rect 30564 36236 30616 36242
rect 30564 36178 30616 36184
rect 30760 36122 30788 53042
rect 30852 51474 30880 53230
rect 30932 53236 30984 53242
rect 30932 53178 30984 53184
rect 31312 52970 31340 53654
rect 31300 52964 31352 52970
rect 31300 52906 31352 52912
rect 30840 51468 30892 51474
rect 30840 51410 30892 51416
rect 30852 46186 30880 51410
rect 31312 51074 31340 52906
rect 31496 52698 31524 54062
rect 32876 54058 32904 54674
rect 32864 54052 32916 54058
rect 32864 53994 32916 54000
rect 32968 53990 32996 54692
rect 33048 54674 33100 54680
rect 33244 54534 33272 55694
rect 33428 55282 33456 56170
rect 33796 55978 33824 57326
rect 33520 55950 33824 55978
rect 33520 55350 33548 55950
rect 34164 55826 34192 57990
rect 34244 57928 34296 57934
rect 34244 57870 34296 57876
rect 35084 57882 35112 59200
rect 34256 57254 34284 57870
rect 35084 57854 35296 57882
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 35268 57390 35296 57854
rect 35256 57384 35308 57390
rect 35256 57326 35308 57332
rect 34244 57248 34296 57254
rect 34244 57190 34296 57196
rect 34612 57248 34664 57254
rect 34612 57190 34664 57196
rect 34428 56840 34480 56846
rect 34428 56782 34480 56788
rect 34336 56772 34388 56778
rect 34336 56714 34388 56720
rect 34348 56488 34376 56714
rect 34440 56710 34468 56782
rect 34428 56704 34480 56710
rect 34428 56646 34480 56652
rect 34256 56460 34376 56488
rect 33692 55820 33744 55826
rect 33692 55762 33744 55768
rect 34152 55820 34204 55826
rect 34152 55762 34204 55768
rect 33508 55344 33560 55350
rect 33508 55286 33560 55292
rect 33416 55276 33468 55282
rect 33704 55264 33732 55762
rect 33876 55276 33928 55282
rect 33704 55236 33876 55264
rect 33416 55218 33468 55224
rect 33876 55218 33928 55224
rect 34060 55276 34112 55282
rect 34060 55218 34112 55224
rect 33508 55208 33560 55214
rect 33508 55150 33560 55156
rect 33416 55072 33468 55078
rect 33416 55014 33468 55020
rect 33232 54528 33284 54534
rect 33232 54470 33284 54476
rect 33048 54120 33100 54126
rect 33048 54062 33100 54068
rect 32956 53984 33008 53990
rect 32956 53926 33008 53932
rect 31760 53508 31812 53514
rect 31760 53450 31812 53456
rect 31772 53122 31800 53450
rect 32036 53440 32088 53446
rect 32036 53382 32088 53388
rect 32220 53440 32272 53446
rect 32220 53382 32272 53388
rect 31680 53094 31800 53122
rect 32048 53106 32076 53382
rect 31680 53038 31708 53094
rect 31668 53032 31720 53038
rect 31668 52974 31720 52980
rect 31484 52692 31536 52698
rect 31484 52634 31536 52640
rect 31772 51950 31800 53094
rect 32036 53100 32088 53106
rect 32036 53042 32088 53048
rect 31944 53032 31996 53038
rect 31942 53000 31944 53009
rect 31996 53000 31998 53009
rect 32232 52970 32260 53382
rect 33060 53174 33088 54062
rect 33140 54052 33192 54058
rect 33140 53994 33192 54000
rect 33048 53168 33100 53174
rect 33048 53110 33100 53116
rect 33060 53038 33088 53110
rect 33048 53032 33100 53038
rect 33048 52974 33100 52980
rect 33152 52970 33180 53994
rect 33244 53650 33272 54470
rect 33324 53984 33376 53990
rect 33324 53926 33376 53932
rect 33232 53644 33284 53650
rect 33232 53586 33284 53592
rect 31942 52935 31998 52944
rect 32220 52964 32272 52970
rect 31760 51944 31812 51950
rect 31760 51886 31812 51892
rect 31956 51406 31984 52935
rect 32220 52906 32272 52912
rect 33140 52964 33192 52970
rect 33140 52906 33192 52912
rect 32128 52896 32180 52902
rect 32128 52838 32180 52844
rect 32036 52556 32088 52562
rect 32036 52498 32088 52504
rect 32048 52154 32076 52498
rect 32036 52148 32088 52154
rect 32036 52090 32088 52096
rect 32140 52086 32168 52838
rect 32588 52556 32640 52562
rect 32588 52498 32640 52504
rect 32128 52080 32180 52086
rect 32128 52022 32180 52028
rect 32600 51882 32628 52498
rect 32588 51876 32640 51882
rect 32588 51818 32640 51824
rect 32600 51474 32628 51818
rect 33152 51610 33180 52906
rect 33244 52698 33272 53586
rect 33336 52902 33364 53926
rect 33324 52896 33376 52902
rect 33324 52838 33376 52844
rect 33232 52692 33284 52698
rect 33232 52634 33284 52640
rect 33428 51950 33456 55014
rect 33520 54058 33548 55150
rect 33692 54596 33744 54602
rect 33692 54538 33744 54544
rect 33704 54330 33732 54538
rect 33876 54528 33928 54534
rect 33876 54470 33928 54476
rect 33692 54324 33744 54330
rect 33692 54266 33744 54272
rect 33600 54120 33652 54126
rect 33600 54062 33652 54068
rect 33508 54052 33560 54058
rect 33508 53994 33560 54000
rect 33612 53786 33640 54062
rect 33784 53984 33836 53990
rect 33784 53926 33836 53932
rect 33600 53780 33652 53786
rect 33600 53722 33652 53728
rect 33508 53032 33560 53038
rect 33508 52974 33560 52980
rect 33520 52358 33548 52974
rect 33508 52352 33560 52358
rect 33508 52294 33560 52300
rect 33612 52018 33640 53722
rect 33796 53718 33824 53926
rect 33784 53712 33836 53718
rect 33784 53654 33836 53660
rect 33888 53446 33916 54470
rect 33876 53440 33928 53446
rect 33876 53382 33928 53388
rect 33784 52896 33836 52902
rect 33784 52838 33836 52844
rect 33796 52630 33824 52838
rect 33784 52624 33836 52630
rect 33784 52566 33836 52572
rect 34072 52562 34100 55218
rect 34256 55146 34284 56460
rect 34428 56432 34480 56438
rect 34428 56374 34480 56380
rect 34624 56386 34652 57190
rect 35622 57080 35678 57089
rect 35912 57050 35940 59200
rect 36268 57792 36320 57798
rect 36268 57734 36320 57740
rect 35622 57015 35678 57024
rect 35900 57044 35952 57050
rect 35440 56908 35492 56914
rect 35440 56850 35492 56856
rect 34716 56766 35296 56794
rect 34716 56506 34744 56766
rect 35268 56710 35296 56766
rect 34796 56704 34848 56710
rect 34796 56646 34848 56652
rect 35256 56704 35308 56710
rect 35256 56646 35308 56652
rect 34704 56500 34756 56506
rect 34704 56442 34756 56448
rect 34440 56302 34468 56374
rect 34624 56358 34744 56386
rect 34428 56296 34480 56302
rect 34428 56238 34480 56244
rect 34520 56228 34572 56234
rect 34520 56170 34572 56176
rect 34532 55350 34560 56170
rect 34520 55344 34572 55350
rect 34716 55298 34744 56358
rect 34808 56302 34836 56646
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 35256 56500 35308 56506
rect 35452 56488 35480 56850
rect 35308 56460 35480 56488
rect 35256 56442 35308 56448
rect 35636 56438 35664 57015
rect 35900 56986 35952 56992
rect 35898 56944 35954 56953
rect 35898 56879 35900 56888
rect 35952 56879 35954 56888
rect 35900 56850 35952 56856
rect 35624 56432 35676 56438
rect 34978 56400 35034 56409
rect 35624 56374 35676 56380
rect 34978 56335 35034 56344
rect 34796 56296 34848 56302
rect 34796 56238 34848 56244
rect 34808 55894 34836 56238
rect 34992 56166 35020 56335
rect 36280 56302 36308 57734
rect 36648 57458 36676 59200
rect 37096 57860 37148 57866
rect 37096 57802 37148 57808
rect 36636 57452 36688 57458
rect 36636 57394 36688 57400
rect 37108 57390 37136 57802
rect 36452 57384 36504 57390
rect 36452 57326 36504 57332
rect 37096 57384 37148 57390
rect 37096 57326 37148 57332
rect 36268 56296 36320 56302
rect 36082 56264 36138 56273
rect 36268 56238 36320 56244
rect 36082 56199 36138 56208
rect 36096 56166 36124 56199
rect 34980 56160 35032 56166
rect 34980 56102 35032 56108
rect 36084 56160 36136 56166
rect 36084 56102 36136 56108
rect 34796 55888 34848 55894
rect 36464 55865 36492 57326
rect 36912 57248 36964 57254
rect 36912 57190 36964 57196
rect 36924 56982 36952 57190
rect 36912 56976 36964 56982
rect 36912 56918 36964 56924
rect 37476 56914 37504 59200
rect 38212 57322 38240 59200
rect 39040 57458 39068 59200
rect 39028 57452 39080 57458
rect 39028 57394 39080 57400
rect 38200 57316 38252 57322
rect 38200 57258 38252 57264
rect 38936 57248 38988 57254
rect 38936 57190 38988 57196
rect 39580 57248 39632 57254
rect 39580 57190 39632 57196
rect 37464 56908 37516 56914
rect 37464 56850 37516 56856
rect 37648 56704 37700 56710
rect 37648 56646 37700 56652
rect 34796 55830 34848 55836
rect 36450 55856 36506 55865
rect 36450 55791 36506 55800
rect 34796 55616 34848 55622
rect 34796 55558 34848 55564
rect 34520 55286 34572 55292
rect 34624 55270 34744 55298
rect 34244 55140 34296 55146
rect 34244 55082 34296 55088
rect 34152 54732 34204 54738
rect 34152 54674 34204 54680
rect 34164 53242 34192 54674
rect 34624 53650 34652 55270
rect 34704 55208 34756 55214
rect 34808 55162 34836 55558
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 34756 55156 34836 55162
rect 34704 55150 34836 55156
rect 34716 55134 34836 55150
rect 34808 54670 34836 55134
rect 35256 55140 35308 55146
rect 35256 55082 35308 55088
rect 34796 54664 34848 54670
rect 34796 54606 34848 54612
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 35268 54330 35296 55082
rect 36176 55072 36228 55078
rect 36176 55014 36228 55020
rect 36188 54738 36216 55014
rect 37660 54806 37688 56646
rect 38948 56506 38976 57190
rect 38936 56500 38988 56506
rect 38936 56442 38988 56448
rect 37648 54800 37700 54806
rect 37648 54742 37700 54748
rect 36176 54732 36228 54738
rect 36176 54674 36228 54680
rect 35440 54596 35492 54602
rect 35440 54538 35492 54544
rect 35256 54324 35308 54330
rect 35256 54266 35308 54272
rect 35452 54126 35480 54538
rect 36188 54482 36216 54674
rect 36096 54454 36216 54482
rect 35900 54188 35952 54194
rect 35900 54130 35952 54136
rect 35440 54120 35492 54126
rect 35440 54062 35492 54068
rect 35912 53650 35940 54130
rect 36096 54058 36124 54454
rect 39592 54262 39620 57190
rect 39776 56914 39804 59200
rect 40604 57390 40632 59200
rect 41432 57458 41460 59200
rect 41420 57452 41472 57458
rect 41420 57394 41472 57400
rect 40592 57384 40644 57390
rect 40592 57326 40644 57332
rect 40408 57248 40460 57254
rect 40408 57190 40460 57196
rect 39764 56908 39816 56914
rect 39764 56850 39816 56856
rect 39580 54256 39632 54262
rect 39580 54198 39632 54204
rect 36176 54120 36228 54126
rect 36176 54062 36228 54068
rect 36360 54120 36412 54126
rect 36360 54062 36412 54068
rect 36084 54052 36136 54058
rect 36084 53994 36136 54000
rect 36188 53650 36216 54062
rect 36372 53990 36400 54062
rect 36360 53984 36412 53990
rect 36360 53926 36412 53932
rect 34612 53644 34664 53650
rect 34612 53586 34664 53592
rect 35900 53644 35952 53650
rect 35900 53586 35952 53592
rect 36176 53644 36228 53650
rect 36176 53586 36228 53592
rect 35716 53440 35768 53446
rect 35716 53382 35768 53388
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34152 53236 34204 53242
rect 34152 53178 34204 53184
rect 35728 53038 35756 53382
rect 36188 53242 36216 53586
rect 36372 53446 36400 53926
rect 36360 53440 36412 53446
rect 36360 53382 36412 53388
rect 36728 53440 36780 53446
rect 36728 53382 36780 53388
rect 36176 53236 36228 53242
rect 36176 53178 36228 53184
rect 34704 53032 34756 53038
rect 34702 53000 34704 53009
rect 35716 53032 35768 53038
rect 34756 53000 34758 53009
rect 35716 52974 35768 52980
rect 34702 52935 34758 52944
rect 36740 52698 36768 53382
rect 40420 53174 40448 57190
rect 42168 56914 42196 59200
rect 42996 57390 43024 59200
rect 43732 57390 43760 59200
rect 44560 57390 44588 59200
rect 45388 57458 45416 59200
rect 45376 57452 45428 57458
rect 45376 57394 45428 57400
rect 46124 57390 46152 59200
rect 46952 57526 46980 59200
rect 46940 57520 46992 57526
rect 46940 57462 46992 57468
rect 47688 57390 47716 59200
rect 48516 57390 48544 59200
rect 49252 57458 49280 59200
rect 50080 57458 50108 59200
rect 49240 57452 49292 57458
rect 49240 57394 49292 57400
rect 50068 57452 50120 57458
rect 50908 57440 50936 59200
rect 50908 57412 51120 57440
rect 50068 57394 50120 57400
rect 42984 57384 43036 57390
rect 42984 57326 43036 57332
rect 43720 57384 43772 57390
rect 43720 57326 43772 57332
rect 44548 57384 44600 57390
rect 44548 57326 44600 57332
rect 46112 57384 46164 57390
rect 46112 57326 46164 57332
rect 47676 57384 47728 57390
rect 47676 57326 47728 57332
rect 48504 57384 48556 57390
rect 48504 57326 48556 57332
rect 50300 57148 50596 57168
rect 50356 57146 50380 57148
rect 50436 57146 50460 57148
rect 50516 57146 50540 57148
rect 50378 57094 50380 57146
rect 50442 57094 50454 57146
rect 50516 57094 50518 57146
rect 50356 57092 50380 57094
rect 50436 57092 50460 57094
rect 50516 57092 50540 57094
rect 50300 57072 50596 57092
rect 51092 56914 51120 57412
rect 51644 56914 51672 59200
rect 42156 56908 42208 56914
rect 42156 56850 42208 56856
rect 51080 56908 51132 56914
rect 51080 56850 51132 56856
rect 51632 56908 51684 56914
rect 51632 56850 51684 56856
rect 52472 56302 52500 59200
rect 53104 57316 53156 57322
rect 53104 57258 53156 57264
rect 53116 57050 53144 57258
rect 53104 57044 53156 57050
rect 53104 56986 53156 56992
rect 52460 56296 52512 56302
rect 52460 56238 52512 56244
rect 50300 56060 50596 56080
rect 50356 56058 50380 56060
rect 50436 56058 50460 56060
rect 50516 56058 50540 56060
rect 50378 56006 50380 56058
rect 50442 56006 50454 56058
rect 50516 56006 50518 56058
rect 50356 56004 50380 56006
rect 50436 56004 50460 56006
rect 50516 56004 50540 56006
rect 50300 55984 50596 56004
rect 53208 55826 53236 59200
rect 53748 58064 53800 58070
rect 53748 58006 53800 58012
rect 53760 57390 53788 58006
rect 53748 57384 53800 57390
rect 53748 57326 53800 57332
rect 53932 56432 53984 56438
rect 53932 56374 53984 56380
rect 53196 55820 53248 55826
rect 53196 55762 53248 55768
rect 53944 55214 53972 56374
rect 54036 55826 54064 59200
rect 54116 57384 54168 57390
rect 54116 57326 54168 57332
rect 54128 56914 54156 57326
rect 54772 56930 54800 59200
rect 55312 58676 55364 58682
rect 55312 58618 55364 58624
rect 55126 58304 55182 58313
rect 55126 58239 55182 58248
rect 55140 57526 55168 58239
rect 55128 57520 55180 57526
rect 55128 57462 55180 57468
rect 54116 56908 54168 56914
rect 54116 56850 54168 56856
rect 54680 56902 54800 56930
rect 54576 56840 54628 56846
rect 54576 56782 54628 56788
rect 54300 56296 54352 56302
rect 54300 56238 54352 56244
rect 54024 55820 54076 55826
rect 54024 55762 54076 55768
rect 53932 55208 53984 55214
rect 53932 55150 53984 55156
rect 50300 54972 50596 54992
rect 50356 54970 50380 54972
rect 50436 54970 50460 54972
rect 50516 54970 50540 54972
rect 50378 54918 50380 54970
rect 50442 54918 50454 54970
rect 50516 54918 50518 54970
rect 50356 54916 50380 54918
rect 50436 54916 50460 54918
rect 50516 54916 50540 54918
rect 50300 54896 50596 54916
rect 50300 53884 50596 53904
rect 50356 53882 50380 53884
rect 50436 53882 50460 53884
rect 50516 53882 50540 53884
rect 50378 53830 50380 53882
rect 50442 53830 50454 53882
rect 50516 53830 50518 53882
rect 50356 53828 50380 53830
rect 50436 53828 50460 53830
rect 50516 53828 50540 53830
rect 50300 53808 50596 53828
rect 40408 53168 40460 53174
rect 40408 53110 40460 53116
rect 50300 52796 50596 52816
rect 50356 52794 50380 52796
rect 50436 52794 50460 52796
rect 50516 52794 50540 52796
rect 50378 52742 50380 52794
rect 50442 52742 50454 52794
rect 50516 52742 50518 52794
rect 50356 52740 50380 52742
rect 50436 52740 50460 52742
rect 50516 52740 50540 52742
rect 50300 52720 50596 52740
rect 36728 52692 36780 52698
rect 36728 52634 36780 52640
rect 34060 52556 34112 52562
rect 34060 52498 34112 52504
rect 34336 52556 34388 52562
rect 34336 52498 34388 52504
rect 36268 52556 36320 52562
rect 36268 52498 36320 52504
rect 33600 52012 33652 52018
rect 33600 51954 33652 51960
rect 34348 51950 34376 52498
rect 36084 52488 36136 52494
rect 36084 52430 36136 52436
rect 35716 52352 35768 52358
rect 35716 52294 35768 52300
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 35728 51950 35756 52294
rect 33416 51944 33468 51950
rect 33416 51886 33468 51892
rect 34336 51944 34388 51950
rect 34336 51886 34388 51892
rect 35716 51944 35768 51950
rect 35716 51886 35768 51892
rect 33508 51808 33560 51814
rect 33508 51750 33560 51756
rect 33520 51610 33548 51750
rect 33140 51604 33192 51610
rect 33140 51546 33192 51552
rect 33508 51604 33560 51610
rect 33508 51546 33560 51552
rect 32312 51468 32364 51474
rect 32312 51410 32364 51416
rect 32588 51468 32640 51474
rect 32588 51410 32640 51416
rect 31944 51400 31996 51406
rect 31944 51342 31996 51348
rect 31220 51046 31340 51074
rect 31116 49836 31168 49842
rect 31116 49778 31168 49784
rect 30932 49700 30984 49706
rect 30932 49642 30984 49648
rect 30944 48890 30972 49642
rect 30932 48884 30984 48890
rect 30932 48826 30984 48832
rect 30944 48278 30972 48826
rect 31128 48686 31156 49778
rect 31116 48680 31168 48686
rect 31116 48622 31168 48628
rect 30932 48272 30984 48278
rect 30932 48214 30984 48220
rect 31220 48226 31248 51046
rect 31484 50924 31536 50930
rect 31484 50866 31536 50872
rect 31392 50720 31444 50726
rect 31392 50662 31444 50668
rect 31404 50454 31432 50662
rect 31392 50448 31444 50454
rect 31392 50390 31444 50396
rect 31496 50318 31524 50866
rect 31852 50856 31904 50862
rect 31852 50798 31904 50804
rect 31864 50522 31892 50798
rect 31852 50516 31904 50522
rect 31852 50458 31904 50464
rect 31956 50386 31984 51342
rect 32324 50522 32352 51410
rect 33232 50856 33284 50862
rect 33232 50798 33284 50804
rect 32956 50788 33008 50794
rect 32956 50730 33008 50736
rect 32312 50516 32364 50522
rect 32312 50458 32364 50464
rect 32968 50386 32996 50730
rect 33244 50522 33272 50798
rect 33232 50516 33284 50522
rect 33232 50458 33284 50464
rect 33520 50454 33548 51546
rect 34152 50720 34204 50726
rect 34152 50662 34204 50668
rect 34164 50454 34192 50662
rect 33508 50448 33560 50454
rect 33508 50390 33560 50396
rect 34152 50448 34204 50454
rect 34152 50390 34204 50396
rect 31944 50380 31996 50386
rect 31944 50322 31996 50328
rect 32496 50380 32548 50386
rect 32496 50322 32548 50328
rect 32956 50380 33008 50386
rect 32956 50322 33008 50328
rect 31484 50312 31536 50318
rect 31484 50254 31536 50260
rect 31496 49978 31524 50254
rect 31956 50250 31984 50322
rect 31944 50244 31996 50250
rect 31944 50186 31996 50192
rect 31484 49972 31536 49978
rect 31484 49914 31536 49920
rect 31484 49768 31536 49774
rect 31484 49710 31536 49716
rect 31668 49768 31720 49774
rect 31668 49710 31720 49716
rect 31300 49292 31352 49298
rect 31300 49234 31352 49240
rect 31312 48346 31340 49234
rect 31300 48340 31352 48346
rect 31300 48282 31352 48288
rect 31220 48198 31340 48226
rect 31496 48210 31524 49710
rect 31680 48890 31708 49710
rect 31760 49700 31812 49706
rect 31760 49642 31812 49648
rect 31772 49094 31800 49642
rect 31760 49088 31812 49094
rect 31760 49030 31812 49036
rect 31668 48884 31720 48890
rect 31668 48826 31720 48832
rect 31680 48210 31708 48826
rect 31772 48210 31800 49030
rect 31024 47524 31076 47530
rect 31024 47466 31076 47472
rect 31036 47258 31064 47466
rect 31024 47252 31076 47258
rect 31024 47194 31076 47200
rect 31208 46436 31260 46442
rect 31208 46378 31260 46384
rect 30852 46158 31064 46186
rect 31220 46170 31248 46378
rect 30840 42560 30892 42566
rect 30840 42502 30892 42508
rect 30852 41070 30880 42502
rect 30932 42288 30984 42294
rect 30932 42230 30984 42236
rect 30840 41064 30892 41070
rect 30840 41006 30892 41012
rect 30944 39914 30972 42230
rect 30932 39908 30984 39914
rect 30932 39850 30984 39856
rect 30944 38894 30972 39850
rect 30932 38888 30984 38894
rect 30932 38830 30984 38836
rect 30944 38418 30972 38830
rect 30932 38412 30984 38418
rect 30932 38354 30984 38360
rect 30944 37330 30972 38354
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30944 36786 30972 37266
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30576 36094 30788 36122
rect 30472 35080 30524 35086
rect 30472 35022 30524 35028
rect 30484 33998 30512 35022
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30484 32434 30512 33934
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30484 31890 30512 32370
rect 30472 31884 30524 31890
rect 30472 31826 30524 31832
rect 30472 30184 30524 30190
rect 30470 30152 30472 30161
rect 30524 30152 30526 30161
rect 30470 30087 30526 30096
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 28724 29096 28776 29102
rect 28724 29038 28776 29044
rect 28828 28994 28856 29242
rect 30392 29102 30420 29582
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 28552 28966 28856 28994
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 28356 28960 28408 28966
rect 28356 28902 28408 28908
rect 28552 28558 28580 28966
rect 29012 28762 29040 28970
rect 30392 28762 30420 29038
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 29000 28620 29052 28626
rect 29000 28562 29052 28568
rect 28540 28552 28592 28558
rect 28540 28494 28592 28500
rect 28080 28144 28132 28150
rect 28080 28086 28132 28092
rect 28092 28014 28120 28086
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 28000 27606 28028 27882
rect 27988 27600 28040 27606
rect 27988 27542 28040 27548
rect 28000 26926 28028 27542
rect 29012 27010 29040 28562
rect 30286 28112 30342 28121
rect 30286 28047 30342 28056
rect 30300 27878 30328 28047
rect 30392 28014 30420 28698
rect 30380 28008 30432 28014
rect 30484 27985 30512 30087
rect 30380 27950 30432 27956
rect 30470 27976 30526 27985
rect 30470 27911 30526 27920
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 29104 27674 29132 27814
rect 29092 27668 29144 27674
rect 29092 27610 29144 27616
rect 30392 27606 30420 27814
rect 30380 27600 30432 27606
rect 30380 27542 30432 27548
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29012 26982 29132 27010
rect 27988 26920 28040 26926
rect 27988 26862 28040 26868
rect 29000 26920 29052 26926
rect 29104 26897 29132 26982
rect 29000 26862 29052 26868
rect 29090 26888 29146 26897
rect 28540 26784 28592 26790
rect 28540 26726 28592 26732
rect 28264 26444 28316 26450
rect 28264 26386 28316 26392
rect 27804 26308 27856 26314
rect 27804 26250 27856 26256
rect 28276 25838 28304 26386
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28276 25498 28304 25774
rect 28264 25492 28316 25498
rect 28264 25434 28316 25440
rect 27988 25356 28040 25362
rect 27988 25298 28040 25304
rect 28000 25158 28028 25298
rect 27988 25152 28040 25158
rect 27988 25094 28040 25100
rect 27804 24812 27856 24818
rect 27804 24754 27856 24760
rect 27816 24721 27844 24754
rect 27802 24712 27858 24721
rect 27802 24647 27858 24656
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 26516 23180 26568 23186
rect 26516 23122 26568 23128
rect 26884 22976 26936 22982
rect 26422 22944 26478 22953
rect 26422 22879 26478 22888
rect 26804 22936 26884 22964
rect 26436 22642 26464 22879
rect 26424 22636 26476 22642
rect 26424 22578 26476 22584
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26608 21344 26660 21350
rect 26608 21286 26660 21292
rect 26620 21010 26648 21286
rect 26516 21004 26568 21010
rect 26516 20946 26568 20952
rect 26608 21004 26660 21010
rect 26608 20946 26660 20952
rect 26528 20602 26556 20946
rect 26712 20913 26740 21490
rect 26804 21486 26832 22936
rect 26884 22918 26936 22924
rect 27066 22536 27122 22545
rect 27066 22471 27122 22480
rect 27080 21486 27108 22471
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 27068 21480 27120 21486
rect 27068 21422 27120 21428
rect 26698 20904 26754 20913
rect 26698 20839 26754 20848
rect 26712 20806 26740 20839
rect 26700 20800 26752 20806
rect 26700 20742 26752 20748
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26424 20324 26476 20330
rect 26424 20266 26476 20272
rect 26436 18630 26464 20266
rect 26608 19984 26660 19990
rect 26608 19926 26660 19932
rect 26620 19310 26648 19926
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26712 19310 26740 19858
rect 26608 19304 26660 19310
rect 26608 19246 26660 19252
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 26528 18766 26556 19110
rect 26608 18828 26660 18834
rect 26712 18816 26740 19246
rect 26660 18788 26740 18816
rect 26608 18770 26660 18776
rect 26516 18760 26568 18766
rect 26516 18702 26568 18708
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 25780 18148 25832 18154
rect 25780 18090 25832 18096
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25780 17672 25832 17678
rect 25780 17614 25832 17620
rect 25792 17338 25820 17614
rect 24768 17332 24820 17338
rect 24768 17274 24820 17280
rect 25780 17332 25832 17338
rect 25780 17274 25832 17280
rect 26068 16658 26096 18158
rect 26160 17542 26188 18226
rect 26620 17882 26648 18770
rect 26804 18222 26832 21422
rect 26976 21412 27028 21418
rect 26976 21354 27028 21360
rect 26884 21344 26936 21350
rect 26884 21286 26936 21292
rect 26896 20942 26924 21286
rect 26988 21049 27016 21354
rect 26974 21040 27030 21049
rect 26974 20975 27030 20984
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 26884 20256 26936 20262
rect 26884 20198 26936 20204
rect 26896 18222 26924 20198
rect 26976 19916 27028 19922
rect 26976 19858 27028 19864
rect 26988 19378 27016 19858
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27080 19514 27108 19790
rect 27068 19508 27120 19514
rect 27068 19450 27120 19456
rect 27172 19378 27200 23462
rect 27356 23050 27384 24210
rect 27816 23730 27844 24647
rect 28000 24614 28028 25094
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27344 23044 27396 23050
rect 27344 22986 27396 22992
rect 27356 22574 27384 22986
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27894 22536 27950 22545
rect 27894 22471 27950 22480
rect 27908 22438 27936 22471
rect 27620 22432 27672 22438
rect 27620 22374 27672 22380
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27632 21962 27660 22374
rect 27908 22166 27936 22374
rect 27896 22160 27948 22166
rect 28000 22137 28028 24550
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 28264 22976 28316 22982
rect 28264 22918 28316 22924
rect 27896 22102 27948 22108
rect 27986 22128 28042 22137
rect 27986 22063 28042 22072
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27620 21956 27672 21962
rect 27620 21898 27672 21904
rect 27342 21856 27398 21865
rect 27342 21791 27398 21800
rect 27356 21690 27384 21791
rect 27252 21684 27304 21690
rect 27252 21626 27304 21632
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27264 21350 27292 21626
rect 27632 21486 27660 21898
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27632 21010 27660 21422
rect 27620 21004 27672 21010
rect 27620 20946 27672 20952
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27724 19990 27752 20470
rect 27816 20466 27844 21966
rect 27804 20460 27856 20466
rect 27804 20402 27856 20408
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 28276 19922 28304 22918
rect 28368 19990 28396 24142
rect 28448 24064 28500 24070
rect 28448 24006 28500 24012
rect 28460 23662 28488 24006
rect 28448 23656 28500 23662
rect 28448 23598 28500 23604
rect 28552 22574 28580 26726
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28630 22672 28686 22681
rect 28630 22607 28686 22616
rect 28644 22574 28672 22607
rect 28540 22568 28592 22574
rect 28540 22510 28592 22516
rect 28632 22568 28684 22574
rect 28632 22510 28684 22516
rect 28540 21480 28592 21486
rect 28540 21422 28592 21428
rect 28552 20874 28580 21422
rect 28540 20868 28592 20874
rect 28540 20810 28592 20816
rect 28356 19984 28408 19990
rect 28356 19926 28408 19932
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 28264 19916 28316 19922
rect 28264 19858 28316 19864
rect 27632 19446 27660 19858
rect 27896 19848 27948 19854
rect 27896 19790 27948 19796
rect 27620 19440 27672 19446
rect 27620 19382 27672 19388
rect 26976 19372 27028 19378
rect 26976 19314 27028 19320
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 26988 19242 27016 19314
rect 26976 19236 27028 19242
rect 26976 19178 27028 19184
rect 26988 18834 27016 19178
rect 27908 19174 27936 19790
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28368 18426 28396 18770
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28552 18290 28580 20810
rect 28644 19922 28672 22510
rect 28736 22250 28764 25230
rect 29012 24290 29040 26862
rect 29090 26823 29146 26832
rect 29104 24342 29132 26823
rect 29184 26240 29236 26246
rect 29184 26182 29236 26188
rect 29196 25344 29224 26182
rect 29380 26042 29408 27066
rect 30024 26926 30052 27270
rect 30208 26926 30236 27474
rect 30392 26926 30420 27542
rect 29460 26920 29512 26926
rect 29460 26862 29512 26868
rect 30012 26920 30064 26926
rect 30012 26862 30064 26868
rect 30196 26920 30248 26926
rect 30196 26862 30248 26868
rect 30380 26920 30432 26926
rect 30380 26862 30432 26868
rect 29368 26036 29420 26042
rect 29368 25978 29420 25984
rect 29276 25356 29328 25362
rect 29196 25316 29276 25344
rect 28828 24262 29040 24290
rect 29092 24336 29144 24342
rect 29092 24278 29144 24284
rect 28828 23225 28856 24262
rect 28908 24200 28960 24206
rect 28908 24142 28960 24148
rect 28814 23216 28870 23225
rect 28814 23151 28816 23160
rect 28868 23151 28870 23160
rect 28816 23122 28868 23128
rect 28920 22778 28948 24142
rect 28908 22772 28960 22778
rect 28908 22714 28960 22720
rect 29000 22772 29052 22778
rect 29000 22714 29052 22720
rect 29012 22574 29040 22714
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 28736 22222 28948 22250
rect 28722 22128 28778 22137
rect 28722 22063 28778 22072
rect 28736 21010 28764 22063
rect 28814 21312 28870 21321
rect 28814 21247 28870 21256
rect 28724 21004 28776 21010
rect 28724 20946 28776 20952
rect 28724 19984 28776 19990
rect 28724 19926 28776 19932
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28736 19514 28764 19926
rect 28828 19922 28856 21247
rect 28920 21078 28948 22222
rect 29012 21690 29040 22510
rect 29196 22420 29224 25316
rect 29276 25298 29328 25304
rect 29368 25152 29420 25158
rect 29368 25094 29420 25100
rect 29380 24750 29408 25094
rect 29368 24744 29420 24750
rect 29368 24686 29420 24692
rect 29368 23860 29420 23866
rect 29368 23802 29420 23808
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29288 22574 29316 23054
rect 29276 22568 29328 22574
rect 29276 22510 29328 22516
rect 29380 22506 29408 23802
rect 29472 23186 29500 26862
rect 29552 26444 29604 26450
rect 29552 26386 29604 26392
rect 29564 24410 29592 26386
rect 29644 25764 29696 25770
rect 29644 25706 29696 25712
rect 29552 24404 29604 24410
rect 29552 24346 29604 24352
rect 29460 23180 29512 23186
rect 29460 23122 29512 23128
rect 29472 23089 29500 23122
rect 29458 23080 29514 23089
rect 29458 23015 29514 23024
rect 29552 23044 29604 23050
rect 29552 22986 29604 22992
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29368 22500 29420 22506
rect 29368 22442 29420 22448
rect 29196 22392 29316 22420
rect 29184 22092 29236 22098
rect 29184 22034 29236 22040
rect 29092 21888 29144 21894
rect 29092 21830 29144 21836
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 29104 21486 29132 21830
rect 29092 21480 29144 21486
rect 29092 21422 29144 21428
rect 29000 21412 29052 21418
rect 29000 21354 29052 21360
rect 28908 21072 28960 21078
rect 28908 21014 28960 21020
rect 29012 20874 29040 21354
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 29012 20602 29040 20810
rect 29000 20596 29052 20602
rect 29000 20538 29052 20544
rect 28816 19916 28868 19922
rect 28816 19858 28868 19864
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 29104 19310 29132 21286
rect 28908 19304 28960 19310
rect 28722 19272 28778 19281
rect 28908 19246 28960 19252
rect 29092 19304 29144 19310
rect 29092 19246 29144 19252
rect 28722 19207 28778 19216
rect 28632 19168 28684 19174
rect 28632 19110 28684 19116
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 28644 18222 28672 19110
rect 28736 18766 28764 19207
rect 28920 18970 28948 19246
rect 29196 18970 29224 22034
rect 29288 21010 29316 22392
rect 29472 21894 29500 22510
rect 29460 21888 29512 21894
rect 29460 21830 29512 21836
rect 29276 21004 29328 21010
rect 29276 20946 29328 20952
rect 29276 20324 29328 20330
rect 29276 20266 29328 20272
rect 28908 18964 28960 18970
rect 28908 18906 28960 18912
rect 29184 18964 29236 18970
rect 29184 18906 29236 18912
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 29288 18426 29316 20266
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29380 18834 29408 20198
rect 29564 19310 29592 22986
rect 29656 20262 29684 25706
rect 29828 25696 29880 25702
rect 29828 25638 29880 25644
rect 29736 24744 29788 24750
rect 29736 24686 29788 24692
rect 29748 23866 29776 24686
rect 29736 23860 29788 23866
rect 29736 23802 29788 23808
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29748 20398 29776 20742
rect 29736 20392 29788 20398
rect 29736 20334 29788 20340
rect 29644 20256 29696 20262
rect 29644 20198 29696 20204
rect 29840 19310 29868 25638
rect 29920 25424 29972 25430
rect 29920 25366 29972 25372
rect 29932 19514 29960 25366
rect 30024 23594 30052 26862
rect 30208 26042 30236 26862
rect 30288 26852 30340 26858
rect 30288 26794 30340 26800
rect 30300 26586 30328 26794
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30300 25838 30328 26522
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30484 25702 30512 27911
rect 30576 26518 30604 36094
rect 30748 35488 30800 35494
rect 30748 35430 30800 35436
rect 30760 35222 30788 35430
rect 30748 35216 30800 35222
rect 30748 35158 30800 35164
rect 31036 34626 31064 46158
rect 31208 46164 31260 46170
rect 31208 46106 31260 46112
rect 31220 45626 31248 46106
rect 31208 45620 31260 45626
rect 31208 45562 31260 45568
rect 31116 42560 31168 42566
rect 31116 42502 31168 42508
rect 31128 42090 31156 42502
rect 31116 42084 31168 42090
rect 31116 42026 31168 42032
rect 31312 41414 31340 48198
rect 31484 48204 31536 48210
rect 31484 48146 31536 48152
rect 31668 48204 31720 48210
rect 31668 48146 31720 48152
rect 31760 48204 31812 48210
rect 31760 48146 31812 48152
rect 31852 48136 31904 48142
rect 31852 48078 31904 48084
rect 31760 48000 31812 48006
rect 31760 47942 31812 47948
rect 31772 46578 31800 47942
rect 31864 47054 31892 48078
rect 31956 48006 31984 50186
rect 32508 49978 32536 50322
rect 32496 49972 32548 49978
rect 32496 49914 32548 49920
rect 33140 49836 33192 49842
rect 33060 49796 33140 49824
rect 33060 48210 33088 49796
rect 33140 49778 33192 49784
rect 33520 49774 33548 50390
rect 34348 49978 34376 51886
rect 36096 51882 36124 52430
rect 36176 52352 36228 52358
rect 36176 52294 36228 52300
rect 36188 51950 36216 52294
rect 36280 52154 36308 52498
rect 36268 52148 36320 52154
rect 36268 52090 36320 52096
rect 36176 51944 36228 51950
rect 36176 51886 36228 51892
rect 36084 51876 36136 51882
rect 36084 51818 36136 51824
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 36188 51066 36216 51886
rect 50300 51708 50596 51728
rect 50356 51706 50380 51708
rect 50436 51706 50460 51708
rect 50516 51706 50540 51708
rect 50378 51654 50380 51706
rect 50442 51654 50454 51706
rect 50516 51654 50518 51706
rect 50356 51652 50380 51654
rect 50436 51652 50460 51654
rect 50516 51652 50540 51654
rect 50300 51632 50596 51652
rect 36176 51060 36228 51066
rect 36176 51002 36228 51008
rect 34796 50924 34848 50930
rect 34796 50866 34848 50872
rect 34704 50856 34756 50862
rect 34704 50798 34756 50804
rect 34336 49972 34388 49978
rect 34336 49914 34388 49920
rect 33508 49768 33560 49774
rect 33508 49710 33560 49716
rect 34244 49768 34296 49774
rect 34244 49710 34296 49716
rect 33692 49224 33744 49230
rect 33692 49166 33744 49172
rect 33324 49088 33376 49094
rect 33324 49030 33376 49036
rect 33336 48686 33364 49030
rect 33324 48680 33376 48686
rect 33324 48622 33376 48628
rect 33704 48346 33732 49166
rect 33692 48340 33744 48346
rect 33692 48282 33744 48288
rect 32220 48204 32272 48210
rect 32220 48146 32272 48152
rect 33048 48204 33100 48210
rect 33048 48146 33100 48152
rect 33692 48204 33744 48210
rect 33692 48146 33744 48152
rect 31944 48000 31996 48006
rect 31944 47942 31996 47948
rect 32232 47802 32260 48146
rect 32220 47796 32272 47802
rect 32220 47738 32272 47744
rect 32036 47456 32088 47462
rect 32036 47398 32088 47404
rect 32048 47122 32076 47398
rect 32036 47116 32088 47122
rect 32036 47058 32088 47064
rect 31852 47048 31904 47054
rect 31852 46990 31904 46996
rect 31864 46714 31892 46990
rect 31944 46980 31996 46986
rect 31944 46922 31996 46928
rect 31852 46708 31904 46714
rect 31852 46650 31904 46656
rect 31760 46572 31812 46578
rect 31760 46514 31812 46520
rect 31956 46510 31984 46922
rect 32048 46510 32076 47058
rect 32312 47048 32364 47054
rect 32312 46990 32364 46996
rect 32324 46578 32352 46990
rect 32404 46640 32456 46646
rect 32404 46582 32456 46588
rect 32312 46572 32364 46578
rect 32312 46514 32364 46520
rect 31484 46504 31536 46510
rect 31484 46446 31536 46452
rect 31944 46504 31996 46510
rect 31944 46446 31996 46452
rect 32036 46504 32088 46510
rect 32036 46446 32088 46452
rect 31392 46368 31444 46374
rect 31392 46310 31444 46316
rect 31404 45354 31432 46310
rect 31496 45354 31524 46446
rect 31956 45558 31984 46446
rect 31944 45552 31996 45558
rect 31944 45494 31996 45500
rect 32416 45422 32444 46582
rect 33060 46102 33088 48146
rect 33508 47592 33560 47598
rect 33508 47534 33560 47540
rect 33140 47456 33192 47462
rect 33140 47398 33192 47404
rect 33152 47190 33180 47398
rect 33520 47258 33548 47534
rect 33704 47530 33732 48146
rect 34256 48074 34284 49710
rect 34348 48754 34376 49914
rect 34716 49774 34744 50798
rect 34808 50522 34836 50866
rect 50300 50620 50596 50640
rect 50356 50618 50380 50620
rect 50436 50618 50460 50620
rect 50516 50618 50540 50620
rect 50378 50566 50380 50618
rect 50442 50566 50454 50618
rect 50516 50566 50518 50618
rect 50356 50564 50380 50566
rect 50436 50564 50460 50566
rect 50516 50564 50540 50566
rect 50300 50544 50596 50564
rect 34796 50516 34848 50522
rect 34796 50458 34848 50464
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34704 49768 34756 49774
rect 34756 49728 34836 49756
rect 34704 49710 34756 49716
rect 34612 49632 34664 49638
rect 34612 49574 34664 49580
rect 34428 49360 34480 49366
rect 34428 49302 34480 49308
rect 34440 48890 34468 49302
rect 34428 48884 34480 48890
rect 34428 48826 34480 48832
rect 34336 48748 34388 48754
rect 34336 48690 34388 48696
rect 34440 48346 34468 48826
rect 34624 48618 34652 49574
rect 34808 49434 34836 49728
rect 50300 49532 50596 49552
rect 50356 49530 50380 49532
rect 50436 49530 50460 49532
rect 50516 49530 50540 49532
rect 50378 49478 50380 49530
rect 50442 49478 50454 49530
rect 50516 49478 50518 49530
rect 50356 49476 50380 49478
rect 50436 49476 50460 49478
rect 50516 49476 50540 49478
rect 50300 49456 50596 49476
rect 34796 49428 34848 49434
rect 34796 49370 34848 49376
rect 35256 49360 35308 49366
rect 35256 49302 35308 49308
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 35268 48890 35296 49302
rect 35256 48884 35308 48890
rect 35256 48826 35308 48832
rect 34612 48612 34664 48618
rect 34612 48554 34664 48560
rect 34428 48340 34480 48346
rect 34428 48282 34480 48288
rect 35268 48278 35296 48826
rect 50300 48444 50596 48464
rect 50356 48442 50380 48444
rect 50436 48442 50460 48444
rect 50516 48442 50540 48444
rect 50378 48390 50380 48442
rect 50442 48390 50454 48442
rect 50516 48390 50518 48442
rect 50356 48388 50380 48390
rect 50436 48388 50460 48390
rect 50516 48388 50540 48390
rect 50300 48368 50596 48388
rect 35256 48272 35308 48278
rect 35256 48214 35308 48220
rect 34244 48068 34296 48074
rect 34244 48010 34296 48016
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 34336 47592 34388 47598
rect 34336 47534 34388 47540
rect 33692 47524 33744 47530
rect 33692 47466 33744 47472
rect 34244 47524 34296 47530
rect 34244 47466 34296 47472
rect 34256 47258 34284 47466
rect 33508 47252 33560 47258
rect 33508 47194 33560 47200
rect 34244 47252 34296 47258
rect 34244 47194 34296 47200
rect 33140 47184 33192 47190
rect 33140 47126 33192 47132
rect 34348 47122 34376 47534
rect 50300 47356 50596 47376
rect 50356 47354 50380 47356
rect 50436 47354 50460 47356
rect 50516 47354 50540 47356
rect 50378 47302 50380 47354
rect 50442 47302 50454 47354
rect 50516 47302 50518 47354
rect 50356 47300 50380 47302
rect 50436 47300 50460 47302
rect 50516 47300 50540 47302
rect 50300 47280 50596 47300
rect 34336 47116 34388 47122
rect 34336 47058 34388 47064
rect 33508 46436 33560 46442
rect 33508 46378 33560 46384
rect 33416 46368 33468 46374
rect 33416 46310 33468 46316
rect 33048 46096 33100 46102
rect 33048 46038 33100 46044
rect 33428 46034 33456 46310
rect 33520 46170 33548 46378
rect 34348 46374 34376 47058
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34336 46368 34388 46374
rect 34336 46310 34388 46316
rect 50300 46268 50596 46288
rect 50356 46266 50380 46268
rect 50436 46266 50460 46268
rect 50516 46266 50540 46268
rect 50378 46214 50380 46266
rect 50442 46214 50454 46266
rect 50516 46214 50518 46266
rect 50356 46212 50380 46214
rect 50436 46212 50460 46214
rect 50516 46212 50540 46214
rect 50300 46192 50596 46212
rect 33508 46164 33560 46170
rect 33508 46106 33560 46112
rect 32956 46028 33008 46034
rect 32956 45970 33008 45976
rect 33416 46028 33468 46034
rect 33416 45970 33468 45976
rect 32968 45490 32996 45970
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 32956 45484 33008 45490
rect 32956 45426 33008 45432
rect 32404 45416 32456 45422
rect 32404 45358 32456 45364
rect 31392 45348 31444 45354
rect 31392 45290 31444 45296
rect 31484 45348 31536 45354
rect 31484 45290 31536 45296
rect 31404 44946 31432 45290
rect 31496 45082 31524 45290
rect 50300 45180 50596 45200
rect 50356 45178 50380 45180
rect 50436 45178 50460 45180
rect 50516 45178 50540 45180
rect 50378 45126 50380 45178
rect 50442 45126 50454 45178
rect 50516 45126 50518 45178
rect 50356 45124 50380 45126
rect 50436 45124 50460 45126
rect 50516 45124 50540 45126
rect 50300 45104 50596 45124
rect 31484 45076 31536 45082
rect 31484 45018 31536 45024
rect 31392 44940 31444 44946
rect 31392 44882 31444 44888
rect 31496 44810 31524 45018
rect 31944 45008 31996 45014
rect 31944 44950 31996 44956
rect 33968 45008 34020 45014
rect 33968 44950 34020 44956
rect 31484 44804 31536 44810
rect 31484 44746 31536 44752
rect 31956 44538 31984 44950
rect 32220 44940 32272 44946
rect 32220 44882 32272 44888
rect 32312 44940 32364 44946
rect 32312 44882 32364 44888
rect 32128 44804 32180 44810
rect 32128 44746 32180 44752
rect 32036 44736 32088 44742
rect 32036 44678 32088 44684
rect 31944 44532 31996 44538
rect 31944 44474 31996 44480
rect 32048 44334 32076 44678
rect 32140 44538 32168 44746
rect 32128 44532 32180 44538
rect 32128 44474 32180 44480
rect 32036 44328 32088 44334
rect 32036 44270 32088 44276
rect 32232 44266 32260 44882
rect 32220 44260 32272 44266
rect 32220 44202 32272 44208
rect 31944 44192 31996 44198
rect 31944 44134 31996 44140
rect 31956 43994 31984 44134
rect 31944 43988 31996 43994
rect 31944 43930 31996 43936
rect 31668 43784 31720 43790
rect 31668 43726 31720 43732
rect 31392 43648 31444 43654
rect 31392 43590 31444 43596
rect 31404 43246 31432 43590
rect 31392 43240 31444 43246
rect 31392 43182 31444 43188
rect 31680 42566 31708 43726
rect 31956 43654 31984 43930
rect 32232 43926 32260 44202
rect 32324 44198 32352 44882
rect 33048 44464 33100 44470
rect 33048 44406 33100 44412
rect 32312 44192 32364 44198
rect 32312 44134 32364 44140
rect 33060 43926 33088 44406
rect 33980 43994 34008 44950
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 33968 43988 34020 43994
rect 33968 43930 34020 43936
rect 32220 43920 32272 43926
rect 32220 43862 32272 43868
rect 33048 43920 33100 43926
rect 33048 43862 33100 43868
rect 32232 43790 32260 43862
rect 32220 43784 32272 43790
rect 32220 43726 32272 43732
rect 31944 43648 31996 43654
rect 31944 43590 31996 43596
rect 32232 43450 32260 43726
rect 32864 43648 32916 43654
rect 32864 43590 32916 43596
rect 32220 43444 32272 43450
rect 32220 43386 32272 43392
rect 32876 42770 32904 43590
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 32864 42764 32916 42770
rect 32864 42706 32916 42712
rect 31668 42560 31720 42566
rect 31668 42502 31720 42508
rect 31680 42294 31708 42502
rect 31668 42288 31720 42294
rect 31668 42230 31720 42236
rect 32680 42220 32732 42226
rect 32680 42162 32732 42168
rect 32128 42152 32180 42158
rect 32128 42094 32180 42100
rect 31484 42016 31536 42022
rect 31484 41958 31536 41964
rect 31496 41750 31524 41958
rect 32140 41818 32168 42094
rect 32128 41812 32180 41818
rect 32128 41754 32180 41760
rect 32692 41750 32720 42162
rect 31484 41744 31536 41750
rect 31484 41686 31536 41692
rect 32680 41744 32732 41750
rect 32680 41686 32732 41692
rect 31312 41386 31432 41414
rect 31300 40384 31352 40390
rect 31300 40326 31352 40332
rect 31312 39982 31340 40326
rect 31300 39976 31352 39982
rect 31300 39918 31352 39924
rect 31116 36032 31168 36038
rect 31116 35974 31168 35980
rect 31128 35834 31156 35974
rect 31116 35828 31168 35834
rect 31116 35770 31168 35776
rect 30944 34598 31064 34626
rect 30840 34400 30892 34406
rect 30840 34342 30892 34348
rect 30852 34134 30880 34342
rect 30840 34128 30892 34134
rect 30840 34070 30892 34076
rect 30944 32842 30972 34598
rect 31024 34536 31076 34542
rect 31024 34478 31076 34484
rect 31208 34536 31260 34542
rect 31208 34478 31260 34484
rect 31300 34536 31352 34542
rect 31300 34478 31352 34484
rect 31036 33590 31064 34478
rect 31024 33584 31076 33590
rect 31024 33526 31076 33532
rect 31220 33454 31248 34478
rect 31312 34202 31340 34478
rect 31300 34196 31352 34202
rect 31300 34138 31352 34144
rect 31312 33454 31340 34138
rect 31208 33448 31260 33454
rect 31208 33390 31260 33396
rect 31300 33448 31352 33454
rect 31300 33390 31352 33396
rect 30932 32836 30984 32842
rect 30932 32778 30984 32784
rect 31116 30388 31168 30394
rect 31116 30330 31168 30336
rect 30656 30184 30708 30190
rect 30656 30126 30708 30132
rect 30668 29510 30696 30126
rect 31128 29782 31156 30330
rect 31116 29776 31168 29782
rect 31116 29718 31168 29724
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 31208 29164 31260 29170
rect 31208 29106 31260 29112
rect 31116 29028 31168 29034
rect 31036 28988 31116 29016
rect 31036 28694 31064 28988
rect 31116 28970 31168 28976
rect 31114 28928 31170 28937
rect 31114 28863 31170 28872
rect 31024 28688 31076 28694
rect 31024 28630 31076 28636
rect 31128 28626 31156 28863
rect 31220 28694 31248 29106
rect 31298 28792 31354 28801
rect 31298 28727 31354 28736
rect 31208 28688 31260 28694
rect 31208 28630 31260 28636
rect 31116 28620 31168 28626
rect 31116 28562 31168 28568
rect 31220 28150 31248 28630
rect 31312 28490 31340 28727
rect 31300 28484 31352 28490
rect 31300 28426 31352 28432
rect 31208 28144 31260 28150
rect 31208 28086 31260 28092
rect 30840 28008 30892 28014
rect 30840 27950 30892 27956
rect 31208 28008 31260 28014
rect 31208 27950 31260 27956
rect 30852 27538 30880 27950
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 30564 26512 30616 26518
rect 30564 26454 30616 26460
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30564 25424 30616 25430
rect 30564 25366 30616 25372
rect 30472 25356 30524 25362
rect 30472 25298 30524 25304
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30392 24954 30420 25230
rect 30380 24948 30432 24954
rect 30380 24890 30432 24896
rect 30484 24410 30512 25298
rect 30472 24404 30524 24410
rect 30472 24346 30524 24352
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30300 23594 30328 24142
rect 30576 23866 30604 25366
rect 30944 25362 30972 27814
rect 31220 27334 31248 27950
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 31404 26926 31432 41386
rect 32692 41290 32720 41686
rect 32876 41546 32904 42706
rect 33232 42696 33284 42702
rect 33232 42638 33284 42644
rect 33140 42560 33192 42566
rect 33140 42502 33192 42508
rect 33152 42158 33180 42502
rect 33140 42152 33192 42158
rect 33140 42094 33192 42100
rect 33048 41608 33100 41614
rect 33048 41550 33100 41556
rect 32864 41540 32916 41546
rect 32864 41482 32916 41488
rect 33060 41414 33088 41550
rect 33244 41546 33272 42638
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 33324 42016 33376 42022
rect 33324 41958 33376 41964
rect 33336 41750 33364 41958
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 33324 41744 33376 41750
rect 33324 41686 33376 41692
rect 33232 41540 33284 41546
rect 33232 41482 33284 41488
rect 32968 41386 33088 41414
rect 32968 41290 32996 41386
rect 32692 41262 32996 41290
rect 31760 41064 31812 41070
rect 31760 41006 31812 41012
rect 32588 41064 32640 41070
rect 32588 41006 32640 41012
rect 33060 41018 33088 41386
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 33140 41064 33192 41070
rect 33060 41012 33140 41018
rect 33060 41006 33192 41012
rect 31576 40588 31628 40594
rect 31576 40530 31628 40536
rect 31588 39642 31616 40530
rect 31772 40526 31800 41006
rect 31852 40928 31904 40934
rect 31852 40870 31904 40876
rect 31864 40594 31892 40870
rect 32600 40730 32628 41006
rect 33060 40990 33180 41006
rect 32588 40724 32640 40730
rect 32588 40666 32640 40672
rect 31852 40588 31904 40594
rect 31852 40530 31904 40536
rect 31760 40520 31812 40526
rect 31760 40462 31812 40468
rect 31772 40186 31800 40462
rect 31852 40384 31904 40390
rect 31852 40326 31904 40332
rect 31760 40180 31812 40186
rect 31760 40122 31812 40128
rect 31864 40066 31892 40326
rect 31772 40038 31892 40066
rect 31576 39636 31628 39642
rect 31576 39578 31628 39584
rect 31772 39506 31800 40038
rect 33060 39642 33088 40990
rect 33140 40928 33192 40934
rect 33140 40870 33192 40876
rect 33152 39982 33180 40870
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 34060 40656 34112 40662
rect 34060 40598 34112 40604
rect 33876 40384 33928 40390
rect 33876 40326 33928 40332
rect 33140 39976 33192 39982
rect 33140 39918 33192 39924
rect 33416 39908 33468 39914
rect 33416 39850 33468 39856
rect 33048 39636 33100 39642
rect 33048 39578 33100 39584
rect 31760 39500 31812 39506
rect 31760 39442 31812 39448
rect 32128 39500 32180 39506
rect 32128 39442 32180 39448
rect 31772 38894 31800 39442
rect 32140 38962 32168 39442
rect 32864 39432 32916 39438
rect 32864 39374 32916 39380
rect 32128 38956 32180 38962
rect 32128 38898 32180 38904
rect 31760 38888 31812 38894
rect 31760 38830 31812 38836
rect 31668 38752 31720 38758
rect 31668 38694 31720 38700
rect 31680 38486 31708 38694
rect 32140 38554 32168 38898
rect 32404 38888 32456 38894
rect 32404 38830 32456 38836
rect 32416 38554 32444 38830
rect 32128 38548 32180 38554
rect 32128 38490 32180 38496
rect 32404 38548 32456 38554
rect 32404 38490 32456 38496
rect 31668 38480 31720 38486
rect 31668 38422 31720 38428
rect 32876 38418 32904 39374
rect 33048 39364 33100 39370
rect 33048 39306 33100 39312
rect 33060 38894 33088 39306
rect 33232 39296 33284 39302
rect 33232 39238 33284 39244
rect 33244 38894 33272 39238
rect 33428 38894 33456 39850
rect 33888 39574 33916 40326
rect 34072 40050 34100 40598
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34060 40044 34112 40050
rect 34060 39986 34112 39992
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50300 39664 50596 39684
rect 33876 39568 33928 39574
rect 33876 39510 33928 39516
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 33692 39024 33744 39030
rect 33692 38966 33744 38972
rect 33048 38888 33100 38894
rect 33048 38830 33100 38836
rect 33232 38888 33284 38894
rect 33232 38830 33284 38836
rect 33416 38888 33468 38894
rect 33416 38830 33468 38836
rect 32864 38412 32916 38418
rect 32864 38354 32916 38360
rect 33060 38282 33088 38830
rect 33244 38418 33272 38830
rect 33232 38412 33284 38418
rect 33232 38354 33284 38360
rect 33048 38276 33100 38282
rect 33048 38218 33100 38224
rect 33060 37738 33088 38218
rect 33324 37800 33376 37806
rect 33324 37742 33376 37748
rect 33048 37732 33100 37738
rect 33048 37674 33100 37680
rect 32220 37324 32272 37330
rect 32220 37266 32272 37272
rect 32232 36378 32260 37266
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32508 36718 32536 37062
rect 32496 36712 32548 36718
rect 32416 36660 32496 36666
rect 32416 36654 32548 36660
rect 32416 36638 32536 36654
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 32416 36242 32444 36638
rect 33060 36582 33088 37674
rect 33140 37324 33192 37330
rect 33140 37266 33192 37272
rect 32772 36576 32824 36582
rect 32772 36518 32824 36524
rect 33048 36576 33100 36582
rect 33048 36518 33100 36524
rect 32784 36242 32812 36518
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 32772 36236 32824 36242
rect 32772 36178 32824 36184
rect 33152 35698 33180 37266
rect 33336 36378 33364 37742
rect 33428 37330 33456 38830
rect 33704 38486 33732 38966
rect 33968 38820 34020 38826
rect 33968 38762 34020 38768
rect 33692 38480 33744 38486
rect 33692 38422 33744 38428
rect 33980 38282 34008 38762
rect 35256 38752 35308 38758
rect 35256 38694 35308 38700
rect 34152 38412 34204 38418
rect 34152 38354 34204 38360
rect 33968 38276 34020 38282
rect 33968 38218 34020 38224
rect 34164 38010 34192 38354
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34152 38004 34204 38010
rect 34152 37946 34204 37952
rect 35268 37806 35296 38694
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 34796 37800 34848 37806
rect 34796 37742 34848 37748
rect 35256 37800 35308 37806
rect 35256 37742 35308 37748
rect 33508 37732 33560 37738
rect 33508 37674 33560 37680
rect 33520 37398 33548 37674
rect 34520 37664 34572 37670
rect 34520 37606 34572 37612
rect 33508 37392 33560 37398
rect 33508 37334 33560 37340
rect 33416 37324 33468 37330
rect 33416 37266 33468 37272
rect 34532 36854 34560 37606
rect 34808 37466 34836 37742
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 34796 37460 34848 37466
rect 34796 37402 34848 37408
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34520 36848 34572 36854
rect 34520 36790 34572 36796
rect 33784 36780 33836 36786
rect 33784 36722 33836 36728
rect 33324 36372 33376 36378
rect 33324 36314 33376 36320
rect 33796 36242 33824 36722
rect 34532 36310 34560 36790
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 34520 36304 34572 36310
rect 34520 36246 34572 36252
rect 33784 36236 33836 36242
rect 33784 36178 33836 36184
rect 33796 36122 33824 36178
rect 33704 36094 33824 36122
rect 34244 36100 34296 36106
rect 33704 36038 33732 36094
rect 34244 36042 34296 36048
rect 33692 36032 33744 36038
rect 33692 35974 33744 35980
rect 33140 35692 33192 35698
rect 33140 35634 33192 35640
rect 31852 35624 31904 35630
rect 31852 35566 31904 35572
rect 31760 35488 31812 35494
rect 31760 35430 31812 35436
rect 31772 34542 31800 35430
rect 31864 35290 31892 35566
rect 31852 35284 31904 35290
rect 31852 35226 31904 35232
rect 33232 35148 33284 35154
rect 33232 35090 33284 35096
rect 33244 34746 33272 35090
rect 33704 35086 33732 35974
rect 34256 35698 34284 36042
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34244 35692 34296 35698
rect 34244 35634 34296 35640
rect 34980 35624 35032 35630
rect 34980 35566 35032 35572
rect 34428 35488 34480 35494
rect 34428 35430 34480 35436
rect 34440 35154 34468 35430
rect 34992 35290 35020 35566
rect 50300 35388 50596 35408
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 34980 35284 35032 35290
rect 34980 35226 35032 35232
rect 33784 35148 33836 35154
rect 33784 35090 33836 35096
rect 34428 35148 34480 35154
rect 34428 35090 34480 35096
rect 33692 35080 33744 35086
rect 33692 35022 33744 35028
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 33796 34678 33824 35090
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34152 34740 34204 34746
rect 34152 34682 34204 34688
rect 33784 34672 33836 34678
rect 33784 34614 33836 34620
rect 33876 34604 33928 34610
rect 33876 34546 33928 34552
rect 31760 34536 31812 34542
rect 31760 34478 31812 34484
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33048 34400 33100 34406
rect 33048 34342 33100 34348
rect 33060 34134 33088 34342
rect 33336 34134 33364 34478
rect 33888 34406 33916 34546
rect 34060 34536 34112 34542
rect 34060 34478 34112 34484
rect 33876 34400 33928 34406
rect 33876 34342 33928 34348
rect 33888 34202 33916 34342
rect 33876 34196 33928 34202
rect 33876 34138 33928 34144
rect 33048 34128 33100 34134
rect 33048 34070 33100 34076
rect 33324 34128 33376 34134
rect 33324 34070 33376 34076
rect 31852 33584 31904 33590
rect 31852 33526 31904 33532
rect 32956 33584 33008 33590
rect 32956 33526 33008 33532
rect 31864 32978 31892 33526
rect 32864 33448 32916 33454
rect 32864 33390 32916 33396
rect 32876 32978 32904 33390
rect 32968 33114 32996 33526
rect 33232 33448 33284 33454
rect 33232 33390 33284 33396
rect 33876 33448 33928 33454
rect 33876 33390 33928 33396
rect 32956 33108 33008 33114
rect 32956 33050 33008 33056
rect 31760 32972 31812 32978
rect 31760 32914 31812 32920
rect 31852 32972 31904 32978
rect 31852 32914 31904 32920
rect 32864 32972 32916 32978
rect 32864 32914 32916 32920
rect 31668 32904 31720 32910
rect 31668 32846 31720 32852
rect 31576 32768 31628 32774
rect 31576 32710 31628 32716
rect 31588 32366 31616 32710
rect 31680 32434 31708 32846
rect 31772 32502 31800 32914
rect 32968 32858 32996 33050
rect 33244 32910 33272 33390
rect 33232 32904 33284 32910
rect 32968 32830 33088 32858
rect 33232 32846 33284 32852
rect 31760 32496 31812 32502
rect 31760 32438 31812 32444
rect 31668 32428 31720 32434
rect 31668 32370 31720 32376
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 32968 31482 32996 31826
rect 33060 31498 33088 32830
rect 33244 32502 33272 32846
rect 33232 32496 33284 32502
rect 33232 32438 33284 32444
rect 33888 32366 33916 33390
rect 34072 33386 34100 34478
rect 34164 34066 34192 34682
rect 34244 34400 34296 34406
rect 34244 34342 34296 34348
rect 34152 34060 34204 34066
rect 34152 34002 34204 34008
rect 34060 33380 34112 33386
rect 34060 33322 34112 33328
rect 34060 32836 34112 32842
rect 34060 32778 34112 32784
rect 33876 32360 33928 32366
rect 33876 32302 33928 32308
rect 33888 32026 33916 32302
rect 33876 32020 33928 32026
rect 33876 31962 33928 31968
rect 33508 31680 33560 31686
rect 33508 31622 33560 31628
rect 33060 31482 33180 31498
rect 32956 31476 33008 31482
rect 33060 31476 33192 31482
rect 33060 31470 33140 31476
rect 32956 31418 33008 31424
rect 33140 31418 33192 31424
rect 33520 31346 33548 31622
rect 34072 31482 34100 32778
rect 34164 32774 34192 34002
rect 34256 33454 34284 34342
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 35348 34060 35400 34066
rect 35348 34002 35400 34008
rect 54116 34060 54168 34066
rect 54116 34002 54168 34008
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 35360 33590 35388 34002
rect 35900 33856 35952 33862
rect 35900 33798 35952 33804
rect 35348 33584 35400 33590
rect 35348 33526 35400 33532
rect 35912 33454 35940 33798
rect 54128 33658 54156 34002
rect 54116 33652 54168 33658
rect 54116 33594 54168 33600
rect 34244 33448 34296 33454
rect 34244 33390 34296 33396
rect 35900 33448 35952 33454
rect 35900 33390 35952 33396
rect 36176 33448 36228 33454
rect 36176 33390 36228 33396
rect 35716 33380 35768 33386
rect 35716 33322 35768 33328
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 34532 32978 34560 33254
rect 35728 33114 35756 33322
rect 35716 33108 35768 33114
rect 35716 33050 35768 33056
rect 34704 33040 34756 33046
rect 34704 32982 34756 32988
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 34152 32768 34204 32774
rect 34152 32710 34204 32716
rect 34244 32292 34296 32298
rect 34244 32234 34296 32240
rect 34256 32026 34284 32234
rect 34428 32224 34480 32230
rect 34428 32166 34480 32172
rect 34244 32020 34296 32026
rect 34244 31962 34296 31968
rect 34440 31890 34468 32166
rect 34428 31884 34480 31890
rect 34428 31826 34480 31832
rect 34520 31884 34572 31890
rect 34520 31826 34572 31832
rect 34532 31482 34560 31826
rect 34716 31822 34744 32982
rect 35912 32978 35940 33390
rect 35900 32972 35952 32978
rect 35900 32914 35952 32920
rect 36188 32910 36216 33390
rect 50300 33212 50596 33232
rect 50356 33210 50380 33212
rect 50436 33210 50460 33212
rect 50516 33210 50540 33212
rect 50378 33158 50380 33210
rect 50442 33158 50454 33210
rect 50516 33158 50518 33210
rect 50356 33156 50380 33158
rect 50436 33156 50460 33158
rect 50516 33156 50540 33158
rect 50300 33136 50596 33156
rect 53840 32972 53892 32978
rect 53840 32914 53892 32920
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 49976 32904 50028 32910
rect 49976 32846 50028 32852
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 35716 32224 35768 32230
rect 35716 32166 35768 32172
rect 35728 31890 35756 32166
rect 35716 31884 35768 31890
rect 35716 31826 35768 31832
rect 36188 31822 36216 32846
rect 49988 32298 50016 32846
rect 50344 32836 50396 32842
rect 50344 32778 50396 32784
rect 50356 32570 50384 32778
rect 50344 32564 50396 32570
rect 50344 32506 50396 32512
rect 53852 32434 53880 32914
rect 53840 32428 53892 32434
rect 53840 32370 53892 32376
rect 49976 32292 50028 32298
rect 49976 32234 50028 32240
rect 50300 32124 50596 32144
rect 50356 32122 50380 32124
rect 50436 32122 50460 32124
rect 50516 32122 50540 32124
rect 50378 32070 50380 32122
rect 50442 32070 50454 32122
rect 50516 32070 50518 32122
rect 50356 32068 50380 32070
rect 50436 32068 50460 32070
rect 50516 32068 50540 32070
rect 50300 32048 50596 32068
rect 53852 31890 53880 32370
rect 53840 31884 53892 31890
rect 53840 31826 53892 31832
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 36176 31816 36228 31822
rect 36176 31758 36228 31764
rect 34060 31476 34112 31482
rect 34060 31418 34112 31424
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 33508 31340 33560 31346
rect 33508 31282 33560 31288
rect 34716 31278 34744 31758
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34704 31272 34756 31278
rect 34704 31214 34756 31220
rect 36544 31204 36596 31210
rect 36544 31146 36596 31152
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 36556 30258 36584 31146
rect 50300 31036 50596 31056
rect 50356 31034 50380 31036
rect 50436 31034 50460 31036
rect 50516 31034 50540 31036
rect 50378 30982 50380 31034
rect 50442 30982 50454 31034
rect 50516 30982 50518 31034
rect 50356 30980 50380 30982
rect 50436 30980 50460 30982
rect 50516 30980 50540 30982
rect 50300 30960 50596 30980
rect 53852 30802 53880 31826
rect 53840 30796 53892 30802
rect 53840 30738 53892 30744
rect 50068 30320 50120 30326
rect 50068 30262 50120 30268
rect 36544 30252 36596 30258
rect 36544 30194 36596 30200
rect 31484 30184 31536 30190
rect 31484 30126 31536 30132
rect 35440 30184 35492 30190
rect 35440 30126 35492 30132
rect 31496 28966 31524 30126
rect 31588 29850 31800 29866
rect 31576 29844 31800 29850
rect 31628 29838 31800 29844
rect 31576 29786 31628 29792
rect 31772 29782 31800 29838
rect 31760 29776 31812 29782
rect 31760 29718 31812 29724
rect 31576 29572 31628 29578
rect 31576 29514 31628 29520
rect 31588 29102 31616 29514
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31576 29096 31628 29102
rect 31576 29038 31628 29044
rect 31484 28960 31536 28966
rect 31588 28937 31616 29038
rect 31484 28902 31536 28908
rect 31574 28928 31630 28937
rect 31496 28014 31524 28902
rect 31574 28863 31630 28872
rect 31772 28778 31800 29446
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 33324 29232 33376 29238
rect 33324 29174 33376 29180
rect 33140 29028 33192 29034
rect 33192 28976 33272 28994
rect 33140 28970 33272 28976
rect 33152 28966 33272 28970
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 31680 28750 31800 28778
rect 31680 28082 31708 28750
rect 32048 28626 32076 28902
rect 33244 28694 33272 28966
rect 33336 28801 33364 29174
rect 35452 29102 35480 30126
rect 50080 29782 50108 30262
rect 50160 30252 50212 30258
rect 50160 30194 50212 30200
rect 50172 29850 50200 30194
rect 50300 29948 50596 29968
rect 50356 29946 50380 29948
rect 50436 29946 50460 29948
rect 50516 29946 50540 29948
rect 50378 29894 50380 29946
rect 50442 29894 50454 29946
rect 50516 29894 50518 29946
rect 50356 29892 50380 29894
rect 50436 29892 50460 29894
rect 50516 29892 50540 29894
rect 50300 29872 50596 29892
rect 50160 29844 50212 29850
rect 50160 29786 50212 29792
rect 50068 29776 50120 29782
rect 50068 29718 50120 29724
rect 50252 29640 50304 29646
rect 50252 29582 50304 29588
rect 35624 29504 35676 29510
rect 35624 29446 35676 29452
rect 35636 29102 35664 29446
rect 50264 29170 50292 29582
rect 50344 29572 50396 29578
rect 50344 29514 50396 29520
rect 50356 29306 50384 29514
rect 50344 29300 50396 29306
rect 50344 29242 50396 29248
rect 50252 29164 50304 29170
rect 50252 29106 50304 29112
rect 33416 29096 33468 29102
rect 33416 29038 33468 29044
rect 33692 29096 33744 29102
rect 33692 29038 33744 29044
rect 35440 29096 35492 29102
rect 35440 29038 35492 29044
rect 35624 29096 35676 29102
rect 35624 29038 35676 29044
rect 36452 29096 36504 29102
rect 36452 29038 36504 29044
rect 33322 28792 33378 28801
rect 33322 28727 33378 28736
rect 32864 28688 32916 28694
rect 32864 28630 32916 28636
rect 33232 28688 33284 28694
rect 33232 28630 33284 28636
rect 31760 28620 31812 28626
rect 31760 28562 31812 28568
rect 31944 28620 31996 28626
rect 31944 28562 31996 28568
rect 32036 28620 32088 28626
rect 32036 28562 32088 28568
rect 31772 28082 31800 28562
rect 31668 28076 31720 28082
rect 31668 28018 31720 28024
rect 31760 28076 31812 28082
rect 31760 28018 31812 28024
rect 31484 28008 31536 28014
rect 31484 27950 31536 27956
rect 31680 27878 31708 28018
rect 31484 27872 31536 27878
rect 31484 27814 31536 27820
rect 31668 27872 31720 27878
rect 31668 27814 31720 27820
rect 31392 26920 31444 26926
rect 31392 26862 31444 26868
rect 31116 26852 31168 26858
rect 31116 26794 31168 26800
rect 31128 26518 31156 26794
rect 31116 26512 31168 26518
rect 31116 26454 31168 26460
rect 31116 25968 31168 25974
rect 31116 25910 31168 25916
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 30748 24268 30800 24274
rect 30748 24210 30800 24216
rect 30564 23860 30616 23866
rect 30564 23802 30616 23808
rect 30380 23724 30432 23730
rect 30380 23666 30432 23672
rect 30012 23588 30064 23594
rect 30012 23530 30064 23536
rect 30288 23588 30340 23594
rect 30288 23530 30340 23536
rect 30300 22574 30328 23530
rect 30392 23118 30420 23666
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30288 22568 30340 22574
rect 30288 22510 30340 22516
rect 30392 22506 30420 23054
rect 30576 22642 30604 23802
rect 30760 23662 30788 24210
rect 30852 24206 30880 24550
rect 30840 24200 30892 24206
rect 30840 24142 30892 24148
rect 31024 24132 31076 24138
rect 31024 24074 31076 24080
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30748 23656 30800 23662
rect 30748 23598 30800 23604
rect 30564 22636 30616 22642
rect 30564 22578 30616 22584
rect 30380 22500 30432 22506
rect 30380 22442 30432 22448
rect 30392 22094 30420 22442
rect 30760 22098 30788 23598
rect 30852 23254 30880 24006
rect 30932 23792 30984 23798
rect 30932 23734 30984 23740
rect 30840 23248 30892 23254
rect 30840 23190 30892 23196
rect 30944 22778 30972 23734
rect 31036 23662 31064 24074
rect 31024 23656 31076 23662
rect 31024 23598 31076 23604
rect 31024 23520 31076 23526
rect 31024 23462 31076 23468
rect 31036 23186 31064 23462
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 30932 22772 30984 22778
rect 30932 22714 30984 22720
rect 30840 22160 30892 22166
rect 30838 22128 30840 22137
rect 30892 22128 30894 22137
rect 30392 22066 30512 22094
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 21078 30420 21286
rect 30380 21072 30432 21078
rect 30380 21014 30432 21020
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29552 19304 29604 19310
rect 29552 19246 29604 19252
rect 29828 19304 29880 19310
rect 29828 19246 29880 19252
rect 30484 18834 30512 22066
rect 30748 22092 30800 22098
rect 31128 22094 31156 25910
rect 31208 25832 31260 25838
rect 31208 25774 31260 25780
rect 31220 25498 31248 25774
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31312 25362 31340 25638
rect 31300 25356 31352 25362
rect 31300 25298 31352 25304
rect 31300 25220 31352 25226
rect 31300 25162 31352 25168
rect 31312 24818 31340 25162
rect 31300 24812 31352 24818
rect 31300 24754 31352 24760
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 31404 23662 31432 24550
rect 31496 24313 31524 27814
rect 31668 27600 31720 27606
rect 31668 27542 31720 27548
rect 31680 27334 31708 27542
rect 31772 27402 31800 28018
rect 31956 27878 31984 28562
rect 32048 28014 32076 28562
rect 32876 28558 32904 28630
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32864 28552 32916 28558
rect 32864 28494 32916 28500
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 31944 27872 31996 27878
rect 31944 27814 31996 27820
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31668 27328 31720 27334
rect 31668 27270 31720 27276
rect 31956 26926 31984 27814
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 31852 26784 31904 26790
rect 32048 26738 32076 27406
rect 32220 27056 32272 27062
rect 32220 26998 32272 27004
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 31852 26726 31904 26732
rect 31864 25838 31892 26726
rect 31956 26710 32076 26738
rect 31956 26586 31984 26710
rect 32140 26586 32168 26930
rect 31944 26580 31996 26586
rect 31944 26522 31996 26528
rect 32128 26580 32180 26586
rect 32128 26522 32180 26528
rect 31852 25832 31904 25838
rect 31852 25774 31904 25780
rect 31864 25362 31892 25774
rect 31852 25356 31904 25362
rect 31852 25298 31904 25304
rect 31760 25220 31812 25226
rect 31760 25162 31812 25168
rect 31668 24812 31720 24818
rect 31668 24754 31720 24760
rect 31680 24410 31708 24754
rect 31668 24404 31720 24410
rect 31668 24346 31720 24352
rect 31482 24304 31538 24313
rect 31482 24239 31538 24248
rect 31772 24206 31800 25162
rect 31484 24200 31536 24206
rect 31484 24142 31536 24148
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 31392 23656 31444 23662
rect 31392 23598 31444 23604
rect 31392 23520 31444 23526
rect 31392 23462 31444 23468
rect 31208 23180 31260 23186
rect 31208 23122 31260 23128
rect 31220 22778 31248 23122
rect 31404 23118 31432 23462
rect 31300 23112 31352 23118
rect 31392 23112 31444 23118
rect 31300 23054 31352 23060
rect 31390 23080 31392 23089
rect 31444 23080 31446 23089
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31220 22574 31248 22714
rect 31208 22568 31260 22574
rect 31208 22510 31260 22516
rect 31312 22098 31340 23054
rect 31390 23015 31446 23024
rect 31392 22772 31444 22778
rect 31392 22714 31444 22720
rect 31404 22166 31432 22714
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 30838 22063 30894 22072
rect 31036 22066 31156 22094
rect 31300 22092 31352 22098
rect 30748 22034 30800 22040
rect 30932 21616 30984 21622
rect 30760 21564 30932 21570
rect 30760 21558 30984 21564
rect 30760 21554 30972 21558
rect 30748 21548 30972 21554
rect 30800 21542 30972 21548
rect 30748 21490 30800 21496
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30656 21480 30708 21486
rect 30656 21422 30708 21428
rect 30576 19242 30604 21422
rect 30668 20602 30696 21422
rect 31036 21146 31064 22066
rect 31300 22034 31352 22040
rect 31116 21956 31168 21962
rect 31116 21898 31168 21904
rect 31128 21570 31156 21898
rect 31312 21894 31340 22034
rect 31300 21888 31352 21894
rect 31300 21830 31352 21836
rect 31404 21690 31432 22102
rect 31392 21684 31444 21690
rect 31392 21626 31444 21632
rect 31128 21542 31248 21570
rect 31220 21486 31248 21542
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31024 21140 31076 21146
rect 31024 21082 31076 21088
rect 31220 21010 31248 21422
rect 31404 21010 31432 21626
rect 31496 21554 31524 24142
rect 31576 23588 31628 23594
rect 31576 23530 31628 23536
rect 31588 23186 31616 23530
rect 31772 23254 31800 24142
rect 31956 23662 31984 26522
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 32048 24954 32076 25094
rect 32036 24948 32088 24954
rect 32036 24890 32088 24896
rect 32140 24834 32168 25842
rect 32048 24806 32168 24834
rect 32048 24274 32076 24806
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 31944 23656 31996 23662
rect 31944 23598 31996 23604
rect 31944 23520 31996 23526
rect 31944 23462 31996 23468
rect 31760 23248 31812 23254
rect 31760 23190 31812 23196
rect 31576 23180 31628 23186
rect 31576 23122 31628 23128
rect 31588 22642 31616 23122
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31772 22506 31800 23054
rect 31760 22500 31812 22506
rect 31760 22442 31812 22448
rect 31956 22438 31984 23462
rect 32048 22438 32076 24210
rect 32232 23866 32260 26998
rect 32600 26450 32628 28494
rect 32876 27470 32904 28494
rect 32956 27532 33008 27538
rect 32956 27474 33008 27480
rect 33048 27532 33100 27538
rect 33048 27474 33100 27480
rect 32864 27464 32916 27470
rect 32864 27406 32916 27412
rect 32864 27328 32916 27334
rect 32864 27270 32916 27276
rect 32772 26784 32824 26790
rect 32772 26726 32824 26732
rect 32784 26450 32812 26726
rect 32876 26450 32904 27270
rect 32968 26518 32996 27474
rect 33060 27130 33088 27474
rect 33048 27124 33100 27130
rect 33048 27066 33100 27072
rect 33336 26926 33364 28727
rect 33428 28694 33456 29038
rect 33508 29006 33560 29012
rect 33508 28948 33560 28954
rect 33416 28688 33468 28694
rect 33416 28630 33468 28636
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33428 27062 33456 27406
rect 33416 27056 33468 27062
rect 33416 26998 33468 27004
rect 33520 26926 33548 28948
rect 33704 28762 33732 29038
rect 33692 28756 33744 28762
rect 33692 28698 33744 28704
rect 33784 28620 33836 28626
rect 33784 28562 33836 28568
rect 33796 28082 33824 28562
rect 35452 28422 35480 29038
rect 35716 28620 35768 28626
rect 35716 28562 35768 28568
rect 35440 28416 35492 28422
rect 35440 28358 35492 28364
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 35452 28014 35480 28358
rect 34336 28008 34388 28014
rect 34334 27976 34336 27985
rect 35440 28008 35492 28014
rect 34388 27976 34390 27985
rect 35440 27950 35492 27956
rect 35532 28008 35584 28014
rect 35532 27950 35584 27956
rect 34334 27911 34390 27920
rect 34612 27940 34664 27946
rect 34612 27882 34664 27888
rect 34624 27674 34652 27882
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34796 27328 34848 27334
rect 34796 27270 34848 27276
rect 33784 26988 33836 26994
rect 33784 26930 33836 26936
rect 34704 26988 34756 26994
rect 34704 26930 34756 26936
rect 33324 26920 33376 26926
rect 33244 26880 33324 26908
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 32956 26512 33008 26518
rect 32956 26454 33008 26460
rect 33060 26450 33088 26794
rect 32312 26444 32364 26450
rect 32588 26444 32640 26450
rect 32312 26386 32364 26392
rect 32508 26404 32588 26432
rect 32324 25498 32352 26386
rect 32404 26376 32456 26382
rect 32404 26318 32456 26324
rect 32416 25838 32444 26318
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32312 25492 32364 25498
rect 32312 25434 32364 25440
rect 32416 25362 32444 25774
rect 32404 25356 32456 25362
rect 32404 25298 32456 25304
rect 32404 24676 32456 24682
rect 32404 24618 32456 24624
rect 32416 24274 32444 24618
rect 32404 24268 32456 24274
rect 32404 24210 32456 24216
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 32508 23746 32536 26404
rect 32588 26386 32640 26392
rect 32772 26444 32824 26450
rect 32772 26386 32824 26392
rect 32864 26444 32916 26450
rect 32864 26386 32916 26392
rect 33048 26444 33100 26450
rect 33048 26386 33100 26392
rect 33060 26042 33088 26386
rect 32588 26036 32640 26042
rect 32588 25978 32640 25984
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 32600 25906 32628 25978
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32600 25294 32628 25842
rect 32680 25764 32732 25770
rect 32680 25706 32732 25712
rect 32692 25294 32720 25706
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25362 33180 25638
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 32588 25288 32640 25294
rect 32588 25230 32640 25236
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 32600 24750 32628 25230
rect 32692 24954 32720 25230
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32600 24410 32628 24686
rect 32680 24608 32732 24614
rect 32680 24550 32732 24556
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32692 24274 32720 24550
rect 32680 24268 32732 24274
rect 32680 24210 32732 24216
rect 33140 24268 33192 24274
rect 33140 24210 33192 24216
rect 33152 23866 33180 24210
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 32232 23718 32536 23746
rect 32232 23186 32260 23718
rect 33244 23662 33272 26880
rect 33508 26920 33560 26926
rect 33324 26862 33376 26868
rect 33506 26888 33508 26897
rect 33692 26920 33744 26926
rect 33560 26888 33562 26897
rect 33692 26862 33744 26868
rect 33506 26823 33562 26832
rect 33324 25968 33376 25974
rect 33324 25910 33376 25916
rect 33336 24886 33364 25910
rect 33324 24880 33376 24886
rect 33324 24822 33376 24828
rect 33336 24682 33364 24822
rect 33324 24676 33376 24682
rect 33324 24618 33376 24624
rect 33520 23662 33548 26823
rect 33704 26586 33732 26862
rect 33692 26580 33744 26586
rect 33692 26522 33744 26528
rect 33796 26518 33824 26930
rect 33784 26512 33836 26518
rect 33784 26454 33836 26460
rect 33968 26444 34020 26450
rect 33968 26386 34020 26392
rect 33980 25974 34008 26386
rect 34520 26308 34572 26314
rect 34520 26250 34572 26256
rect 33968 25968 34020 25974
rect 33968 25910 34020 25916
rect 34244 25968 34296 25974
rect 34244 25910 34296 25916
rect 34060 25832 34112 25838
rect 34060 25774 34112 25780
rect 34072 25362 34100 25774
rect 34256 25362 34284 25910
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 34348 25498 34376 25842
rect 34532 25702 34560 26250
rect 34428 25696 34480 25702
rect 34428 25638 34480 25644
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34440 25498 34468 25638
rect 34336 25492 34388 25498
rect 34336 25434 34388 25440
rect 34428 25492 34480 25498
rect 34428 25434 34480 25440
rect 33692 25356 33744 25362
rect 33692 25298 33744 25304
rect 33968 25356 34020 25362
rect 33968 25298 34020 25304
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 34244 25356 34296 25362
rect 34244 25298 34296 25304
rect 33704 24750 33732 25298
rect 33980 24818 34008 25298
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 33692 24744 33744 24750
rect 33692 24686 33744 24692
rect 33980 23662 34008 24754
rect 34440 24750 34468 25434
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34152 24064 34204 24070
rect 34152 24006 34204 24012
rect 33232 23656 33284 23662
rect 33508 23656 33560 23662
rect 33284 23616 33364 23644
rect 33232 23598 33284 23604
rect 32220 23180 32272 23186
rect 32140 23140 32220 23168
rect 31944 22432 31996 22438
rect 31944 22374 31996 22380
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 32036 22092 32088 22098
rect 32140 22080 32168 23140
rect 32220 23122 32272 23128
rect 32404 23180 32456 23186
rect 32404 23122 32456 23128
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32324 22658 32352 22918
rect 32416 22778 32444 23122
rect 32404 22772 32456 22778
rect 32404 22714 32456 22720
rect 32220 22636 32272 22642
rect 32324 22630 32444 22658
rect 32220 22578 32272 22584
rect 32232 22234 32260 22578
rect 32416 22506 32444 22630
rect 33232 22568 33284 22574
rect 33232 22510 33284 22516
rect 32404 22500 32456 22506
rect 32404 22442 32456 22448
rect 32312 22432 32364 22438
rect 32312 22374 32364 22380
rect 32220 22228 32272 22234
rect 32220 22170 32272 22176
rect 32324 22166 32352 22374
rect 33244 22234 33272 22510
rect 33232 22228 33284 22234
rect 33232 22170 33284 22176
rect 32312 22160 32364 22166
rect 32312 22102 32364 22108
rect 32088 22052 32168 22080
rect 32220 22092 32272 22098
rect 32036 22034 32088 22040
rect 32220 22034 32272 22040
rect 32496 22092 32548 22098
rect 32496 22034 32548 22040
rect 32232 21622 32260 22034
rect 32220 21616 32272 21622
rect 32220 21558 32272 21564
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31484 21412 31536 21418
rect 31484 21354 31536 21360
rect 31496 21146 31524 21354
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 32508 21049 32536 22034
rect 32956 21888 33008 21894
rect 32956 21830 33008 21836
rect 33140 21888 33192 21894
rect 33140 21830 33192 21836
rect 32968 21146 32996 21830
rect 33048 21412 33100 21418
rect 33048 21354 33100 21360
rect 32956 21140 33008 21146
rect 32956 21082 33008 21088
rect 32494 21040 32550 21049
rect 31208 21004 31260 21010
rect 31208 20946 31260 20952
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31576 21004 31628 21010
rect 32494 20975 32550 20984
rect 32588 21004 32640 21010
rect 31576 20946 31628 20952
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30656 20596 30708 20602
rect 30656 20538 30708 20544
rect 30944 20534 30972 20878
rect 30932 20528 30984 20534
rect 30932 20470 30984 20476
rect 30932 20324 30984 20330
rect 30932 20266 30984 20272
rect 30944 19854 30972 20266
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 30932 19848 30984 19854
rect 30932 19790 30984 19796
rect 30944 19514 30972 19790
rect 30932 19508 30984 19514
rect 30932 19450 30984 19456
rect 30564 19236 30616 19242
rect 30564 19178 30616 19184
rect 31036 18970 31064 19858
rect 31220 19310 31248 20946
rect 31588 20466 31616 20946
rect 32508 20874 32536 20975
rect 32588 20946 32640 20952
rect 32496 20868 32548 20874
rect 32496 20810 32548 20816
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31956 20466 31984 20742
rect 31576 20460 31628 20466
rect 31576 20402 31628 20408
rect 31944 20460 31996 20466
rect 31944 20402 31996 20408
rect 31484 20392 31536 20398
rect 31484 20334 31536 20340
rect 31496 19310 31524 20334
rect 31208 19304 31260 19310
rect 31208 19246 31260 19252
rect 31484 19304 31536 19310
rect 31484 19246 31536 19252
rect 31588 19174 31616 20402
rect 31116 19168 31168 19174
rect 31116 19110 31168 19116
rect 31576 19168 31628 19174
rect 31576 19110 31628 19116
rect 31024 18964 31076 18970
rect 31024 18906 31076 18912
rect 31128 18834 31156 19110
rect 29368 18828 29420 18834
rect 29368 18770 29420 18776
rect 30472 18828 30524 18834
rect 30472 18770 30524 18776
rect 30932 18828 30984 18834
rect 30932 18770 30984 18776
rect 31116 18828 31168 18834
rect 31116 18770 31168 18776
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26884 18216 26936 18222
rect 26884 18158 26936 18164
rect 28632 18216 28684 18222
rect 28632 18158 28684 18164
rect 30944 18154 30972 18770
rect 31956 18766 31984 20402
rect 32600 20330 32628 20946
rect 32864 20460 32916 20466
rect 32864 20402 32916 20408
rect 32588 20324 32640 20330
rect 32588 20266 32640 20272
rect 32600 19922 32628 20266
rect 32876 19922 32904 20402
rect 33060 20398 33088 21354
rect 33152 20398 33180 21830
rect 33244 21690 33272 22170
rect 33336 22166 33364 23616
rect 33508 23598 33560 23604
rect 33692 23656 33744 23662
rect 33692 23598 33744 23604
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33520 22760 33548 23598
rect 33704 23050 33732 23598
rect 34060 23588 34112 23594
rect 34164 23576 34192 24006
rect 34440 23798 34468 24686
rect 34428 23792 34480 23798
rect 34428 23734 34480 23740
rect 34244 23656 34296 23662
rect 34244 23598 34296 23604
rect 34112 23548 34192 23576
rect 34060 23530 34112 23536
rect 34164 23186 34192 23548
rect 34152 23180 34204 23186
rect 34152 23122 34204 23128
rect 33692 23044 33744 23050
rect 33692 22986 33744 22992
rect 33520 22732 33732 22760
rect 33600 22636 33652 22642
rect 33600 22578 33652 22584
rect 33612 22234 33640 22578
rect 33600 22228 33652 22234
rect 33600 22170 33652 22176
rect 33324 22160 33376 22166
rect 33324 22102 33376 22108
rect 33324 22024 33376 22030
rect 33324 21966 33376 21972
rect 33232 21684 33284 21690
rect 33232 21626 33284 21632
rect 33336 21486 33364 21966
rect 33612 21690 33640 22170
rect 33704 22098 33732 22732
rect 34164 22574 34192 23122
rect 34152 22568 34204 22574
rect 34152 22510 34204 22516
rect 33692 22092 33744 22098
rect 33692 22034 33744 22040
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 33796 21894 33824 22034
rect 33784 21888 33836 21894
rect 33784 21830 33836 21836
rect 33600 21684 33652 21690
rect 33600 21626 33652 21632
rect 33692 21684 33744 21690
rect 33692 21626 33744 21632
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 33600 21480 33652 21486
rect 33704 21468 33732 21626
rect 34152 21616 34204 21622
rect 34152 21558 34204 21564
rect 33652 21440 33732 21468
rect 33600 21422 33652 21428
rect 33336 21078 33364 21422
rect 33324 21072 33376 21078
rect 33324 21014 33376 21020
rect 33336 20602 33364 21014
rect 33704 20942 33732 21440
rect 33876 21480 33928 21486
rect 33928 21440 34100 21468
rect 33876 21422 33928 21428
rect 34072 21350 34100 21440
rect 33968 21344 34020 21350
rect 33968 21286 34020 21292
rect 34060 21344 34112 21350
rect 34060 21286 34112 21292
rect 33980 21078 34008 21286
rect 34164 21146 34192 21558
rect 34256 21418 34284 23598
rect 34532 23526 34560 25638
rect 34612 25152 34664 25158
rect 34612 25094 34664 25100
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34520 23180 34572 23186
rect 34520 23122 34572 23128
rect 34426 23080 34482 23089
rect 34426 23015 34428 23024
rect 34480 23015 34482 23024
rect 34428 22986 34480 22992
rect 34532 22710 34560 23122
rect 34520 22704 34572 22710
rect 34520 22646 34572 22652
rect 34624 22506 34652 25094
rect 34716 24750 34744 26930
rect 34808 26518 34836 27270
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 35544 27130 35572 27950
rect 35728 27538 35756 28562
rect 36464 28121 36492 29038
rect 50300 28860 50596 28880
rect 50356 28858 50380 28860
rect 50436 28858 50460 28860
rect 50516 28858 50540 28860
rect 50378 28806 50380 28858
rect 50442 28806 50454 28858
rect 50516 28806 50518 28858
rect 50356 28804 50380 28806
rect 50436 28804 50460 28806
rect 50516 28804 50540 28806
rect 50300 28784 50596 28804
rect 36450 28112 36506 28121
rect 36450 28047 36506 28056
rect 36268 28008 36320 28014
rect 36320 27968 36400 27996
rect 36268 27950 36320 27956
rect 35716 27532 35768 27538
rect 35716 27474 35768 27480
rect 35532 27124 35584 27130
rect 35532 27066 35584 27072
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 34796 26512 34848 26518
rect 34796 26454 34848 26460
rect 34808 25838 34836 26454
rect 35256 26376 35308 26382
rect 35256 26318 35308 26324
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 35268 26042 35296 26318
rect 35256 26036 35308 26042
rect 35256 25978 35308 25984
rect 35636 25974 35664 26726
rect 35624 25968 35676 25974
rect 35624 25910 35676 25916
rect 35636 25838 35664 25910
rect 34796 25832 34848 25838
rect 34796 25774 34848 25780
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34704 24744 34756 24750
rect 34704 24686 34756 24692
rect 34716 24138 34744 24686
rect 34704 24132 34756 24138
rect 34704 24074 34756 24080
rect 34716 23730 34744 24074
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 35348 23656 35400 23662
rect 35348 23598 35400 23604
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 35360 22778 35388 23598
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 35348 22568 35400 22574
rect 35348 22510 35400 22516
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34520 21888 34572 21894
rect 34520 21830 34572 21836
rect 34244 21412 34296 21418
rect 34244 21354 34296 21360
rect 34532 21350 34560 21830
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 35360 21690 35388 22510
rect 35440 22432 35492 22438
rect 35440 22374 35492 22380
rect 35452 22234 35480 22374
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35452 21962 35480 22170
rect 35440 21956 35492 21962
rect 35440 21898 35492 21904
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 34612 21412 34664 21418
rect 34612 21354 34664 21360
rect 34520 21344 34572 21350
rect 34520 21286 34572 21292
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 33968 21072 34020 21078
rect 33968 21014 34020 21020
rect 34334 21040 34390 21049
rect 34334 20975 34336 20984
rect 34388 20975 34390 20984
rect 34336 20946 34388 20952
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33968 20936 34020 20942
rect 33968 20878 34020 20884
rect 33324 20596 33376 20602
rect 33324 20538 33376 20544
rect 33048 20392 33100 20398
rect 33048 20334 33100 20340
rect 33140 20392 33192 20398
rect 33140 20334 33192 20340
rect 32588 19916 32640 19922
rect 32588 19858 32640 19864
rect 32864 19916 32916 19922
rect 32864 19858 32916 19864
rect 33060 19514 33088 20334
rect 33980 19922 34008 20878
rect 34532 20466 34560 21286
rect 34624 20602 34652 21354
rect 35728 21078 35756 27474
rect 36372 27334 36400 27968
rect 50300 27772 50596 27792
rect 50356 27770 50380 27772
rect 50436 27770 50460 27772
rect 50516 27770 50540 27772
rect 50378 27718 50380 27770
rect 50442 27718 50454 27770
rect 50516 27718 50518 27770
rect 50356 27716 50380 27718
rect 50436 27716 50460 27718
rect 50516 27716 50540 27718
rect 50300 27696 50596 27716
rect 36360 27328 36412 27334
rect 36360 27270 36412 27276
rect 35808 26512 35860 26518
rect 35808 26454 35860 26460
rect 35820 25702 35848 26454
rect 36372 26450 36400 27270
rect 37188 26852 37240 26858
rect 37188 26794 37240 26800
rect 37200 26586 37228 26794
rect 50300 26684 50596 26704
rect 50356 26682 50380 26684
rect 50436 26682 50460 26684
rect 50516 26682 50540 26684
rect 50378 26630 50380 26682
rect 50442 26630 50454 26682
rect 50516 26630 50518 26682
rect 50356 26628 50380 26630
rect 50436 26628 50460 26630
rect 50516 26628 50540 26630
rect 50300 26608 50596 26628
rect 37188 26580 37240 26586
rect 37188 26522 37240 26528
rect 36636 26512 36688 26518
rect 36636 26454 36688 26460
rect 36360 26444 36412 26450
rect 36360 26386 36412 26392
rect 36372 25838 36400 26386
rect 36648 25906 36676 26454
rect 37096 26444 37148 26450
rect 37096 26386 37148 26392
rect 36636 25900 36688 25906
rect 36636 25842 36688 25848
rect 36360 25832 36412 25838
rect 36360 25774 36412 25780
rect 35992 25764 36044 25770
rect 35992 25706 36044 25712
rect 35808 25696 35860 25702
rect 35808 25638 35860 25644
rect 35900 25152 35952 25158
rect 35900 25094 35952 25100
rect 35912 24750 35940 25094
rect 36004 24954 36032 25706
rect 36372 25344 36400 25774
rect 37108 25362 37136 26386
rect 50300 25596 50596 25616
rect 50356 25594 50380 25596
rect 50436 25594 50460 25596
rect 50516 25594 50540 25596
rect 50378 25542 50380 25594
rect 50442 25542 50454 25594
rect 50516 25542 50518 25594
rect 50356 25540 50380 25542
rect 50436 25540 50460 25542
rect 50516 25540 50540 25542
rect 50300 25520 50596 25540
rect 36452 25356 36504 25362
rect 36372 25316 36452 25344
rect 36452 25298 36504 25304
rect 36544 25356 36596 25362
rect 36544 25298 36596 25304
rect 37096 25356 37148 25362
rect 37096 25298 37148 25304
rect 36084 25220 36136 25226
rect 36084 25162 36136 25168
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35900 24744 35952 24750
rect 35900 24686 35952 24692
rect 35808 24608 35860 24614
rect 35808 24550 35860 24556
rect 35820 24274 35848 24550
rect 36004 24410 36032 24890
rect 35992 24404 36044 24410
rect 35992 24346 36044 24352
rect 35808 24268 35860 24274
rect 35808 24210 35860 24216
rect 35992 23588 36044 23594
rect 35992 23530 36044 23536
rect 36004 22778 36032 23530
rect 35992 22772 36044 22778
rect 35992 22714 36044 22720
rect 36096 22658 36124 25162
rect 36464 24750 36492 25298
rect 36452 24744 36504 24750
rect 36452 24686 36504 24692
rect 36176 23520 36228 23526
rect 36176 23462 36228 23468
rect 36188 23254 36216 23462
rect 36176 23248 36228 23254
rect 36176 23190 36228 23196
rect 36556 23186 36584 25298
rect 36728 25288 36780 25294
rect 36728 25230 36780 25236
rect 36740 24750 36768 25230
rect 36636 24744 36688 24750
rect 36636 24686 36688 24692
rect 36728 24744 36780 24750
rect 36728 24686 36780 24692
rect 36648 23866 36676 24686
rect 50300 24508 50596 24528
rect 50356 24506 50380 24508
rect 50436 24506 50460 24508
rect 50516 24506 50540 24508
rect 50378 24454 50380 24506
rect 50442 24454 50454 24506
rect 50516 24454 50518 24506
rect 50356 24452 50380 24454
rect 50436 24452 50460 24454
rect 50516 24452 50540 24454
rect 50300 24432 50596 24452
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36544 23180 36596 23186
rect 36544 23122 36596 23128
rect 36556 23050 36584 23122
rect 36740 23118 36768 23462
rect 50300 23420 50596 23440
rect 50356 23418 50380 23420
rect 50436 23418 50460 23420
rect 50516 23418 50540 23420
rect 50378 23366 50380 23418
rect 50442 23366 50454 23418
rect 50516 23366 50518 23418
rect 50356 23364 50380 23366
rect 50436 23364 50460 23366
rect 50516 23364 50540 23366
rect 50300 23344 50596 23364
rect 54312 23322 54340 56238
rect 54588 55826 54616 56782
rect 54680 56438 54708 56902
rect 54760 56840 54812 56846
rect 54760 56782 54812 56788
rect 54772 56506 54800 56782
rect 55218 56536 55274 56545
rect 54760 56500 54812 56506
rect 55218 56471 55274 56480
rect 54760 56442 54812 56448
rect 54668 56432 54720 56438
rect 54668 56374 54720 56380
rect 54576 55820 54628 55826
rect 54576 55762 54628 55768
rect 55232 55214 55260 56471
rect 55220 55208 55272 55214
rect 55220 55150 55272 55156
rect 55324 54738 55352 58618
rect 55600 55214 55628 59200
rect 55678 59120 55734 59129
rect 55678 59055 55734 59064
rect 55692 57526 55720 59055
rect 56428 58682 56456 59200
rect 56416 58676 56468 58682
rect 56416 58618 56468 58624
rect 56414 58576 56470 58585
rect 56414 58511 56470 58520
rect 55680 57520 55732 57526
rect 55680 57462 55732 57468
rect 56428 57458 56456 58511
rect 56520 58313 56548 59599
rect 57150 59200 57206 60000
rect 57978 59200 58034 60000
rect 58714 59200 58770 60000
rect 59542 59200 59598 60000
rect 56506 58304 56562 58313
rect 56506 58239 56562 58248
rect 56508 58064 56560 58070
rect 56506 58032 56508 58041
rect 56560 58032 56562 58041
rect 56506 57967 56562 57976
rect 56416 57452 56468 57458
rect 56416 57394 56468 57400
rect 56784 57384 56836 57390
rect 56784 57326 56836 57332
rect 57164 57338 57192 59200
rect 57992 57474 58020 59200
rect 58162 57488 58218 57497
rect 57992 57446 58112 57474
rect 56600 56840 56652 56846
rect 56600 56782 56652 56788
rect 55772 56772 55824 56778
rect 55772 56714 55824 56720
rect 56416 56772 56468 56778
rect 56416 56714 56468 56720
rect 55784 56370 55812 56714
rect 56428 56506 56456 56714
rect 56416 56500 56468 56506
rect 56416 56442 56468 56448
rect 56508 56500 56560 56506
rect 56508 56442 56560 56448
rect 56140 56432 56192 56438
rect 56140 56374 56192 56380
rect 55772 56364 55824 56370
rect 55772 56306 55824 56312
rect 56048 55752 56100 55758
rect 56048 55694 56100 55700
rect 56060 55418 56088 55694
rect 56048 55412 56100 55418
rect 56048 55354 56100 55360
rect 55600 55186 55720 55214
rect 55586 54904 55642 54913
rect 55586 54839 55642 54848
rect 55600 54738 55628 54839
rect 55312 54732 55364 54738
rect 55312 54674 55364 54680
rect 55588 54732 55640 54738
rect 55588 54674 55640 54680
rect 55692 54126 55720 55186
rect 56152 54806 56180 56374
rect 56232 56364 56284 56370
rect 56232 56306 56284 56312
rect 56244 55690 56272 56306
rect 56232 55684 56284 55690
rect 56232 55626 56284 55632
rect 56140 54800 56192 54806
rect 56140 54742 56192 54748
rect 55680 54120 55732 54126
rect 55680 54062 55732 54068
rect 56520 53650 56548 56442
rect 56612 55826 56640 56782
rect 56692 56228 56744 56234
rect 56692 56170 56744 56176
rect 56704 55826 56732 56170
rect 56796 55962 56824 57326
rect 57164 57310 57284 57338
rect 57060 56976 57112 56982
rect 57058 56944 57060 56953
rect 57112 56944 57114 56953
rect 57058 56879 57114 56888
rect 57152 56908 57204 56914
rect 57152 56850 57204 56856
rect 56784 55956 56836 55962
rect 56784 55898 56836 55904
rect 56600 55820 56652 55826
rect 56600 55762 56652 55768
rect 56692 55820 56744 55826
rect 56692 55762 56744 55768
rect 56704 55214 56732 55762
rect 56612 55208 56744 55214
rect 56612 55186 56692 55208
rect 56508 53644 56560 53650
rect 56508 53586 56560 53592
rect 56506 53408 56562 53417
rect 56506 53343 56562 53352
rect 56520 53038 56548 53343
rect 56508 53032 56560 53038
rect 56508 52974 56560 52980
rect 56508 51944 56560 51950
rect 56508 51886 56560 51892
rect 56520 51785 56548 51886
rect 56506 51776 56562 51785
rect 56506 51711 56562 51720
rect 55036 49292 55088 49298
rect 55036 49234 55088 49240
rect 54944 43852 54996 43858
rect 54944 43794 54996 43800
rect 54484 33380 54536 33386
rect 54484 33322 54536 33328
rect 54496 32570 54524 33322
rect 54576 33040 54628 33046
rect 54576 32982 54628 32988
rect 54484 32564 54536 32570
rect 54484 32506 54536 32512
rect 54588 31754 54616 32982
rect 54956 32842 54984 43794
rect 55048 33522 55076 49234
rect 56508 48680 56560 48686
rect 56506 48648 56508 48657
rect 56560 48648 56562 48657
rect 56506 48583 56562 48592
rect 55680 47524 55732 47530
rect 55680 47466 55732 47472
rect 55310 34640 55366 34649
rect 55310 34575 55366 34584
rect 55324 34542 55352 34575
rect 55312 34536 55364 34542
rect 55312 34478 55364 34484
rect 55220 34060 55272 34066
rect 55220 34002 55272 34008
rect 55036 33516 55088 33522
rect 55036 33458 55088 33464
rect 55232 33017 55260 34002
rect 55218 33008 55274 33017
rect 55218 32943 55274 32952
rect 54944 32836 54996 32842
rect 54944 32778 54996 32784
rect 55496 32496 55548 32502
rect 55496 32438 55548 32444
rect 54668 32360 54720 32366
rect 54668 32302 54720 32308
rect 55036 32360 55088 32366
rect 55036 32302 55088 32308
rect 54680 31890 54708 32302
rect 54668 31884 54720 31890
rect 54668 31826 54720 31832
rect 54576 31748 54628 31754
rect 54576 31690 54628 31696
rect 54576 31204 54628 31210
rect 54576 31146 54628 31152
rect 54588 30938 54616 31146
rect 55048 31142 55076 32302
rect 55220 31952 55272 31958
rect 55220 31894 55272 31900
rect 55232 31822 55260 31894
rect 55220 31816 55272 31822
rect 55220 31758 55272 31764
rect 55036 31136 55088 31142
rect 55036 31078 55088 31084
rect 54576 30932 54628 30938
rect 54576 30874 54628 30880
rect 55048 30802 55076 31078
rect 55036 30796 55088 30802
rect 55036 30738 55088 30744
rect 55508 30326 55536 32438
rect 55692 32026 55720 47466
rect 56506 45520 56562 45529
rect 56506 45455 56562 45464
rect 56520 45422 56548 45455
rect 56508 45416 56560 45422
rect 56508 45358 56560 45364
rect 56506 44024 56562 44033
rect 56506 43959 56562 43968
rect 56520 43246 56548 43959
rect 56508 43240 56560 43246
rect 56508 43182 56560 43188
rect 56506 42392 56562 42401
rect 56506 42327 56562 42336
rect 56520 42158 56548 42327
rect 56508 42152 56560 42158
rect 56508 42094 56560 42100
rect 56508 41064 56560 41070
rect 56508 41006 56560 41012
rect 56520 40905 56548 41006
rect 56506 40896 56562 40905
rect 56506 40831 56562 40840
rect 56508 37800 56560 37806
rect 56506 37768 56508 37777
rect 56560 37768 56562 37777
rect 56506 37703 56562 37712
rect 56230 36136 56286 36145
rect 56230 36071 56286 36080
rect 56244 35630 56272 36071
rect 56232 35624 56284 35630
rect 56232 35566 56284 35572
rect 55864 34060 55916 34066
rect 55864 34002 55916 34008
rect 55772 33856 55824 33862
rect 55772 33798 55824 33804
rect 55784 33386 55812 33798
rect 55772 33380 55824 33386
rect 55772 33322 55824 33328
rect 55876 33114 55904 34002
rect 55864 33108 55916 33114
rect 55864 33050 55916 33056
rect 55876 32434 55904 33050
rect 56232 32972 56284 32978
rect 56232 32914 56284 32920
rect 55864 32428 55916 32434
rect 55864 32370 55916 32376
rect 55680 32020 55732 32026
rect 55680 31962 55732 31968
rect 56244 31278 56272 32914
rect 56416 32020 56468 32026
rect 56416 31962 56468 31968
rect 56232 31272 56284 31278
rect 56232 31214 56284 31220
rect 55772 31136 55824 31142
rect 55772 31078 55824 31084
rect 55784 30870 55812 31078
rect 55772 30864 55824 30870
rect 55772 30806 55824 30812
rect 55680 30592 55732 30598
rect 55680 30534 55732 30540
rect 55496 30320 55548 30326
rect 55496 30262 55548 30268
rect 55692 30258 55720 30534
rect 55680 30252 55732 30258
rect 55680 30194 55732 30200
rect 54944 30184 54996 30190
rect 54944 30126 54996 30132
rect 56140 30184 56192 30190
rect 56140 30126 56192 30132
rect 54852 29776 54904 29782
rect 54852 29718 54904 29724
rect 54484 29708 54536 29714
rect 54484 29650 54536 29656
rect 54496 29510 54524 29650
rect 54484 29504 54536 29510
rect 54484 29446 54536 29452
rect 54864 29306 54892 29718
rect 54956 29714 54984 30126
rect 55404 30116 55456 30122
rect 55404 30058 55456 30064
rect 55416 29850 55444 30058
rect 56048 30048 56100 30054
rect 56048 29990 56100 29996
rect 55404 29844 55456 29850
rect 55404 29786 55456 29792
rect 56060 29782 56088 29990
rect 56048 29776 56100 29782
rect 56048 29718 56100 29724
rect 54944 29708 54996 29714
rect 54996 29668 55260 29696
rect 54944 29650 54996 29656
rect 54852 29300 54904 29306
rect 54852 29242 54904 29248
rect 55232 29238 55260 29668
rect 56152 29306 56180 30126
rect 56140 29300 56192 29306
rect 56140 29242 56192 29248
rect 55220 29232 55272 29238
rect 55220 29174 55272 29180
rect 55232 29102 55260 29174
rect 56244 29102 56272 31214
rect 56428 30938 56456 31962
rect 56506 31512 56562 31521
rect 56506 31447 56562 31456
rect 56520 31414 56548 31447
rect 56508 31408 56560 31414
rect 56508 31350 56560 31356
rect 56416 30932 56468 30938
rect 56416 30874 56468 30880
rect 56506 29880 56562 29889
rect 56506 29815 56562 29824
rect 56520 29510 56548 29815
rect 56508 29504 56560 29510
rect 56508 29446 56560 29452
rect 55220 29096 55272 29102
rect 55220 29038 55272 29044
rect 55680 29096 55732 29102
rect 55680 29038 55732 29044
rect 56232 29096 56284 29102
rect 56232 29038 56284 29044
rect 55128 28552 55180 28558
rect 55128 28494 55180 28500
rect 55140 27946 55168 28494
rect 55232 28014 55260 29038
rect 55312 28688 55364 28694
rect 55312 28630 55364 28636
rect 55324 28218 55352 28630
rect 55588 28484 55640 28490
rect 55588 28426 55640 28432
rect 55600 28393 55628 28426
rect 55586 28384 55642 28393
rect 55586 28319 55642 28328
rect 55312 28212 55364 28218
rect 55312 28154 55364 28160
rect 55220 28008 55272 28014
rect 55220 27950 55272 27956
rect 55128 27940 55180 27946
rect 55128 27882 55180 27888
rect 55588 27532 55640 27538
rect 55588 27474 55640 27480
rect 55404 26852 55456 26858
rect 55404 26794 55456 26800
rect 55496 26852 55548 26858
rect 55496 26794 55548 26800
rect 55416 26314 55444 26794
rect 55404 26308 55456 26314
rect 55404 26250 55456 26256
rect 55508 26042 55536 26794
rect 55600 26761 55628 27474
rect 55586 26752 55642 26761
rect 55586 26687 55642 26696
rect 55692 26234 55720 29038
rect 56232 28688 56284 28694
rect 56232 28630 56284 28636
rect 56244 28218 56272 28630
rect 56232 28212 56284 28218
rect 56232 28154 56284 28160
rect 56048 27532 56100 27538
rect 56048 27474 56100 27480
rect 55956 26376 56008 26382
rect 55956 26318 56008 26324
rect 55600 26206 55720 26234
rect 55496 26036 55548 26042
rect 55496 25978 55548 25984
rect 55600 25498 55628 26206
rect 55968 26042 55996 26318
rect 55956 26036 56008 26042
rect 55956 25978 56008 25984
rect 55680 25832 55732 25838
rect 55680 25774 55732 25780
rect 55588 25492 55640 25498
rect 55588 25434 55640 25440
rect 55692 25362 55720 25774
rect 55680 25356 55732 25362
rect 55680 25298 55732 25304
rect 55404 25152 55456 25158
rect 55404 25094 55456 25100
rect 55416 24818 55444 25094
rect 55404 24812 55456 24818
rect 55404 24754 55456 24760
rect 55692 24274 55720 25298
rect 55772 24744 55824 24750
rect 55772 24686 55824 24692
rect 55784 24410 55812 24686
rect 55772 24404 55824 24410
rect 55772 24346 55824 24352
rect 55680 24268 55732 24274
rect 55680 24210 55732 24216
rect 55588 23656 55640 23662
rect 55588 23598 55640 23604
rect 55220 23520 55272 23526
rect 55220 23462 55272 23468
rect 54300 23316 54352 23322
rect 54300 23258 54352 23264
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36544 23044 36596 23050
rect 36544 22986 36596 22992
rect 36004 22630 36124 22658
rect 36004 22574 36032 22630
rect 35992 22568 36044 22574
rect 35992 22510 36044 22516
rect 35716 21072 35768 21078
rect 35716 21014 35768 21020
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 36004 20330 36032 22510
rect 50300 22332 50596 22352
rect 50356 22330 50380 22332
rect 50436 22330 50460 22332
rect 50516 22330 50540 22332
rect 50378 22278 50380 22330
rect 50442 22278 50454 22330
rect 50516 22278 50518 22330
rect 50356 22276 50380 22278
rect 50436 22276 50460 22278
rect 50516 22276 50540 22278
rect 50300 22256 50596 22276
rect 38764 22234 39160 22250
rect 38752 22228 39160 22234
rect 38804 22222 39160 22228
rect 38752 22170 38804 22176
rect 39132 22166 39160 22222
rect 39120 22160 39172 22166
rect 36266 22128 36322 22137
rect 36084 22092 36136 22098
rect 39120 22102 39172 22108
rect 36266 22063 36268 22072
rect 36084 22034 36136 22040
rect 36320 22063 36322 22072
rect 36268 22034 36320 22040
rect 36096 21486 36124 22034
rect 48044 22024 48096 22030
rect 48044 21966 48096 21972
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 36096 21010 36124 21422
rect 48056 21418 48084 21966
rect 48044 21412 48096 21418
rect 48044 21354 48096 21360
rect 50300 21244 50596 21264
rect 50356 21242 50380 21244
rect 50436 21242 50460 21244
rect 50516 21242 50540 21244
rect 50378 21190 50380 21242
rect 50442 21190 50454 21242
rect 50516 21190 50518 21242
rect 50356 21188 50380 21190
rect 50436 21188 50460 21190
rect 50516 21188 50540 21190
rect 50300 21168 50596 21188
rect 36084 21004 36136 21010
rect 36084 20946 36136 20952
rect 36096 20806 36124 20946
rect 36452 20936 36504 20942
rect 36452 20878 36504 20884
rect 36084 20800 36136 20806
rect 36084 20742 36136 20748
rect 36096 20398 36124 20742
rect 36464 20466 36492 20878
rect 36452 20460 36504 20466
rect 36452 20402 36504 20408
rect 36084 20392 36136 20398
rect 36084 20334 36136 20340
rect 36268 20392 36320 20398
rect 36268 20334 36320 20340
rect 35992 20324 36044 20330
rect 35992 20266 36044 20272
rect 36280 19990 36308 20334
rect 50300 20156 50596 20176
rect 50356 20154 50380 20156
rect 50436 20154 50460 20156
rect 50516 20154 50540 20156
rect 50378 20102 50380 20154
rect 50442 20102 50454 20154
rect 50516 20102 50518 20154
rect 50356 20100 50380 20102
rect 50436 20100 50460 20102
rect 50516 20100 50540 20102
rect 50300 20080 50596 20100
rect 50988 20052 51040 20058
rect 50988 19994 51040 20000
rect 36268 19984 36320 19990
rect 36268 19926 36320 19932
rect 33968 19916 34020 19922
rect 33968 19858 34020 19864
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 33048 19508 33100 19514
rect 33048 19450 33100 19456
rect 50300 19068 50596 19088
rect 50356 19066 50380 19068
rect 50436 19066 50460 19068
rect 50516 19066 50540 19068
rect 50378 19014 50380 19066
rect 50442 19014 50454 19066
rect 50516 19014 50518 19066
rect 50356 19012 50380 19014
rect 50436 19012 50460 19014
rect 50516 19012 50540 19014
rect 50300 18992 50596 19012
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 30932 18148 30984 18154
rect 30932 18090 30984 18096
rect 50300 17980 50596 18000
rect 50356 17978 50380 17980
rect 50436 17978 50460 17980
rect 50516 17978 50540 17980
rect 50378 17926 50380 17978
rect 50442 17926 50454 17978
rect 50516 17926 50518 17978
rect 50356 17924 50380 17926
rect 50436 17924 50460 17926
rect 50516 17924 50540 17926
rect 50300 17904 50596 17924
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 50300 16892 50596 16912
rect 50356 16890 50380 16892
rect 50436 16890 50460 16892
rect 50516 16890 50540 16892
rect 50378 16838 50380 16890
rect 50442 16838 50454 16890
rect 50516 16838 50518 16890
rect 50356 16836 50380 16838
rect 50436 16836 50460 16838
rect 50516 16836 50540 16838
rect 50300 16816 50596 16836
rect 24216 16652 24268 16658
rect 24216 16594 24268 16600
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 34940 16348 35236 16368
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 50300 15804 50596 15824
rect 50356 15802 50380 15804
rect 50436 15802 50460 15804
rect 50516 15802 50540 15804
rect 50378 15750 50380 15802
rect 50442 15750 50454 15802
rect 50516 15750 50518 15802
rect 50356 15748 50380 15750
rect 50436 15748 50460 15750
rect 50516 15748 50540 15750
rect 50300 15728 50596 15748
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 50300 14716 50596 14736
rect 50356 14714 50380 14716
rect 50436 14714 50460 14716
rect 50516 14714 50540 14716
rect 50378 14662 50380 14714
rect 50442 14662 50454 14714
rect 50516 14662 50518 14714
rect 50356 14660 50380 14662
rect 50436 14660 50460 14662
rect 50516 14660 50540 14662
rect 50300 14640 50596 14660
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 50300 13628 50596 13648
rect 50356 13626 50380 13628
rect 50436 13626 50460 13628
rect 50516 13626 50540 13628
rect 50378 13574 50380 13626
rect 50442 13574 50454 13626
rect 50516 13574 50518 13626
rect 50356 13572 50380 13574
rect 50436 13572 50460 13574
rect 50516 13572 50540 13574
rect 50300 13552 50596 13572
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 50300 12540 50596 12560
rect 50356 12538 50380 12540
rect 50436 12538 50460 12540
rect 50516 12538 50540 12540
rect 50378 12486 50380 12538
rect 50442 12486 50454 12538
rect 50516 12486 50518 12538
rect 50356 12484 50380 12486
rect 50436 12484 50460 12486
rect 50516 12484 50540 12486
rect 50300 12464 50596 12484
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 50300 11452 50596 11472
rect 50356 11450 50380 11452
rect 50436 11450 50460 11452
rect 50516 11450 50540 11452
rect 50378 11398 50380 11450
rect 50442 11398 50454 11450
rect 50516 11398 50518 11450
rect 50356 11396 50380 11398
rect 50436 11396 50460 11398
rect 50516 11396 50540 11398
rect 50300 11376 50596 11396
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 50300 10364 50596 10384
rect 50356 10362 50380 10364
rect 50436 10362 50460 10364
rect 50516 10362 50540 10364
rect 50378 10310 50380 10362
rect 50442 10310 50454 10362
rect 50516 10310 50518 10362
rect 50356 10308 50380 10310
rect 50436 10308 50460 10310
rect 50516 10308 50540 10310
rect 50300 10288 50596 10308
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 50300 9276 50596 9296
rect 50356 9274 50380 9276
rect 50436 9274 50460 9276
rect 50516 9274 50540 9276
rect 50378 9222 50380 9274
rect 50442 9222 50454 9274
rect 50516 9222 50518 9274
rect 50356 9220 50380 9222
rect 50436 9220 50460 9222
rect 50516 9220 50540 9222
rect 50300 9200 50596 9220
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 50300 8188 50596 8208
rect 50356 8186 50380 8188
rect 50436 8186 50460 8188
rect 50516 8186 50540 8188
rect 50378 8134 50380 8186
rect 50442 8134 50454 8186
rect 50516 8134 50518 8186
rect 50356 8132 50380 8134
rect 50436 8132 50460 8134
rect 50516 8132 50540 8134
rect 50300 8112 50596 8132
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34940 7568 35236 7588
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 50300 7100 50596 7120
rect 50356 7098 50380 7100
rect 50436 7098 50460 7100
rect 50516 7098 50540 7100
rect 50378 7046 50380 7098
rect 50442 7046 50454 7098
rect 50516 7046 50518 7098
rect 50356 7044 50380 7046
rect 50436 7044 50460 7046
rect 50516 7044 50540 7046
rect 50300 7024 50596 7044
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 50300 6012 50596 6032
rect 50356 6010 50380 6012
rect 50436 6010 50460 6012
rect 50516 6010 50540 6012
rect 50378 5958 50380 6010
rect 50442 5958 50454 6010
rect 50516 5958 50518 6010
rect 50356 5956 50380 5958
rect 50436 5956 50460 5958
rect 50516 5956 50540 5958
rect 50300 5936 50596 5956
rect 29552 5772 29604 5778
rect 29552 5714 29604 5720
rect 29564 5574 29592 5714
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 28080 2984 28132 2990
rect 28080 2926 28132 2932
rect 29000 2984 29052 2990
rect 29000 2926 29052 2932
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 20720 2508 20772 2514
rect 20720 2450 20772 2456
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 23480 2508 23532 2514
rect 23480 2450 23532 2456
rect 24400 2508 24452 2514
rect 24400 2450 24452 2456
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 27160 2508 27212 2514
rect 27160 2450 27212 2456
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19812 800 19840 2450
rect 20732 800 20760 2450
rect 21652 800 21680 2450
rect 22572 800 22600 2450
rect 23492 800 23520 2450
rect 24412 800 24440 2450
rect 25332 800 25360 2450
rect 26252 800 26280 2450
rect 27172 800 27200 2450
rect 28092 800 28120 2926
rect 29012 800 29040 2926
rect 29104 2514 29132 3334
rect 29564 2990 29592 5510
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 51000 5234 51028 19994
rect 53748 19916 53800 19922
rect 53748 19858 53800 19864
rect 53760 17066 53788 19858
rect 54312 19854 54340 23258
rect 55036 22568 55088 22574
rect 55036 22510 55088 22516
rect 55048 22098 55076 22510
rect 55232 22234 55260 23462
rect 55600 23322 55628 23598
rect 55588 23316 55640 23322
rect 55588 23258 55640 23264
rect 55404 23180 55456 23186
rect 55404 23122 55456 23128
rect 55220 22228 55272 22234
rect 55220 22170 55272 22176
rect 55036 22092 55088 22098
rect 55036 22034 55088 22040
rect 55220 21480 55272 21486
rect 55220 21422 55272 21428
rect 55232 21350 55260 21422
rect 55220 21344 55272 21350
rect 55220 21286 55272 21292
rect 55232 21010 55260 21286
rect 55220 21004 55272 21010
rect 55220 20946 55272 20952
rect 55416 20398 55444 23122
rect 55692 23050 55720 24210
rect 56060 23866 56088 27474
rect 56508 25832 56560 25838
rect 56508 25774 56560 25780
rect 56324 25424 56376 25430
rect 56324 25366 56376 25372
rect 56048 23860 56100 23866
rect 56048 23802 56100 23808
rect 55680 23044 55732 23050
rect 55680 22986 55732 22992
rect 55496 22568 55548 22574
rect 55496 22510 55548 22516
rect 55508 22166 55536 22510
rect 55496 22160 55548 22166
rect 55496 22102 55548 22108
rect 55772 22092 55824 22098
rect 55772 22034 55824 22040
rect 55680 21480 55732 21486
rect 55680 21422 55732 21428
rect 55692 20874 55720 21422
rect 55680 20868 55732 20874
rect 55680 20810 55732 20816
rect 55220 20392 55272 20398
rect 55220 20334 55272 20340
rect 55404 20392 55456 20398
rect 55404 20334 55456 20340
rect 55232 20262 55260 20334
rect 55784 20262 55812 22034
rect 55864 21888 55916 21894
rect 55864 21830 55916 21836
rect 55876 21554 55904 21830
rect 55864 21548 55916 21554
rect 55864 21490 55916 21496
rect 56048 21004 56100 21010
rect 56048 20946 56100 20952
rect 56060 20602 56088 20946
rect 56048 20596 56100 20602
rect 56048 20538 56100 20544
rect 56048 20392 56100 20398
rect 56048 20334 56100 20340
rect 55220 20256 55272 20262
rect 55220 20198 55272 20204
rect 55772 20256 55824 20262
rect 55772 20198 55824 20204
rect 54300 19848 54352 19854
rect 54300 19790 54352 19796
rect 55586 19000 55642 19009
rect 55586 18935 55642 18944
rect 55600 18834 55628 18935
rect 55588 18828 55640 18834
rect 55588 18770 55640 18776
rect 55404 17672 55456 17678
rect 55404 17614 55456 17620
rect 55416 17338 55444 17614
rect 55220 17332 55272 17338
rect 55220 17274 55272 17280
rect 55404 17332 55456 17338
rect 55404 17274 55456 17280
rect 53748 17060 53800 17066
rect 53748 17002 53800 17008
rect 55232 15162 55260 17274
rect 55772 17128 55824 17134
rect 55772 17070 55824 17076
rect 55784 16658 55812 17070
rect 55772 16652 55824 16658
rect 55772 16594 55824 16600
rect 55588 16040 55640 16046
rect 55588 15982 55640 15988
rect 55600 15881 55628 15982
rect 55586 15872 55642 15881
rect 55586 15807 55642 15816
rect 55220 15156 55272 15162
rect 55220 15098 55272 15104
rect 55784 14958 55812 16594
rect 55772 14952 55824 14958
rect 55772 14894 55824 14900
rect 55588 14476 55640 14482
rect 55588 14418 55640 14424
rect 53840 14340 53892 14346
rect 53840 14282 53892 14288
rect 52552 7540 52604 7546
rect 52552 7482 52604 7488
rect 52564 6866 52592 7482
rect 53748 6928 53800 6934
rect 53748 6870 53800 6876
rect 52552 6860 52604 6866
rect 52552 6802 52604 6808
rect 52460 6384 52512 6390
rect 52460 6326 52512 6332
rect 52368 6248 52420 6254
rect 52368 6190 52420 6196
rect 50988 5228 51040 5234
rect 50988 5170 51040 5176
rect 49976 5160 50028 5166
rect 49976 5102 50028 5108
rect 50620 5160 50672 5166
rect 50620 5102 50672 5108
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 49148 4684 49200 4690
rect 49148 4626 49200 4632
rect 33600 4480 33652 4486
rect 33600 4422 33652 4428
rect 36268 4480 36320 4486
rect 36268 4422 36320 4428
rect 37280 4480 37332 4486
rect 37280 4422 37332 4428
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 33048 4072 33100 4078
rect 33048 4014 33100 4020
rect 30024 3058 30052 4014
rect 30656 3596 30708 3602
rect 30656 3538 30708 3544
rect 30196 3392 30248 3398
rect 30196 3334 30248 3340
rect 30208 3058 30236 3334
rect 30668 3126 30696 3538
rect 30932 3392 30984 3398
rect 30932 3334 30984 3340
rect 32128 3392 32180 3398
rect 32128 3334 32180 3340
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 30656 3120 30708 3126
rect 30656 3062 30708 3068
rect 30012 3052 30064 3058
rect 30012 2994 30064 3000
rect 30196 3052 30248 3058
rect 30196 2994 30248 3000
rect 29552 2984 29604 2990
rect 29552 2926 29604 2932
rect 29368 2848 29420 2854
rect 29368 2790 29420 2796
rect 29380 2514 29408 2790
rect 30944 2514 30972 3334
rect 32140 3058 32168 3334
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31944 2916 31996 2922
rect 31944 2858 31996 2864
rect 31116 2848 31168 2854
rect 31116 2790 31168 2796
rect 31128 2514 31156 2790
rect 31772 2582 31800 2858
rect 31852 2848 31904 2854
rect 31852 2790 31904 2796
rect 31760 2576 31812 2582
rect 31760 2518 31812 2524
rect 29092 2508 29144 2514
rect 29092 2450 29144 2456
rect 29368 2508 29420 2514
rect 29368 2450 29420 2456
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 31116 2508 31168 2514
rect 31116 2450 31168 2456
rect 29920 2372 29972 2378
rect 29920 2314 29972 2320
rect 29932 800 29960 2314
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30944 800 30972 2246
rect 31864 800 31892 2790
rect 31956 2650 31984 2858
rect 31944 2644 31996 2650
rect 31944 2586 31996 2592
rect 32784 800 32812 3334
rect 33060 2990 33088 4014
rect 33416 3596 33468 3602
rect 33416 3538 33468 3544
rect 33428 3194 33456 3538
rect 33416 3188 33468 3194
rect 33416 3130 33468 3136
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 33612 2514 33640 4422
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 33784 3936 33836 3942
rect 33784 3878 33836 3884
rect 34520 3936 34572 3942
rect 34520 3878 34572 3884
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33600 2508 33652 2514
rect 33600 2450 33652 2456
rect 33704 800 33732 3334
rect 33796 2514 33824 3878
rect 33968 3596 34020 3602
rect 33968 3538 34020 3544
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 33784 2508 33836 2514
rect 33784 2450 33836 2456
rect 33980 2378 34008 3538
rect 34348 2990 34376 3538
rect 34336 2984 34388 2990
rect 34336 2926 34388 2932
rect 34532 2446 34560 3878
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 3058 34652 3334
rect 34612 3052 34664 3058
rect 34612 2994 34664 3000
rect 34612 2916 34664 2922
rect 34612 2858 34664 2864
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 33968 2372 34020 2378
rect 33968 2314 34020 2320
rect 34624 800 34652 2858
rect 34808 2514 34836 4150
rect 35256 4072 35308 4078
rect 35256 4014 35308 4020
rect 36084 4072 36136 4078
rect 36084 4014 36136 4020
rect 34888 3936 34940 3942
rect 34888 3878 34940 3884
rect 34900 3602 34928 3878
rect 34888 3596 34940 3602
rect 34888 3538 34940 3544
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 35268 2990 35296 4014
rect 36096 3602 36124 4014
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35452 3194 35480 3538
rect 35532 3392 35584 3398
rect 35532 3334 35584 3340
rect 35440 3188 35492 3194
rect 35440 3130 35492 3136
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 34980 2848 35032 2854
rect 34980 2790 35032 2796
rect 34992 2514 35020 2790
rect 34796 2508 34848 2514
rect 34796 2450 34848 2456
rect 34980 2508 35032 2514
rect 34980 2450 35032 2456
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35544 800 35572 3334
rect 35992 2916 36044 2922
rect 35992 2858 36044 2864
rect 36004 2650 36032 2858
rect 35992 2644 36044 2650
rect 35992 2586 36044 2592
rect 36280 2446 36308 4422
rect 36728 2916 36780 2922
rect 36728 2858 36780 2864
rect 36452 2848 36504 2854
rect 36452 2790 36504 2796
rect 36268 2440 36320 2446
rect 36268 2382 36320 2388
rect 36464 800 36492 2790
rect 36740 2650 36768 2858
rect 36728 2644 36780 2650
rect 36728 2586 36780 2592
rect 37292 2514 37320 4422
rect 37384 4078 37412 4626
rect 46940 4548 46992 4554
rect 46940 4490 46992 4496
rect 38384 4480 38436 4486
rect 38384 4422 38436 4428
rect 38568 4480 38620 4486
rect 38568 4422 38620 4428
rect 39396 4480 39448 4486
rect 39396 4422 39448 4428
rect 39488 4480 39540 4486
rect 39488 4422 39540 4428
rect 41512 4480 41564 4486
rect 41512 4422 41564 4428
rect 42340 4480 42392 4486
rect 42340 4422 42392 4428
rect 43444 4480 43496 4486
rect 43444 4422 43496 4428
rect 37372 4072 37424 4078
rect 37372 4014 37424 4020
rect 37384 3738 37412 4014
rect 37556 3936 37608 3942
rect 37556 3878 37608 3884
rect 37372 3732 37424 3738
rect 37372 3674 37424 3680
rect 37372 3392 37424 3398
rect 37372 3334 37424 3340
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37384 800 37412 3334
rect 37568 2514 37596 3878
rect 37740 3596 37792 3602
rect 37740 3538 37792 3544
rect 37556 2508 37608 2514
rect 37556 2450 37608 2456
rect 37752 2378 37780 3538
rect 38292 3392 38344 3398
rect 38292 3334 38344 3340
rect 37740 2372 37792 2378
rect 37740 2314 37792 2320
rect 38304 800 38332 3334
rect 38396 2990 38424 4422
rect 38580 3058 38608 4422
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 39304 3596 39356 3602
rect 39304 3538 39356 3544
rect 38672 3194 38700 3538
rect 39212 3392 39264 3398
rect 39212 3334 39264 3340
rect 38660 3188 38712 3194
rect 38660 3130 38712 3136
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 38384 2984 38436 2990
rect 38384 2926 38436 2932
rect 39224 800 39252 3334
rect 39316 3194 39344 3538
rect 39304 3188 39356 3194
rect 39304 3130 39356 3136
rect 39408 3058 39436 4422
rect 39396 3052 39448 3058
rect 39396 2994 39448 3000
rect 39500 2514 39528 4422
rect 41236 4072 41288 4078
rect 41236 4014 41288 4020
rect 39580 3936 39632 3942
rect 39580 3878 39632 3884
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 40408 3936 40460 3942
rect 40408 3878 40460 3884
rect 39592 3058 39620 3878
rect 39776 3058 39804 3878
rect 40132 3392 40184 3398
rect 40132 3334 40184 3340
rect 39580 3052 39632 3058
rect 39580 2994 39632 3000
rect 39764 3052 39816 3058
rect 39764 2994 39816 3000
rect 39488 2508 39540 2514
rect 39488 2450 39540 2456
rect 40144 800 40172 3334
rect 40420 2514 40448 3878
rect 41052 3596 41104 3602
rect 41052 3538 41104 3544
rect 40960 2848 41012 2854
rect 40960 2790 41012 2796
rect 40408 2508 40460 2514
rect 40408 2450 40460 2456
rect 40972 1442 41000 2790
rect 41064 2650 41092 3538
rect 41248 2990 41276 4014
rect 41236 2984 41288 2990
rect 41236 2926 41288 2932
rect 41052 2644 41104 2650
rect 41052 2586 41104 2592
rect 41524 2514 41552 4422
rect 41880 3936 41932 3942
rect 41880 3878 41932 3884
rect 41892 2514 41920 3878
rect 41972 2848 42024 2854
rect 41972 2790 42024 2796
rect 41512 2508 41564 2514
rect 41512 2450 41564 2456
rect 41880 2508 41932 2514
rect 41880 2450 41932 2456
rect 40972 1414 41092 1442
rect 41064 800 41092 1414
rect 41984 800 42012 2790
rect 42352 2514 42380 4422
rect 42432 4072 42484 4078
rect 42432 4014 42484 4020
rect 42444 3602 42472 4014
rect 42432 3596 42484 3602
rect 42432 3538 42484 3544
rect 43076 3596 43128 3602
rect 43076 3538 43128 3544
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42892 3392 42944 3398
rect 42892 3334 42944 3340
rect 42432 2916 42484 2922
rect 42432 2858 42484 2864
rect 42444 2650 42472 2858
rect 42432 2644 42484 2650
rect 42432 2586 42484 2592
rect 42812 2514 42840 3334
rect 42340 2508 42392 2514
rect 42340 2450 42392 2456
rect 42800 2508 42852 2514
rect 42800 2450 42852 2456
rect 42904 800 42932 3334
rect 43088 2378 43116 3538
rect 43456 3058 43484 4422
rect 44272 4208 44324 4214
rect 44272 4150 44324 4156
rect 45744 4208 45796 4214
rect 45744 4150 45796 4156
rect 43904 4072 43956 4078
rect 43904 4014 43956 4020
rect 43720 3936 43772 3942
rect 43720 3878 43772 3884
rect 43732 3058 43760 3878
rect 43916 3738 43944 4014
rect 43904 3732 43956 3738
rect 43904 3674 43956 3680
rect 43444 3052 43496 3058
rect 43444 2994 43496 3000
rect 43720 3052 43772 3058
rect 43720 2994 43772 3000
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 43076 2372 43128 2378
rect 43076 2314 43128 2320
rect 43824 800 43852 2790
rect 44284 2514 44312 4150
rect 44456 3936 44508 3942
rect 44456 3878 44508 3884
rect 44468 2514 44496 3878
rect 45560 3392 45612 3398
rect 45560 3334 45612 3340
rect 44732 3052 44784 3058
rect 44732 2994 44784 3000
rect 44272 2508 44324 2514
rect 44272 2450 44324 2456
rect 44456 2508 44508 2514
rect 44456 2450 44508 2456
rect 44744 800 44772 2994
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45480 2650 45508 2858
rect 45468 2644 45520 2650
rect 45468 2586 45520 2592
rect 45572 2446 45600 3334
rect 45652 2848 45704 2854
rect 45652 2790 45704 2796
rect 45560 2440 45612 2446
rect 45560 2382 45612 2388
rect 45664 800 45692 2790
rect 45756 2514 45784 4150
rect 46204 2916 46256 2922
rect 46204 2858 46256 2864
rect 46216 2650 46244 2858
rect 46204 2644 46256 2650
rect 46204 2586 46256 2592
rect 46952 2514 46980 4490
rect 47032 4480 47084 4486
rect 47032 4422 47084 4428
rect 48044 4480 48096 4486
rect 48044 4422 48096 4428
rect 48964 4480 49016 4486
rect 48964 4422 49016 4428
rect 49056 4480 49108 4486
rect 49056 4422 49108 4428
rect 47044 2990 47072 4422
rect 47676 4072 47728 4078
rect 47676 4014 47728 4020
rect 47216 4004 47268 4010
rect 47216 3946 47268 3952
rect 47124 3936 47176 3942
rect 47124 3878 47176 3884
rect 47136 3058 47164 3878
rect 47228 3602 47256 3946
rect 47216 3596 47268 3602
rect 47216 3538 47268 3544
rect 47584 3596 47636 3602
rect 47584 3538 47636 3544
rect 47216 3460 47268 3466
rect 47216 3402 47268 3408
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 47032 2984 47084 2990
rect 47032 2926 47084 2932
rect 47228 2514 47256 3402
rect 47400 3392 47452 3398
rect 47400 3334 47452 3340
rect 47492 3392 47544 3398
rect 47492 3334 47544 3340
rect 45744 2508 45796 2514
rect 45744 2450 45796 2456
rect 46940 2508 46992 2514
rect 46940 2450 46992 2456
rect 47216 2508 47268 2514
rect 47216 2450 47268 2456
rect 47412 2446 47440 3334
rect 47400 2440 47452 2446
rect 47400 2382 47452 2388
rect 46572 2304 46624 2310
rect 46572 2246 46624 2252
rect 46584 800 46612 2246
rect 47504 800 47532 3334
rect 47596 3194 47624 3538
rect 47688 3534 47716 4014
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 47584 3188 47636 3194
rect 47584 3130 47636 3136
rect 48056 2514 48084 4422
rect 48504 3596 48556 3602
rect 48504 3538 48556 3544
rect 48412 3392 48464 3398
rect 48412 3334 48464 3340
rect 48044 2508 48096 2514
rect 48044 2450 48096 2456
rect 48424 800 48452 3334
rect 48516 2650 48544 3538
rect 48976 3058 49004 4422
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 49068 2990 49096 4422
rect 49160 4078 49188 4626
rect 49700 4480 49752 4486
rect 49700 4422 49752 4428
rect 49148 4072 49200 4078
rect 49148 4014 49200 4020
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 49620 3126 49648 3334
rect 49608 3120 49660 3126
rect 49608 3062 49660 3068
rect 49056 2984 49108 2990
rect 49056 2926 49108 2932
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 48504 2644 48556 2650
rect 48504 2586 48556 2592
rect 49344 800 49372 2790
rect 49712 2446 49740 4422
rect 49792 4072 49844 4078
rect 49792 4014 49844 4020
rect 49804 2514 49832 4014
rect 49884 3936 49936 3942
rect 49884 3878 49936 3884
rect 49896 3602 49924 3878
rect 49884 3596 49936 3602
rect 49884 3538 49936 3544
rect 49792 2508 49844 2514
rect 49792 2450 49844 2456
rect 49700 2440 49752 2446
rect 49700 2382 49752 2388
rect 49988 1766 50016 5102
rect 50300 4924 50596 4944
rect 50356 4922 50380 4924
rect 50436 4922 50460 4924
rect 50516 4922 50540 4924
rect 50378 4870 50380 4922
rect 50442 4870 50454 4922
rect 50516 4870 50518 4922
rect 50356 4868 50380 4870
rect 50436 4868 50460 4870
rect 50516 4868 50540 4870
rect 50300 4848 50596 4868
rect 50300 3836 50596 3856
rect 50356 3834 50380 3836
rect 50436 3834 50460 3836
rect 50516 3834 50540 3836
rect 50378 3782 50380 3834
rect 50442 3782 50454 3834
rect 50516 3782 50518 3834
rect 50356 3780 50380 3782
rect 50436 3780 50460 3782
rect 50516 3780 50540 3782
rect 50300 3760 50596 3780
rect 50160 3596 50212 3602
rect 50160 3538 50212 3544
rect 50068 3392 50120 3398
rect 50068 3334 50120 3340
rect 49976 1760 50028 1766
rect 49976 1702 50028 1708
rect 50080 1714 50108 3334
rect 50172 2650 50200 3538
rect 50632 3058 50660 5102
rect 51000 4078 51028 5170
rect 51632 5160 51684 5166
rect 51632 5102 51684 5108
rect 50988 4072 51040 4078
rect 50988 4014 51040 4020
rect 51540 3936 51592 3942
rect 51540 3878 51592 3884
rect 51448 3596 51500 3602
rect 51448 3538 51500 3544
rect 51172 3392 51224 3398
rect 51172 3334 51224 3340
rect 50620 3052 50672 3058
rect 50620 2994 50672 3000
rect 50300 2748 50596 2768
rect 50356 2746 50380 2748
rect 50436 2746 50460 2748
rect 50516 2746 50540 2748
rect 50378 2694 50380 2746
rect 50442 2694 50454 2746
rect 50516 2694 50518 2746
rect 50356 2692 50380 2694
rect 50436 2692 50460 2694
rect 50516 2692 50540 2694
rect 50300 2672 50596 2692
rect 50160 2644 50212 2650
rect 50160 2586 50212 2592
rect 50080 1686 50292 1714
rect 50264 800 50292 1686
rect 51184 800 51212 3334
rect 51460 3194 51488 3538
rect 51448 3188 51500 3194
rect 51448 3130 51500 3136
rect 51552 2446 51580 3878
rect 51644 2514 51672 5102
rect 51908 5092 51960 5098
rect 51908 5034 51960 5040
rect 51920 4690 51948 5034
rect 51908 4684 51960 4690
rect 51908 4626 51960 4632
rect 51724 4480 51776 4486
rect 51724 4422 51776 4428
rect 51736 2990 51764 4422
rect 51920 4078 51948 4626
rect 51908 4072 51960 4078
rect 51908 4014 51960 4020
rect 52000 3936 52052 3942
rect 52000 3878 52052 3884
rect 52012 3126 52040 3878
rect 52092 3392 52144 3398
rect 52092 3334 52144 3340
rect 52000 3120 52052 3126
rect 52000 3062 52052 3068
rect 51724 2984 51776 2990
rect 51724 2926 51776 2932
rect 51632 2508 51684 2514
rect 51632 2450 51684 2456
rect 51540 2440 51592 2446
rect 51540 2382 51592 2388
rect 52104 800 52132 3334
rect 52380 814 52408 6190
rect 52472 5778 52500 6326
rect 53760 5778 53788 6870
rect 52460 5772 52512 5778
rect 52460 5714 52512 5720
rect 53748 5772 53800 5778
rect 53748 5714 53800 5720
rect 53104 5568 53156 5574
rect 53104 5510 53156 5516
rect 52460 5160 52512 5166
rect 52460 5102 52512 5108
rect 52472 3058 52500 5102
rect 52828 3936 52880 3942
rect 52828 3878 52880 3884
rect 52644 3596 52696 3602
rect 52644 3538 52696 3544
rect 52460 3052 52512 3058
rect 52460 2994 52512 3000
rect 52656 2378 52684 3538
rect 52840 2446 52868 3878
rect 53116 3602 53144 5510
rect 53196 5364 53248 5370
rect 53196 5306 53248 5312
rect 53208 4690 53236 5306
rect 53288 5024 53340 5030
rect 53288 4966 53340 4972
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 53208 4078 53236 4626
rect 53196 4072 53248 4078
rect 53196 4014 53248 4020
rect 53300 3602 53328 4966
rect 53748 4480 53800 4486
rect 53748 4422 53800 4428
rect 53104 3596 53156 3602
rect 53104 3538 53156 3544
rect 53288 3596 53340 3602
rect 53288 3538 53340 3544
rect 53012 3392 53064 3398
rect 53012 3334 53064 3340
rect 52828 2440 52880 2446
rect 52828 2382 52880 2388
rect 52644 2372 52696 2378
rect 52644 2314 52696 2320
rect 52368 808 52420 814
rect 2870 504 2926 513
rect 2870 439 2926 448
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 13358 0 13414 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17958 0 18014 800
rect 18878 0 18934 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22558 0 22614 800
rect 23478 0 23534 800
rect 24398 0 24454 800
rect 25318 0 25374 800
rect 26238 0 26294 800
rect 27158 0 27214 800
rect 28078 0 28134 800
rect 28998 0 29054 800
rect 29918 0 29974 800
rect 30930 0 30986 800
rect 31850 0 31906 800
rect 32770 0 32826 800
rect 33690 0 33746 800
rect 34610 0 34666 800
rect 35530 0 35586 800
rect 36450 0 36506 800
rect 37370 0 37426 800
rect 38290 0 38346 800
rect 39210 0 39266 800
rect 40130 0 40186 800
rect 41050 0 41106 800
rect 41970 0 42026 800
rect 42890 0 42946 800
rect 43810 0 43866 800
rect 44730 0 44786 800
rect 45650 0 45706 800
rect 46570 0 46626 800
rect 47490 0 47546 800
rect 48410 0 48466 800
rect 49330 0 49386 800
rect 50250 0 50306 800
rect 51170 0 51226 800
rect 52090 0 52146 800
rect 53024 800 53052 3334
rect 53760 2990 53788 4422
rect 53748 2984 53800 2990
rect 53748 2926 53800 2932
rect 53852 2582 53880 14282
rect 55600 14249 55628 14418
rect 55772 14408 55824 14414
rect 55772 14350 55824 14356
rect 55586 14240 55642 14249
rect 55586 14175 55642 14184
rect 55784 14074 55812 14350
rect 55772 14068 55824 14074
rect 55772 14010 55824 14016
rect 56060 12782 56088 20334
rect 56140 20256 56192 20262
rect 56140 20198 56192 20204
rect 56152 19310 56180 20198
rect 56140 19304 56192 19310
rect 56140 19246 56192 19252
rect 56232 18216 56284 18222
rect 56232 18158 56284 18164
rect 56244 17377 56272 18158
rect 56230 17368 56286 17377
rect 56230 17303 56286 17312
rect 56336 17270 56364 25366
rect 56520 25265 56548 25774
rect 56506 25256 56562 25265
rect 56506 25191 56562 25200
rect 56508 23656 56560 23662
rect 56506 23624 56508 23633
rect 56560 23624 56562 23633
rect 56506 23559 56562 23568
rect 56416 22568 56468 22574
rect 56416 22510 56468 22516
rect 56428 21690 56456 22510
rect 56416 21684 56468 21690
rect 56416 21626 56468 21632
rect 56506 20496 56562 20505
rect 56506 20431 56562 20440
rect 56520 20330 56548 20431
rect 56508 20324 56560 20330
rect 56508 20266 56560 20272
rect 56324 17264 56376 17270
rect 56324 17206 56376 17212
rect 56336 16046 56364 17206
rect 56612 16250 56640 55186
rect 56692 55150 56744 55156
rect 56966 53816 57022 53825
rect 56966 53751 56968 53760
rect 57020 53751 57022 53760
rect 56968 53722 57020 53728
rect 57058 49192 57114 49201
rect 57058 49127 57060 49136
rect 57112 49127 57114 49136
rect 57060 49098 57112 49104
rect 56874 47152 56930 47161
rect 56874 47087 56876 47096
rect 56928 47087 56930 47096
rect 56876 47058 56928 47064
rect 56968 44940 57020 44946
rect 56968 44882 57020 44888
rect 56876 42764 56928 42770
rect 56876 42706 56928 42712
rect 56784 37324 56836 37330
rect 56784 37266 56836 37272
rect 56796 33590 56824 37266
rect 56784 33584 56836 33590
rect 56784 33526 56836 33532
rect 56784 33380 56836 33386
rect 56784 33322 56836 33328
rect 56692 31884 56744 31890
rect 56692 31826 56744 31832
rect 56704 26586 56732 31826
rect 56796 30172 56824 33322
rect 56888 31346 56916 42706
rect 56980 37330 57008 44882
rect 57058 42936 57114 42945
rect 57058 42871 57114 42880
rect 57072 42770 57100 42871
rect 57060 42764 57112 42770
rect 57060 42706 57112 42712
rect 57060 41676 57112 41682
rect 57060 41618 57112 41624
rect 57072 40594 57100 41618
rect 57060 40588 57112 40594
rect 57060 40530 57112 40536
rect 56968 37324 57020 37330
rect 56968 37266 57020 37272
rect 57058 36680 57114 36689
rect 57058 36615 57060 36624
rect 57112 36615 57114 36624
rect 57060 36586 57112 36592
rect 56968 36576 57020 36582
rect 56968 36518 57020 36524
rect 56980 33658 57008 36518
rect 57060 34468 57112 34474
rect 57060 34410 57112 34416
rect 57072 34066 57100 34410
rect 57060 34060 57112 34066
rect 57060 34002 57112 34008
rect 56968 33652 57020 33658
rect 56968 33594 57020 33600
rect 57058 33552 57114 33561
rect 57058 33487 57060 33496
rect 57112 33487 57114 33496
rect 57060 33458 57112 33464
rect 57164 32434 57192 56850
rect 57256 55894 57284 57310
rect 57980 57316 58032 57322
rect 57980 57258 58032 57264
rect 57992 57050 58020 57258
rect 57980 57044 58032 57050
rect 57980 56986 58032 56992
rect 58084 56438 58112 57446
rect 58162 57423 58164 57432
rect 58216 57423 58218 57432
rect 58164 57394 58216 57400
rect 58348 57248 58400 57254
rect 58348 57190 58400 57196
rect 58072 56432 58124 56438
rect 58072 56374 58124 56380
rect 58162 55992 58218 56001
rect 58162 55927 58218 55936
rect 57244 55888 57296 55894
rect 57244 55830 57296 55836
rect 57704 55752 57756 55758
rect 57704 55694 57756 55700
rect 57334 55448 57390 55457
rect 57334 55383 57336 55392
rect 57388 55383 57390 55392
rect 57336 55354 57388 55360
rect 57716 55350 57744 55694
rect 57980 55616 58032 55622
rect 57980 55558 58032 55564
rect 57704 55344 57756 55350
rect 57704 55286 57756 55292
rect 57992 55214 58020 55558
rect 58176 55350 58204 55927
rect 58164 55344 58216 55350
rect 58164 55286 58216 55292
rect 57980 55208 58032 55214
rect 57980 55150 58032 55156
rect 58360 54874 58388 57190
rect 58728 56166 58756 59200
rect 59556 56506 59584 59200
rect 59544 56500 59596 56506
rect 59544 56442 59596 56448
rect 58716 56160 58768 56166
rect 58716 56102 58768 56108
rect 58532 55140 58584 55146
rect 58532 55082 58584 55088
rect 58348 54868 58400 54874
rect 58348 54810 58400 54816
rect 57704 54664 57756 54670
rect 57704 54606 57756 54612
rect 57716 54330 57744 54606
rect 58162 54360 58218 54369
rect 57704 54324 57756 54330
rect 58162 54295 58218 54304
rect 57704 54266 57756 54272
rect 58176 54262 58204 54295
rect 58164 54256 58216 54262
rect 58164 54198 58216 54204
rect 57336 54120 57388 54126
rect 57336 54062 57388 54068
rect 57428 54120 57480 54126
rect 57428 54062 57480 54068
rect 57348 53650 57376 54062
rect 57336 53644 57388 53650
rect 57336 53586 57388 53592
rect 57440 51354 57468 54062
rect 57980 54052 58032 54058
rect 57980 53994 58032 54000
rect 57992 53786 58020 53994
rect 57980 53780 58032 53786
rect 57980 53722 58032 53728
rect 57796 53712 57848 53718
rect 57796 53654 57848 53660
rect 57704 53576 57756 53582
rect 57704 53518 57756 53524
rect 57716 53242 57744 53518
rect 57704 53236 57756 53242
rect 57704 53178 57756 53184
rect 57520 53032 57572 53038
rect 57520 52974 57572 52980
rect 57532 51950 57560 52974
rect 57704 52488 57756 52494
rect 57704 52430 57756 52436
rect 57716 52154 57744 52430
rect 57704 52148 57756 52154
rect 57704 52090 57756 52096
rect 57520 51944 57572 51950
rect 57520 51886 57572 51892
rect 57348 51326 57468 51354
rect 57244 50380 57296 50386
rect 57244 50322 57296 50328
rect 57256 50289 57284 50322
rect 57242 50280 57298 50289
rect 57242 50215 57298 50224
rect 57244 49632 57296 49638
rect 57244 49574 57296 49580
rect 57256 49298 57284 49574
rect 57244 49292 57296 49298
rect 57244 49234 57296 49240
rect 57348 45554 57376 51326
rect 57428 51264 57480 51270
rect 57428 51206 57480 51212
rect 57440 50930 57468 51206
rect 57428 50924 57480 50930
rect 57428 50866 57480 50872
rect 57532 50794 57560 51886
rect 57520 50788 57572 50794
rect 57520 50730 57572 50736
rect 57532 49774 57560 50730
rect 57520 49768 57572 49774
rect 57520 49710 57572 49716
rect 57428 49224 57480 49230
rect 57428 49166 57480 49172
rect 57440 48890 57468 49166
rect 57428 48884 57480 48890
rect 57428 48826 57480 48832
rect 57532 47598 57560 49710
rect 57704 48136 57756 48142
rect 57704 48078 57756 48084
rect 57716 47802 57744 48078
rect 57704 47796 57756 47802
rect 57704 47738 57756 47744
rect 57520 47592 57572 47598
rect 57520 47534 57572 47540
rect 57704 47592 57756 47598
rect 57704 47534 57756 47540
rect 57716 47258 57744 47534
rect 57704 47252 57756 47258
rect 57704 47194 57756 47200
rect 57612 47116 57664 47122
rect 57612 47058 57664 47064
rect 57256 45526 57376 45554
rect 57256 41414 57284 45526
rect 57336 45416 57388 45422
rect 57336 45358 57388 45364
rect 57348 44742 57376 45358
rect 57624 44946 57652 47058
rect 57704 45960 57756 45966
rect 57704 45902 57756 45908
rect 57716 45626 57744 45902
rect 57704 45620 57756 45626
rect 57704 45562 57756 45568
rect 57612 44940 57664 44946
rect 57612 44882 57664 44888
rect 57336 44736 57388 44742
rect 57336 44678 57388 44684
rect 57348 44334 57376 44678
rect 57336 44328 57388 44334
rect 57336 44270 57388 44276
rect 57348 43246 57376 44270
rect 57428 43648 57480 43654
rect 57428 43590 57480 43596
rect 57336 43240 57388 43246
rect 57336 43182 57388 43188
rect 57348 41682 57376 43182
rect 57440 42770 57468 43590
rect 57704 43104 57756 43110
rect 57704 43046 57756 43052
rect 57716 42770 57744 43046
rect 57428 42764 57480 42770
rect 57428 42706 57480 42712
rect 57704 42764 57756 42770
rect 57704 42706 57756 42712
rect 57520 42152 57572 42158
rect 57520 42094 57572 42100
rect 57532 41682 57560 42094
rect 57336 41676 57388 41682
rect 57336 41618 57388 41624
rect 57520 41676 57572 41682
rect 57520 41618 57572 41624
rect 57256 41386 57652 41414
rect 57334 41304 57390 41313
rect 57334 41239 57336 41248
rect 57388 41239 57390 41248
rect 57336 41210 57388 41216
rect 57520 40996 57572 41002
rect 57520 40938 57572 40944
rect 57428 40520 57480 40526
rect 57428 40462 57480 40468
rect 57440 40186 57468 40462
rect 57428 40180 57480 40186
rect 57428 40122 57480 40128
rect 57428 37800 57480 37806
rect 57428 37742 57480 37748
rect 57440 37126 57468 37742
rect 57428 37120 57480 37126
rect 57428 37062 57480 37068
rect 57440 36242 57468 37062
rect 57428 36236 57480 36242
rect 57428 36178 57480 36184
rect 57440 35154 57468 36178
rect 57532 35154 57560 40938
rect 57428 35148 57480 35154
rect 57428 35090 57480 35096
rect 57520 35148 57572 35154
rect 57520 35090 57572 35096
rect 57440 34542 57468 35090
rect 57520 34604 57572 34610
rect 57520 34546 57572 34552
rect 57336 34536 57388 34542
rect 57336 34478 57388 34484
rect 57428 34536 57480 34542
rect 57428 34478 57480 34484
rect 57244 34400 57296 34406
rect 57244 34342 57296 34348
rect 57256 33522 57284 34342
rect 57244 33516 57296 33522
rect 57244 33458 57296 33464
rect 57348 33454 57376 34478
rect 57532 34066 57560 34546
rect 57520 34060 57572 34066
rect 57520 34002 57572 34008
rect 57624 33946 57652 41386
rect 57704 38344 57756 38350
rect 57704 38286 57756 38292
rect 57716 38010 57744 38286
rect 57704 38004 57756 38010
rect 57704 37946 57756 37952
rect 57704 36712 57756 36718
rect 57704 36654 57756 36660
rect 57716 36378 57744 36654
rect 57704 36372 57756 36378
rect 57704 36314 57756 36320
rect 57704 35624 57756 35630
rect 57704 35566 57756 35572
rect 57716 35290 57744 35566
rect 57704 35284 57756 35290
rect 57704 35226 57756 35232
rect 57704 35148 57756 35154
rect 57704 35090 57756 35096
rect 57440 33918 57652 33946
rect 57336 33448 57388 33454
rect 57336 33390 57388 33396
rect 57152 32428 57204 32434
rect 57152 32370 57204 32376
rect 56966 31920 57022 31929
rect 56966 31855 56968 31864
rect 57020 31855 57022 31864
rect 56968 31826 57020 31832
rect 57440 31754 57468 33918
rect 57716 33810 57744 35090
rect 57348 31726 57468 31754
rect 57532 33782 57744 33810
rect 56876 31340 56928 31346
rect 56876 31282 56928 31288
rect 57244 31204 57296 31210
rect 57244 31146 57296 31152
rect 56876 31136 56928 31142
rect 56876 31078 56928 31084
rect 56888 30326 56916 31078
rect 57058 30968 57114 30977
rect 57058 30903 57114 30912
rect 56968 30728 57020 30734
rect 56968 30670 57020 30676
rect 56980 30598 57008 30670
rect 56968 30592 57020 30598
rect 56968 30534 57020 30540
rect 56876 30320 56928 30326
rect 56876 30262 56928 30268
rect 56796 30144 56916 30172
rect 56784 28552 56836 28558
rect 56784 28494 56836 28500
rect 56796 28082 56824 28494
rect 56784 28076 56836 28082
rect 56784 28018 56836 28024
rect 56784 27464 56836 27470
rect 56784 27406 56836 27412
rect 56796 27130 56824 27406
rect 56784 27124 56836 27130
rect 56784 27066 56836 27072
rect 56888 26994 56916 30144
rect 56980 28665 57008 30534
rect 57072 30326 57100 30903
rect 57256 30666 57284 31146
rect 57244 30660 57296 30666
rect 57244 30602 57296 30608
rect 57348 30546 57376 31726
rect 57256 30518 57376 30546
rect 57150 30424 57206 30433
rect 57150 30359 57206 30368
rect 57060 30320 57112 30326
rect 57060 30262 57112 30268
rect 57164 29238 57192 30359
rect 57152 29232 57204 29238
rect 57152 29174 57204 29180
rect 56966 28656 57022 28665
rect 56966 28591 57022 28600
rect 56968 27328 57020 27334
rect 56966 27296 56968 27305
rect 57020 27296 57022 27305
rect 56966 27231 57022 27240
rect 56876 26988 56928 26994
rect 56876 26930 56928 26936
rect 56692 26580 56744 26586
rect 56692 26522 56744 26528
rect 56876 25832 56928 25838
rect 56876 25774 56928 25780
rect 56888 21486 56916 25774
rect 57060 25696 57112 25702
rect 57060 25638 57112 25644
rect 57072 24750 57100 25638
rect 57256 25158 57284 30518
rect 57532 30054 57560 33782
rect 57704 33652 57756 33658
rect 57704 33594 57756 33600
rect 57612 33584 57664 33590
rect 57612 33526 57664 33532
rect 57520 30048 57572 30054
rect 57520 29990 57572 29996
rect 57428 29096 57480 29102
rect 57428 29038 57480 29044
rect 57336 29028 57388 29034
rect 57336 28970 57388 28976
rect 57244 25152 57296 25158
rect 57244 25094 57296 25100
rect 57060 24744 57112 24750
rect 57060 24686 57112 24692
rect 57058 22536 57114 22545
rect 57058 22471 57060 22480
rect 57112 22471 57114 22480
rect 57060 22442 57112 22448
rect 56876 21480 56928 21486
rect 56876 21422 56928 21428
rect 56888 20602 56916 21422
rect 56876 20596 56928 20602
rect 56876 20538 56928 20544
rect 56968 20392 57020 20398
rect 56968 20334 57020 20340
rect 56784 20324 56836 20330
rect 56784 20266 56836 20272
rect 56796 19990 56824 20266
rect 56784 19984 56836 19990
rect 56784 19926 56836 19932
rect 56692 19848 56744 19854
rect 56692 19790 56744 19796
rect 56876 19848 56928 19854
rect 56876 19790 56928 19796
rect 56704 18902 56732 19790
rect 56888 19174 56916 19790
rect 56980 19514 57008 20334
rect 56968 19508 57020 19514
rect 56968 19450 57020 19456
rect 56876 19168 56928 19174
rect 56876 19110 56928 19116
rect 56692 18896 56744 18902
rect 56692 18838 56744 18844
rect 57060 18216 57112 18222
rect 57060 18158 57112 18164
rect 57072 17134 57100 18158
rect 57060 17128 57112 17134
rect 57060 17070 57112 17076
rect 57256 16574 57284 25094
rect 57348 24682 57376 28970
rect 57440 28014 57468 29038
rect 57428 28008 57480 28014
rect 57428 27950 57480 27956
rect 57440 26926 57468 27950
rect 57428 26920 57480 26926
rect 57428 26862 57480 26868
rect 57440 25702 57468 26862
rect 57624 25838 57652 33526
rect 57716 29782 57744 33594
rect 57808 30870 57836 53654
rect 57980 52964 58032 52970
rect 57980 52906 58032 52912
rect 58164 52964 58216 52970
rect 58164 52906 58216 52912
rect 57992 52698 58020 52906
rect 58176 52873 58204 52906
rect 58162 52864 58218 52873
rect 58162 52799 58218 52808
rect 57980 52692 58032 52698
rect 57980 52634 58032 52640
rect 58162 52320 58218 52329
rect 58162 52255 58218 52264
rect 58176 52086 58204 52255
rect 58164 52080 58216 52086
rect 58164 52022 58216 52028
rect 58348 51876 58400 51882
rect 58348 51818 58400 51824
rect 57980 51468 58032 51474
rect 57980 51410 58032 51416
rect 57992 51066 58020 51410
rect 58164 51332 58216 51338
rect 58164 51274 58216 51280
rect 58176 51241 58204 51274
rect 58162 51232 58218 51241
rect 58162 51167 58218 51176
rect 57980 51060 58032 51066
rect 57980 51002 58032 51008
rect 58162 50688 58218 50697
rect 58162 50623 58218 50632
rect 58176 50454 58204 50623
rect 58164 50448 58216 50454
rect 58164 50390 58216 50396
rect 58256 50380 58308 50386
rect 58256 50322 58308 50328
rect 58164 49768 58216 49774
rect 58162 49736 58164 49745
rect 58216 49736 58218 49745
rect 57980 49700 58032 49706
rect 58162 49671 58218 49680
rect 57980 49642 58032 49648
rect 57992 49434 58020 49642
rect 57980 49428 58032 49434
rect 57980 49370 58032 49376
rect 57980 48612 58032 48618
rect 57980 48554 58032 48560
rect 57888 48544 57940 48550
rect 57888 48486 57940 48492
rect 57900 48113 57928 48486
rect 57992 48346 58020 48554
rect 57980 48340 58032 48346
rect 57980 48282 58032 48288
rect 57886 48104 57942 48113
rect 57886 48039 57942 48048
rect 58162 47560 58218 47569
rect 58162 47495 58164 47504
rect 58216 47495 58218 47504
rect 58164 47466 58216 47472
rect 58162 46608 58218 46617
rect 58162 46543 58164 46552
rect 58216 46543 58218 46552
rect 58164 46514 58216 46520
rect 57980 46436 58032 46442
rect 57980 46378 58032 46384
rect 57992 46170 58020 46378
rect 57980 46164 58032 46170
rect 57980 46106 58032 46112
rect 58162 46064 58218 46073
rect 58162 45999 58218 46008
rect 58176 45558 58204 45999
rect 58164 45552 58216 45558
rect 58164 45494 58216 45500
rect 58162 44976 58218 44985
rect 57980 44940 58032 44946
rect 58162 44911 58164 44920
rect 57980 44882 58032 44888
rect 58216 44911 58218 44920
rect 58164 44882 58216 44888
rect 57992 44538 58020 44882
rect 57980 44532 58032 44538
rect 57980 44474 58032 44480
rect 58162 44432 58218 44441
rect 58162 44367 58218 44376
rect 58176 43926 58204 44367
rect 58164 43920 58216 43926
rect 58164 43862 58216 43868
rect 58162 43480 58218 43489
rect 58162 43415 58218 43424
rect 58176 43382 58204 43415
rect 58164 43376 58216 43382
rect 58164 43318 58216 43324
rect 57980 43172 58032 43178
rect 57980 43114 58032 43120
rect 57992 42906 58020 43114
rect 57980 42900 58032 42906
rect 57980 42842 58032 42848
rect 57980 42084 58032 42090
rect 57980 42026 58032 42032
rect 58164 42084 58216 42090
rect 58164 42026 58216 42032
rect 57992 41818 58020 42026
rect 58176 41857 58204 42026
rect 58162 41848 58218 41857
rect 57980 41812 58032 41818
rect 58162 41783 58218 41792
rect 57980 41754 58032 41760
rect 57980 40996 58032 41002
rect 57980 40938 58032 40944
rect 58164 40996 58216 41002
rect 58164 40938 58216 40944
rect 57992 40730 58020 40938
rect 57980 40724 58032 40730
rect 57980 40666 58032 40672
rect 58176 40361 58204 40938
rect 58162 40352 58218 40361
rect 58162 40287 58218 40296
rect 58164 39908 58216 39914
rect 58164 39850 58216 39856
rect 58176 39817 58204 39850
rect 58162 39808 58218 39817
rect 58162 39743 58218 39752
rect 57980 39500 58032 39506
rect 57980 39442 58032 39448
rect 57992 39273 58020 39442
rect 57978 39264 58034 39273
rect 57978 39199 58034 39208
rect 57980 38820 58032 38826
rect 57980 38762 58032 38768
rect 58164 38820 58216 38826
rect 58164 38762 58216 38768
rect 57992 38554 58020 38762
rect 58176 38729 58204 38762
rect 58162 38720 58218 38729
rect 58162 38655 58218 38664
rect 57980 38548 58032 38554
rect 57980 38490 58032 38496
rect 58162 38176 58218 38185
rect 58162 38111 58218 38120
rect 58176 37942 58204 38111
rect 58164 37936 58216 37942
rect 58164 37878 58216 37884
rect 57888 37460 57940 37466
rect 57888 37402 57940 37408
rect 57900 37233 57928 37402
rect 57980 37324 58032 37330
rect 57980 37266 58032 37272
rect 57886 37224 57942 37233
rect 57886 37159 57942 37168
rect 57992 36922 58020 37266
rect 57980 36916 58032 36922
rect 57980 36858 58032 36864
rect 57980 36236 58032 36242
rect 57980 36178 58032 36184
rect 57888 36032 57940 36038
rect 57888 35974 57940 35980
rect 57900 35601 57928 35974
rect 57992 35834 58020 36178
rect 57980 35828 58032 35834
rect 57980 35770 58032 35776
rect 57886 35592 57942 35601
rect 57886 35527 57942 35536
rect 58072 35148 58124 35154
rect 58072 35090 58124 35096
rect 57888 34536 57940 34542
rect 57888 34478 57940 34484
rect 57900 34105 57928 34478
rect 57980 34468 58032 34474
rect 57980 34410 58032 34416
rect 57992 34202 58020 34410
rect 57980 34196 58032 34202
rect 57980 34138 58032 34144
rect 57886 34096 57942 34105
rect 57886 34031 57942 34040
rect 57888 31816 57940 31822
rect 57888 31758 57940 31764
rect 57796 30864 57848 30870
rect 57796 30806 57848 30812
rect 57704 29776 57756 29782
rect 57704 29718 57756 29724
rect 57704 29096 57756 29102
rect 57704 29038 57756 29044
rect 57716 28218 57744 29038
rect 57900 28529 57928 31758
rect 57980 29708 58032 29714
rect 57980 29650 58032 29656
rect 57992 29306 58020 29650
rect 57980 29300 58032 29306
rect 57980 29242 58032 29248
rect 58084 28762 58112 35090
rect 58162 35048 58218 35057
rect 58162 34983 58164 34992
rect 58216 34983 58218 34992
rect 58164 34954 58216 34960
rect 58164 33312 58216 33318
rect 58164 33254 58216 33260
rect 58176 32366 58204 33254
rect 58268 33046 58296 50322
rect 58256 33040 58308 33046
rect 58256 32982 58308 32988
rect 58164 32360 58216 32366
rect 58164 32302 58216 32308
rect 58360 31958 58388 51818
rect 58544 41414 58572 55082
rect 58808 45348 58860 45354
rect 58808 45290 58860 45296
rect 58452 41386 58572 41414
rect 58348 31952 58400 31958
rect 58348 31894 58400 31900
rect 58452 31346 58480 41386
rect 58624 39976 58676 39982
rect 58624 39918 58676 39924
rect 58532 32496 58584 32502
rect 58530 32464 58532 32473
rect 58584 32464 58586 32473
rect 58530 32399 58586 32408
rect 58440 31340 58492 31346
rect 58440 31282 58492 31288
rect 58636 29850 58664 39918
rect 58716 37732 58768 37738
rect 58716 37674 58768 37680
rect 58624 29844 58676 29850
rect 58624 29786 58676 29792
rect 58164 29572 58216 29578
rect 58164 29514 58216 29520
rect 58176 29345 58204 29514
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 58162 28792 58218 28801
rect 58072 28756 58124 28762
rect 58162 28727 58218 28736
rect 58072 28698 58124 28704
rect 58176 28694 58204 28727
rect 58164 28688 58216 28694
rect 58164 28630 58216 28636
rect 58072 28620 58124 28626
rect 58072 28562 58124 28568
rect 57886 28520 57942 28529
rect 57886 28455 57942 28464
rect 57704 28212 57756 28218
rect 57704 28154 57756 28160
rect 57980 27940 58032 27946
rect 57980 27882 58032 27888
rect 57992 27674 58020 27882
rect 57980 27668 58032 27674
rect 57980 27610 58032 27616
rect 57704 27464 57756 27470
rect 57704 27406 57756 27412
rect 57716 27130 57744 27406
rect 57704 27124 57756 27130
rect 57704 27066 57756 27072
rect 57980 26852 58032 26858
rect 57980 26794 58032 26800
rect 57992 26586 58020 26794
rect 57980 26580 58032 26586
rect 57980 26522 58032 26528
rect 57980 26376 58032 26382
rect 57980 26318 58032 26324
rect 57612 25832 57664 25838
rect 57612 25774 57664 25780
rect 57428 25696 57480 25702
rect 57428 25638 57480 25644
rect 57440 25362 57468 25638
rect 57992 25498 58020 26318
rect 57980 25492 58032 25498
rect 57980 25434 58032 25440
rect 57428 25356 57480 25362
rect 57428 25298 57480 25304
rect 58084 24818 58112 28562
rect 58728 28558 58756 37674
rect 58820 33386 58848 45290
rect 58808 33380 58860 33386
rect 58808 33322 58860 33328
rect 58716 28552 58768 28558
rect 58716 28494 58768 28500
rect 58164 27940 58216 27946
rect 58164 27882 58216 27888
rect 58176 27849 58204 27882
rect 58162 27840 58218 27849
rect 58162 27775 58218 27784
rect 58348 26784 58400 26790
rect 58348 26726 58400 26732
rect 58360 26217 58388 26726
rect 58346 26208 58402 26217
rect 58346 26143 58402 26152
rect 58256 25832 58308 25838
rect 58256 25774 58308 25780
rect 58164 25764 58216 25770
rect 58164 25706 58216 25712
rect 58176 25673 58204 25706
rect 58162 25664 58218 25673
rect 58162 25599 58218 25608
rect 58072 24812 58124 24818
rect 58072 24754 58124 24760
rect 57428 24744 57480 24750
rect 57428 24686 57480 24692
rect 58162 24712 58218 24721
rect 57336 24676 57388 24682
rect 57336 24618 57388 24624
rect 57440 24274 57468 24686
rect 58162 24647 58218 24656
rect 57980 24608 58032 24614
rect 57980 24550 58032 24556
rect 57992 24342 58020 24550
rect 58176 24342 58204 24647
rect 57980 24336 58032 24342
rect 57980 24278 58032 24284
rect 58164 24336 58216 24342
rect 58164 24278 58216 24284
rect 57428 24268 57480 24274
rect 57428 24210 57480 24216
rect 58162 24168 58218 24177
rect 58162 24103 58218 24112
rect 58176 23798 58204 24103
rect 58164 23792 58216 23798
rect 58164 23734 58216 23740
rect 57336 23656 57388 23662
rect 57336 23598 57388 23604
rect 57348 22137 57376 23598
rect 58072 23588 58124 23594
rect 58072 23530 58124 23536
rect 57980 23180 58032 23186
rect 57980 23122 58032 23128
rect 57520 22976 57572 22982
rect 57520 22918 57572 22924
rect 57532 22642 57560 22918
rect 57992 22778 58020 23122
rect 57980 22772 58032 22778
rect 57980 22714 58032 22720
rect 57520 22636 57572 22642
rect 57520 22578 57572 22584
rect 57334 22128 57390 22137
rect 57334 22063 57390 22072
rect 57980 22092 58032 22098
rect 57980 22034 58032 22040
rect 57992 21690 58020 22034
rect 58084 22030 58112 23530
rect 58162 23080 58218 23089
rect 58162 23015 58164 23024
rect 58216 23015 58218 23024
rect 58164 22986 58216 22992
rect 58072 22024 58124 22030
rect 58072 21966 58124 21972
rect 58164 21956 58216 21962
rect 58164 21898 58216 21904
rect 57980 21684 58032 21690
rect 57980 21626 58032 21632
rect 58176 21593 58204 21898
rect 58268 21622 58296 25774
rect 58256 21616 58308 21622
rect 58162 21584 58218 21593
rect 58256 21558 58308 21564
rect 58162 21519 58218 21528
rect 57520 21480 57572 21486
rect 57520 21422 57572 21428
rect 57704 21480 57756 21486
rect 57704 21422 57756 21428
rect 57428 21344 57480 21350
rect 57428 21286 57480 21292
rect 57440 19310 57468 21286
rect 57532 21078 57560 21422
rect 57716 21146 57744 21422
rect 57704 21140 57756 21146
rect 57704 21082 57756 21088
rect 57520 21072 57572 21078
rect 57520 21014 57572 21020
rect 58162 21040 58218 21049
rect 58162 20975 58164 20984
rect 58216 20975 58218 20984
rect 58164 20946 58216 20952
rect 57704 20392 57756 20398
rect 57704 20334 57756 20340
rect 57716 19514 57744 20334
rect 57980 20256 58032 20262
rect 57980 20198 58032 20204
rect 57992 19990 58020 20198
rect 57980 19984 58032 19990
rect 57980 19926 58032 19932
rect 58162 19952 58218 19961
rect 58162 19887 58164 19896
rect 58216 19887 58218 19896
rect 58164 19858 58216 19864
rect 57980 19712 58032 19718
rect 57980 19654 58032 19660
rect 57704 19508 57756 19514
rect 57704 19450 57756 19456
rect 57992 19310 58020 19654
rect 58162 19408 58218 19417
rect 58162 19343 58218 19352
rect 58176 19310 58204 19343
rect 57428 19304 57480 19310
rect 57428 19246 57480 19252
rect 57980 19304 58032 19310
rect 57980 19246 58032 19252
rect 58164 19304 58216 19310
rect 58164 19246 58216 19252
rect 57440 18222 57468 19246
rect 57980 18828 58032 18834
rect 57980 18770 58032 18776
rect 57520 18624 57572 18630
rect 57520 18566 57572 18572
rect 57532 18290 57560 18566
rect 57992 18426 58020 18770
rect 58164 18692 58216 18698
rect 58164 18634 58216 18640
rect 58176 18465 58204 18634
rect 58162 18456 58218 18465
rect 57980 18420 58032 18426
rect 58162 18391 58218 18400
rect 57980 18362 58032 18368
rect 57520 18284 57572 18290
rect 57520 18226 57572 18232
rect 57428 18216 57480 18222
rect 57428 18158 57480 18164
rect 58162 17912 58218 17921
rect 58162 17847 58218 17856
rect 58176 17814 58204 17847
rect 58164 17808 58216 17814
rect 58164 17750 58216 17756
rect 57520 17128 57572 17134
rect 57520 17070 57572 17076
rect 57256 16546 57468 16574
rect 56600 16244 56652 16250
rect 56600 16186 56652 16192
rect 56324 16040 56376 16046
rect 56324 15982 56376 15988
rect 56324 15904 56376 15910
rect 56324 15846 56376 15852
rect 56336 15570 56364 15846
rect 56324 15564 56376 15570
rect 56324 15506 56376 15512
rect 56140 14952 56192 14958
rect 56140 14894 56192 14900
rect 56152 13870 56180 14894
rect 56612 14482 56640 16186
rect 57060 15972 57112 15978
rect 57060 15914 57112 15920
rect 56692 15564 56744 15570
rect 56692 15506 56744 15512
rect 56876 15564 56928 15570
rect 56876 15506 56928 15512
rect 56600 14476 56652 14482
rect 56600 14418 56652 14424
rect 56704 13870 56732 15506
rect 56888 15162 56916 15506
rect 56968 15360 57020 15366
rect 56968 15302 57020 15308
rect 56876 15156 56928 15162
rect 56876 15098 56928 15104
rect 56980 14793 57008 15302
rect 56966 14784 57022 14793
rect 56966 14719 57022 14728
rect 56784 14000 56836 14006
rect 56784 13942 56836 13948
rect 56140 13864 56192 13870
rect 56140 13806 56192 13812
rect 56692 13864 56744 13870
rect 56692 13806 56744 13812
rect 56152 12986 56180 13806
rect 56796 13394 56824 13942
rect 56784 13388 56836 13394
rect 56784 13330 56836 13336
rect 56140 12980 56192 12986
rect 56140 12922 56192 12928
rect 55404 12776 55456 12782
rect 55402 12744 55404 12753
rect 56048 12776 56100 12782
rect 55456 12744 55458 12753
rect 56048 12718 56100 12724
rect 55402 12679 55458 12688
rect 55588 12232 55640 12238
rect 55588 12174 55640 12180
rect 55600 11898 55628 12174
rect 55588 11892 55640 11898
rect 55588 11834 55640 11840
rect 55588 11212 55640 11218
rect 55588 11154 55640 11160
rect 55600 11121 55628 11154
rect 55586 11112 55642 11121
rect 55586 11047 55642 11056
rect 55588 10124 55640 10130
rect 55588 10066 55640 10072
rect 55600 9625 55628 10066
rect 55586 9616 55642 9625
rect 55586 9551 55642 9560
rect 55680 9512 55732 9518
rect 55680 9454 55732 9460
rect 55692 7993 55720 9454
rect 56060 8430 56088 12718
rect 56152 11694 56180 12922
rect 56876 12300 56928 12306
rect 56876 12242 56928 12248
rect 56508 12096 56560 12102
rect 56508 12038 56560 12044
rect 56140 11688 56192 11694
rect 56520 11665 56548 12038
rect 56888 11898 56916 12242
rect 56876 11892 56928 11898
rect 56876 11834 56928 11840
rect 56140 11630 56192 11636
rect 56506 11656 56562 11665
rect 56506 11591 56562 11600
rect 56784 9512 56836 9518
rect 56784 9454 56836 9460
rect 56968 9512 57020 9518
rect 56968 9454 57020 9460
rect 56140 9104 56192 9110
rect 56140 9046 56192 9052
rect 56152 8634 56180 9046
rect 56140 8628 56192 8634
rect 56140 8570 56192 8576
rect 56048 8424 56100 8430
rect 56048 8366 56100 8372
rect 55772 8356 55824 8362
rect 55772 8298 55824 8304
rect 55678 7984 55734 7993
rect 55128 7948 55180 7954
rect 55678 7919 55734 7928
rect 55128 7890 55180 7896
rect 54300 6656 54352 6662
rect 54300 6598 54352 6604
rect 54484 6656 54536 6662
rect 54484 6598 54536 6604
rect 54024 6248 54076 6254
rect 54024 6190 54076 6196
rect 53932 3936 53984 3942
rect 53932 3878 53984 3884
rect 53840 2576 53892 2582
rect 53840 2518 53892 2524
rect 53944 800 53972 3878
rect 54036 3058 54064 6190
rect 54312 4622 54340 6598
rect 54300 4616 54352 4622
rect 54300 4558 54352 4564
rect 54392 4480 54444 4486
rect 54392 4422 54444 4428
rect 54404 4214 54432 4422
rect 54392 4208 54444 4214
rect 54392 4150 54444 4156
rect 54116 4004 54168 4010
rect 54116 3946 54168 3952
rect 54128 3738 54156 3946
rect 54116 3732 54168 3738
rect 54116 3674 54168 3680
rect 54300 3596 54352 3602
rect 54300 3538 54352 3544
rect 54312 3194 54340 3538
rect 54300 3188 54352 3194
rect 54300 3130 54352 3136
rect 54496 3058 54524 6598
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 54760 6112 54812 6118
rect 54760 6054 54812 6060
rect 54576 4684 54628 4690
rect 54576 4626 54628 4632
rect 54588 4078 54616 4626
rect 54576 4072 54628 4078
rect 54576 4014 54628 4020
rect 54668 4004 54720 4010
rect 54668 3946 54720 3952
rect 54680 3194 54708 3946
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54772 3126 54800 6054
rect 54956 5370 54984 6190
rect 54944 5364 54996 5370
rect 54944 5306 54996 5312
rect 55036 4548 55088 4554
rect 55036 4490 55088 4496
rect 55048 4146 55076 4490
rect 55036 4140 55088 4146
rect 55036 4082 55088 4088
rect 54852 3936 54904 3942
rect 54852 3878 54904 3884
rect 54760 3120 54812 3126
rect 54760 3062 54812 3068
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 54484 3052 54536 3058
rect 54484 2994 54536 3000
rect 54864 800 54892 3878
rect 55140 3369 55168 7890
rect 55680 7744 55732 7750
rect 55680 7686 55732 7692
rect 55220 7404 55272 7410
rect 55220 7346 55272 7352
rect 55232 4865 55260 7346
rect 55404 7336 55456 7342
rect 55404 7278 55456 7284
rect 55588 7336 55640 7342
rect 55588 7278 55640 7284
rect 55218 4856 55274 4865
rect 55218 4791 55274 4800
rect 55312 4480 55364 4486
rect 55312 4422 55364 4428
rect 55324 3602 55352 4422
rect 55312 3596 55364 3602
rect 55312 3538 55364 3544
rect 55126 3360 55182 3369
rect 55126 3295 55182 3304
rect 55416 3058 55444 7278
rect 55496 6724 55548 6730
rect 55496 6666 55548 6672
rect 55508 6497 55536 6666
rect 55494 6488 55550 6497
rect 55494 6423 55550 6432
rect 55494 6352 55550 6361
rect 55494 6287 55496 6296
rect 55548 6287 55550 6296
rect 55496 6258 55548 6264
rect 55600 6254 55628 7278
rect 55692 7206 55720 7686
rect 55680 7200 55732 7206
rect 55680 7142 55732 7148
rect 55784 6866 55812 8298
rect 56060 7426 56088 8366
rect 56152 8362 56180 8570
rect 56416 8492 56468 8498
rect 56416 8434 56468 8440
rect 56140 8356 56192 8362
rect 56140 8298 56192 8304
rect 56232 7744 56284 7750
rect 56232 7686 56284 7692
rect 55968 7398 56088 7426
rect 55772 6860 55824 6866
rect 55772 6802 55824 6808
rect 55588 6248 55640 6254
rect 55588 6190 55640 6196
rect 55600 4570 55628 6190
rect 55784 6066 55812 6802
rect 55864 6656 55916 6662
rect 55864 6598 55916 6604
rect 55876 6118 55904 6598
rect 55692 6038 55812 6066
rect 55864 6112 55916 6118
rect 55864 6054 55916 6060
rect 55692 5846 55720 6038
rect 55680 5840 55732 5846
rect 55680 5782 55732 5788
rect 55968 5234 55996 7398
rect 56048 7268 56100 7274
rect 56048 7210 56100 7216
rect 55956 5228 56008 5234
rect 55956 5170 56008 5176
rect 55864 5092 55916 5098
rect 55864 5034 55916 5040
rect 55772 5024 55824 5030
rect 55772 4966 55824 4972
rect 55600 4542 55720 4570
rect 55588 4480 55640 4486
rect 55588 4422 55640 4428
rect 55600 3670 55628 4422
rect 55692 4078 55720 4542
rect 55680 4072 55732 4078
rect 55680 4014 55732 4020
rect 55692 3670 55720 4014
rect 55588 3664 55640 3670
rect 55588 3606 55640 3612
rect 55680 3664 55732 3670
rect 55680 3606 55732 3612
rect 55404 3052 55456 3058
rect 55404 2994 55456 3000
rect 55220 2916 55272 2922
rect 55220 2858 55272 2864
rect 55232 2582 55260 2858
rect 55220 2576 55272 2582
rect 55220 2518 55272 2524
rect 55588 2372 55640 2378
rect 55588 2314 55640 2320
rect 52368 750 52420 756
rect 53010 0 53066 800
rect 53930 0 53986 800
rect 54850 0 54906 800
rect 55600 649 55628 2314
rect 55784 800 55812 4966
rect 55876 3194 55904 5034
rect 55956 3460 56008 3466
rect 55956 3402 56008 3408
rect 55864 3188 55916 3194
rect 55864 3130 55916 3136
rect 55968 2281 55996 3402
rect 56060 2514 56088 7210
rect 56140 6656 56192 6662
rect 56140 6598 56192 6604
rect 56152 6254 56180 6598
rect 56140 6248 56192 6254
rect 56140 6190 56192 6196
rect 56244 4078 56272 7686
rect 56428 7342 56456 8434
rect 56796 7954 56824 9454
rect 56980 9042 57008 9454
rect 56968 9036 57020 9042
rect 56968 8978 57020 8984
rect 56784 7948 56836 7954
rect 56784 7890 56836 7896
rect 56416 7336 56468 7342
rect 56416 7278 56468 7284
rect 56508 7200 56560 7206
rect 56508 7142 56560 7148
rect 56414 6896 56470 6905
rect 56414 6831 56470 6840
rect 56428 6390 56456 6831
rect 56416 6384 56468 6390
rect 56416 6326 56468 6332
rect 56520 6322 56548 7142
rect 57072 7002 57100 15914
rect 57152 13864 57204 13870
rect 57152 13806 57204 13812
rect 57164 11218 57192 13806
rect 57244 13184 57296 13190
rect 57244 13126 57296 13132
rect 57334 13152 57390 13161
rect 57256 12782 57284 13126
rect 57334 13087 57390 13096
rect 57348 12986 57376 13087
rect 57336 12980 57388 12986
rect 57336 12922 57388 12928
rect 57244 12776 57296 12782
rect 57244 12718 57296 12724
rect 57152 11212 57204 11218
rect 57152 11154 57204 11160
rect 57164 10606 57192 11154
rect 57152 10600 57204 10606
rect 57152 10542 57204 10548
rect 57244 10600 57296 10606
rect 57244 10542 57296 10548
rect 57164 10130 57192 10542
rect 57256 10266 57284 10542
rect 57244 10260 57296 10266
rect 57244 10202 57296 10208
rect 57152 10124 57204 10130
rect 57152 10066 57204 10072
rect 57152 9512 57204 9518
rect 57152 9454 57204 9460
rect 57164 9178 57192 9454
rect 57152 9172 57204 9178
rect 57152 9114 57204 9120
rect 57440 8650 57468 16546
rect 57532 16182 57560 17070
rect 57980 16992 58032 16998
rect 57980 16934 58032 16940
rect 57992 16726 58020 16934
rect 58162 16824 58218 16833
rect 58162 16759 58218 16768
rect 58176 16726 58204 16759
rect 57980 16720 58032 16726
rect 57980 16662 58032 16668
rect 58164 16720 58216 16726
rect 58164 16662 58216 16668
rect 57980 16584 58032 16590
rect 57980 16526 58032 16532
rect 57520 16176 57572 16182
rect 57520 16118 57572 16124
rect 57992 14958 58020 16526
rect 58254 16280 58310 16289
rect 58254 16215 58310 16224
rect 58164 15972 58216 15978
rect 58164 15914 58216 15920
rect 58072 15904 58124 15910
rect 58072 15846 58124 15852
rect 58084 15337 58112 15846
rect 58176 15706 58204 15914
rect 58164 15700 58216 15706
rect 58164 15642 58216 15648
rect 58070 15328 58126 15337
rect 58070 15263 58126 15272
rect 58268 15094 58296 16215
rect 58256 15088 58308 15094
rect 58256 15030 58308 15036
rect 57980 14952 58032 14958
rect 57980 14894 58032 14900
rect 57520 13864 57572 13870
rect 57520 13806 57572 13812
rect 57532 13462 57560 13806
rect 58164 13728 58216 13734
rect 58070 13696 58126 13705
rect 58164 13670 58216 13676
rect 58070 13631 58126 13640
rect 58084 13530 58112 13631
rect 58072 13524 58124 13530
rect 58072 13466 58124 13472
rect 58176 13462 58204 13670
rect 57520 13456 57572 13462
rect 57520 13398 57572 13404
rect 58164 13456 58216 13462
rect 58164 13398 58216 13404
rect 57980 12708 58032 12714
rect 57980 12650 58032 12656
rect 57888 12640 57940 12646
rect 57888 12582 57940 12588
rect 57704 12232 57756 12238
rect 57900 12209 57928 12582
rect 57992 12442 58020 12650
rect 57980 12436 58032 12442
rect 57980 12378 58032 12384
rect 57704 12174 57756 12180
rect 57886 12200 57942 12209
rect 57716 11354 57744 12174
rect 57886 12135 57942 12144
rect 57704 11348 57756 11354
rect 57704 11290 57756 11296
rect 57980 11212 58032 11218
rect 57980 11154 58032 11160
rect 57888 11076 57940 11082
rect 57888 11018 57940 11024
rect 57900 10577 57928 11018
rect 57992 10810 58020 11154
rect 57980 10804 58032 10810
rect 57980 10746 58032 10752
rect 57886 10568 57942 10577
rect 57886 10503 57942 10512
rect 57704 10464 57756 10470
rect 57704 10406 57756 10412
rect 57612 10124 57664 10130
rect 57612 10066 57664 10072
rect 57624 9654 57652 10066
rect 57612 9648 57664 9654
rect 57612 9590 57664 9596
rect 57716 9042 57744 10406
rect 58162 10024 58218 10033
rect 58162 9959 58164 9968
rect 58216 9959 58218 9968
rect 58164 9930 58216 9936
rect 58162 9072 58218 9081
rect 57704 9036 57756 9042
rect 58162 9007 58218 9016
rect 57704 8978 57756 8984
rect 57980 8832 58032 8838
rect 57980 8774 58032 8780
rect 57256 8622 57468 8650
rect 57256 7274 57284 8622
rect 57336 8560 57388 8566
rect 57336 8502 57388 8508
rect 57426 8528 57482 8537
rect 57348 7954 57376 8502
rect 57426 8463 57428 8472
rect 57480 8463 57482 8472
rect 57428 8434 57480 8440
rect 57992 8430 58020 8774
rect 58176 8566 58204 9007
rect 58164 8560 58216 8566
rect 58164 8502 58216 8508
rect 57980 8424 58032 8430
rect 57980 8366 58032 8372
rect 57520 8356 57572 8362
rect 57520 8298 57572 8304
rect 57336 7948 57388 7954
rect 57336 7890 57388 7896
rect 57532 7818 57560 8298
rect 57336 7812 57388 7818
rect 57336 7754 57388 7760
rect 57520 7812 57572 7818
rect 57520 7754 57572 7760
rect 57244 7268 57296 7274
rect 57244 7210 57296 7216
rect 57060 6996 57112 7002
rect 57060 6938 57112 6944
rect 56600 6384 56652 6390
rect 56598 6352 56600 6361
rect 56652 6352 56654 6361
rect 56508 6316 56560 6322
rect 56598 6287 56654 6296
rect 56508 6258 56560 6264
rect 56968 6248 57020 6254
rect 56968 6190 57020 6196
rect 56692 6180 56744 6186
rect 56692 6122 56744 6128
rect 56704 5778 56732 6122
rect 56980 5914 57008 6190
rect 57152 6180 57204 6186
rect 57152 6122 57204 6128
rect 56968 5908 57020 5914
rect 56968 5850 57020 5856
rect 56508 5772 56560 5778
rect 56508 5714 56560 5720
rect 56692 5772 56744 5778
rect 56692 5714 56744 5720
rect 56416 4752 56468 4758
rect 56416 4694 56468 4700
rect 56232 4072 56284 4078
rect 56232 4014 56284 4020
rect 56428 3194 56456 4694
rect 56520 4146 56548 5714
rect 56784 5704 56836 5710
rect 56784 5646 56836 5652
rect 56692 4820 56744 4826
rect 56692 4762 56744 4768
rect 56600 4684 56652 4690
rect 56600 4626 56652 4632
rect 56508 4140 56560 4146
rect 56508 4082 56560 4088
rect 56612 3942 56640 4626
rect 56600 3936 56652 3942
rect 56600 3878 56652 3884
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 56600 3120 56652 3126
rect 56600 3062 56652 3068
rect 56612 2582 56640 3062
rect 56704 2650 56732 4762
rect 56796 4622 56824 5646
rect 56876 5568 56928 5574
rect 56876 5510 56928 5516
rect 57060 5568 57112 5574
rect 57060 5510 57112 5516
rect 56784 4616 56836 4622
rect 56784 4558 56836 4564
rect 56888 3618 56916 5510
rect 57072 5166 57100 5510
rect 57060 5160 57112 5166
rect 57060 5102 57112 5108
rect 57060 5024 57112 5030
rect 57060 4966 57112 4972
rect 56968 4480 57020 4486
rect 56968 4422 57020 4428
rect 56980 4321 57008 4422
rect 56966 4312 57022 4321
rect 56966 4247 57022 4256
rect 57072 3777 57100 4966
rect 57058 3768 57114 3777
rect 57058 3703 57114 3712
rect 56888 3602 57008 3618
rect 56784 3596 56836 3602
rect 56888 3596 57020 3602
rect 56888 3590 56968 3596
rect 56784 3538 56836 3544
rect 56968 3538 57020 3544
rect 56692 2644 56744 2650
rect 56692 2586 56744 2592
rect 56600 2576 56652 2582
rect 56600 2518 56652 2524
rect 56048 2508 56100 2514
rect 56048 2450 56100 2456
rect 55954 2272 56010 2281
rect 56796 2258 56824 3538
rect 57164 2990 57192 6122
rect 57244 6112 57296 6118
rect 57244 6054 57296 6060
rect 57256 3058 57284 6054
rect 57348 5234 57376 7754
rect 58162 7440 58218 7449
rect 58162 7375 58218 7384
rect 57704 7336 57756 7342
rect 57704 7278 57756 7284
rect 57716 6458 57744 7278
rect 57980 7200 58032 7206
rect 57980 7142 58032 7148
rect 58072 7200 58124 7206
rect 58072 7142 58124 7148
rect 57992 6866 58020 7142
rect 57980 6860 58032 6866
rect 57980 6802 58032 6808
rect 57704 6452 57756 6458
rect 57704 6394 57756 6400
rect 57428 6384 57480 6390
rect 57428 6326 57480 6332
rect 57336 5228 57388 5234
rect 57336 5170 57388 5176
rect 57440 3534 57468 6326
rect 57888 6112 57940 6118
rect 57888 6054 57940 6060
rect 57612 5840 57664 5846
rect 57612 5782 57664 5788
rect 57428 3528 57480 3534
rect 57428 3470 57480 3476
rect 57244 3052 57296 3058
rect 57244 2994 57296 3000
rect 57152 2984 57204 2990
rect 57152 2926 57204 2932
rect 55954 2207 56010 2216
rect 56704 2230 56824 2258
rect 56508 1760 56560 1766
rect 56506 1728 56508 1737
rect 56560 1728 56562 1737
rect 56506 1663 56562 1672
rect 56324 808 56376 814
rect 55586 640 55642 649
rect 55586 575 55642 584
rect 55770 0 55826 800
rect 56704 800 56732 2230
rect 57624 800 57652 5782
rect 57900 5409 57928 6054
rect 58084 5778 58112 7142
rect 58176 6866 58204 7375
rect 58164 6860 58216 6866
rect 58164 6802 58216 6808
rect 58162 5944 58218 5953
rect 58162 5879 58218 5888
rect 58176 5846 58204 5879
rect 58164 5840 58216 5846
rect 58164 5782 58216 5788
rect 58072 5772 58124 5778
rect 58072 5714 58124 5720
rect 57886 5400 57942 5409
rect 57886 5335 57942 5344
rect 57704 5160 57756 5166
rect 57704 5102 57756 5108
rect 57716 3738 57744 5102
rect 58164 5024 58216 5030
rect 58164 4966 58216 4972
rect 58176 4758 58204 4966
rect 58164 4752 58216 4758
rect 58164 4694 58216 4700
rect 57980 4480 58032 4486
rect 57980 4422 58032 4428
rect 57992 4078 58020 4422
rect 58532 4140 58584 4146
rect 58532 4082 58584 4088
rect 57980 4072 58032 4078
rect 57980 4014 58032 4020
rect 58164 4004 58216 4010
rect 58164 3946 58216 3952
rect 57704 3732 57756 3738
rect 57704 3674 57756 3680
rect 57980 3392 58032 3398
rect 57980 3334 58032 3340
rect 57992 2582 58020 3334
rect 58176 2825 58204 3946
rect 58162 2816 58218 2825
rect 58162 2751 58218 2760
rect 57980 2576 58032 2582
rect 57980 2518 58032 2524
rect 57888 2304 57940 2310
rect 57888 2246 57940 2252
rect 57900 1193 57928 2246
rect 57886 1184 57942 1193
rect 57886 1119 57942 1128
rect 58544 800 58572 4082
rect 59452 2916 59504 2922
rect 59452 2858 59504 2864
rect 59464 800 59492 2858
rect 56324 750 56376 756
rect 56336 241 56364 750
rect 56322 232 56378 241
rect 56322 167 56378 176
rect 56690 0 56746 800
rect 57610 0 57666 800
rect 58530 0 58586 800
rect 59450 0 59506 800
<< via2 >>
rect 2778 59472 2834 59528
rect 1214 58520 1270 58576
rect 1398 56616 1454 56672
rect 1398 55820 1454 55856
rect 1398 55800 1400 55820
rect 1400 55800 1452 55820
rect 1452 55800 1454 55820
rect 2134 57568 2190 57624
rect 56506 59608 56562 59664
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 1398 54848 1454 54904
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 1398 53896 1454 53952
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 1398 52980 1400 53000
rect 1400 52980 1452 53000
rect 1452 52980 1454 53000
rect 1398 52944 1454 52980
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 1398 51992 1454 52048
rect 1398 51176 1454 51232
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 1398 50224 1454 50280
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 1398 49292 1454 49328
rect 1398 49272 1400 49292
rect 1400 49272 1452 49292
rect 1452 49272 1454 49292
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 1398 48320 1454 48376
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 1398 47540 1400 47560
rect 1400 47540 1452 47560
rect 1452 47540 1454 47560
rect 1398 47504 1454 47540
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 1398 46552 1454 46608
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 1398 45600 1454 45656
rect 1398 44648 1454 44704
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 1398 43696 1454 43752
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 1398 42880 1454 42936
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 1398 41928 1454 41984
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 1398 41012 1400 41032
rect 1400 41012 1452 41032
rect 1452 41012 1454 41032
rect 1398 40976 1454 41012
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 1398 40024 1454 40080
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 1398 39072 1454 39128
rect 1398 38256 1454 38312
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 1398 37324 1454 37360
rect 1398 37304 1400 37324
rect 1400 37304 1452 37324
rect 1452 37304 1454 37324
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 1398 36352 1454 36408
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 1398 35400 1454 35456
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 1398 34584 1454 34640
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 1398 33632 1454 33688
rect 1398 32680 1454 32736
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 1398 31728 1454 31784
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 1398 30796 1454 30832
rect 1398 30776 1400 30796
rect 1400 30776 1452 30796
rect 1452 30776 1454 30796
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 1398 29960 1454 30016
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 1950 29008 2006 29064
rect 2042 28056 2098 28112
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 5078 28464 5134 28520
rect 1950 27104 2006 27160
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 1398 26152 1454 26208
rect 1950 24384 2006 24440
rect 1582 23468 1584 23488
rect 1584 23468 1636 23488
rect 1636 23468 1638 23488
rect 1582 23432 1638 23468
rect 1950 22480 2006 22536
rect 1950 21684 2006 21720
rect 1950 21664 1952 21684
rect 1952 21664 2004 21684
rect 2004 21664 2006 21684
rect 1950 20748 1952 20768
rect 1952 20748 2004 20768
rect 2004 20748 2006 20768
rect 1950 20712 2006 20748
rect 1858 19780 1914 19816
rect 1858 19760 1860 19780
rect 1860 19760 1912 19780
rect 1912 19760 1914 19780
rect 2042 18844 2044 18864
rect 2044 18844 2096 18864
rect 2096 18844 2098 18864
rect 2042 18808 2098 18844
rect 1950 17876 2006 17912
rect 1950 17856 1952 17876
rect 1952 17856 2004 17876
rect 2004 17856 2006 17876
rect 3146 25336 3202 25392
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 2042 17060 2098 17096
rect 2042 17040 2044 17060
rect 2044 17040 2096 17060
rect 2096 17040 2098 17060
rect 2042 16108 2098 16144
rect 2042 16088 2044 16108
rect 2044 16088 2096 16108
rect 2096 16088 2098 16108
rect 1950 15156 2006 15192
rect 1950 15136 1952 15156
rect 1952 15136 2004 15156
rect 2004 15136 2006 15156
rect 1950 14220 1952 14240
rect 1952 14220 2004 14240
rect 2004 14220 2006 14240
rect 1950 14184 2006 14220
rect 2042 13252 2098 13288
rect 2042 13232 2044 13252
rect 2044 13232 2096 13252
rect 2096 13232 2098 13252
rect 1950 12436 2006 12472
rect 1950 12416 1952 12436
rect 1952 12416 2004 12436
rect 2004 12416 2006 12436
rect 1950 11500 1952 11520
rect 1952 11500 2004 11520
rect 2004 11500 2006 11520
rect 1950 11464 2006 11500
rect 2042 10532 2098 10568
rect 2042 10512 2044 10532
rect 2044 10512 2096 10532
rect 2096 10512 2098 10532
rect 2042 9596 2044 9616
rect 2044 9596 2096 9616
rect 2096 9596 2098 9616
rect 2042 9560 2098 9596
rect 1950 8780 1952 8800
rect 1952 8780 2004 8800
rect 2004 8780 2006 8800
rect 1950 8744 2006 8780
rect 2042 7812 2098 7848
rect 2042 7792 2044 7812
rect 2044 7792 2096 7812
rect 2096 7792 2098 7812
rect 2042 6840 2098 6896
rect 1950 5908 2006 5944
rect 1950 5888 1952 5908
rect 1952 5888 2004 5908
rect 2004 5888 2006 5908
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 1950 4972 1952 4992
rect 1952 4972 2004 4992
rect 2004 4972 2006 4992
rect 1950 4936 2006 4972
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 2042 4140 2098 4176
rect 2042 4120 2044 4140
rect 2044 4120 2096 4140
rect 2096 4120 2098 4140
rect 1950 2216 2006 2272
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 3054 3188 3110 3224
rect 3054 3168 3056 3188
rect 3056 3168 3108 3188
rect 3108 3168 3110 3188
rect 2778 1264 2834 1320
rect 8206 28464 8262 28520
rect 7470 24268 7526 24304
rect 7470 24248 7472 24268
rect 7472 24248 7524 24268
rect 7524 24248 7526 24268
rect 9678 28756 9734 28792
rect 9678 28736 9680 28756
rect 9680 28736 9732 28756
rect 9732 28736 9734 28756
rect 10138 26968 10194 27024
rect 10690 26968 10746 27024
rect 10782 26444 10838 26480
rect 10782 26424 10784 26444
rect 10784 26424 10836 26444
rect 10836 26424 10838 26444
rect 9586 24112 9642 24168
rect 10138 24384 10194 24440
rect 10782 24384 10838 24440
rect 10782 23976 10838 24032
rect 11334 24384 11390 24440
rect 11978 26444 12034 26480
rect 11978 26424 11980 26444
rect 11980 26424 12032 26444
rect 12032 26424 12034 26444
rect 12254 27276 12256 27296
rect 12256 27276 12308 27296
rect 12308 27276 12310 27296
rect 12254 27240 12310 27276
rect 12714 26868 12716 26888
rect 12716 26868 12768 26888
rect 12768 26868 12770 26888
rect 12714 26832 12770 26868
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 25594 57568 25650 57624
rect 28354 57024 28410 57080
rect 29274 57568 29330 57624
rect 29274 57024 29330 57080
rect 29550 56888 29606 56944
rect 29090 56772 29146 56808
rect 31114 57024 31170 57080
rect 29090 56752 29092 56772
rect 29092 56752 29144 56772
rect 29144 56752 29146 56772
rect 29642 56752 29698 56808
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 32954 56344 33010 56400
rect 31942 55800 31998 55856
rect 33046 56228 33102 56264
rect 33046 56208 33048 56228
rect 33048 56208 33100 56228
rect 33100 56208 33102 56228
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 11978 23724 12034 23760
rect 11978 23704 11980 23724
rect 11980 23704 12032 23724
rect 12032 23704 12034 23724
rect 12438 24112 12494 24168
rect 13266 21800 13322 21856
rect 13818 27240 13874 27296
rect 12254 18672 12310 18728
rect 14186 26696 14242 26752
rect 14462 27784 14518 27840
rect 14002 26016 14058 26072
rect 15842 28736 15898 28792
rect 15106 25780 15108 25800
rect 15108 25780 15160 25800
rect 15160 25780 15162 25800
rect 15106 25744 15162 25780
rect 12438 18148 12494 18184
rect 12438 18128 12440 18148
rect 12440 18128 12492 18148
rect 12492 18128 12494 18148
rect 15566 25608 15622 25664
rect 15566 22072 15622 22128
rect 15106 19216 15162 19272
rect 16118 26968 16174 27024
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 16578 26968 16634 27024
rect 16486 26424 16542 26480
rect 16670 26016 16726 26072
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 17866 28600 17922 28656
rect 17038 27104 17094 27160
rect 16946 26832 17002 26888
rect 18050 28464 18106 28520
rect 17958 27956 17960 27976
rect 17960 27956 18012 27976
rect 18012 27956 18014 27976
rect 17958 27920 18014 27956
rect 18142 27784 18198 27840
rect 17590 26868 17592 26888
rect 17592 26868 17644 26888
rect 17644 26868 17646 26888
rect 17590 26832 17646 26868
rect 17958 26696 18014 26752
rect 17866 26424 17922 26480
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19614 30132 19616 30152
rect 19616 30132 19668 30152
rect 19668 30132 19670 30152
rect 19614 30096 19670 30132
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19430 29044 19432 29064
rect 19432 29044 19484 29064
rect 19484 29044 19486 29064
rect 19430 29008 19486 29044
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 18694 27920 18750 27976
rect 19154 27920 19210 27976
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 18786 27104 18842 27160
rect 18418 26852 18474 26888
rect 18418 26832 18420 26852
rect 18420 26832 18472 26852
rect 18472 26832 18474 26852
rect 18510 26016 18566 26072
rect 18418 25880 18474 25936
rect 18142 25608 18198 25664
rect 16118 19252 16120 19272
rect 16120 19252 16172 19272
rect 16172 19252 16174 19272
rect 16118 19216 16174 19252
rect 16486 22072 16542 22128
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 17130 18672 17186 18728
rect 17958 23976 18014 24032
rect 17682 21020 17684 21040
rect 17684 21020 17736 21040
rect 17736 21020 17738 21040
rect 17682 20984 17738 21020
rect 19062 25744 19118 25800
rect 18970 25608 19026 25664
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 18694 23704 18750 23760
rect 18234 22092 18290 22128
rect 18234 22072 18236 22092
rect 18236 22072 18288 22092
rect 18288 22072 18290 22092
rect 18142 21836 18144 21856
rect 18144 21836 18196 21856
rect 18196 21836 18198 21856
rect 18142 21800 18198 21836
rect 19338 22652 19340 22672
rect 19340 22652 19392 22672
rect 19392 22652 19394 22672
rect 19338 22616 19394 22652
rect 19338 22072 19394 22128
rect 19246 21004 19302 21040
rect 19246 20984 19248 21004
rect 19248 20984 19300 21004
rect 19300 20984 19302 21004
rect 18050 18128 18106 18184
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 20074 22888 20130 22944
rect 19798 22480 19854 22536
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19798 20868 19854 20904
rect 19798 20848 19800 20868
rect 19800 20848 19852 20868
rect 19852 20848 19854 20868
rect 19614 20440 19670 20496
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 20074 21292 20076 21312
rect 20076 21292 20128 21312
rect 20128 21292 20130 21312
rect 20074 21256 20130 21292
rect 20258 20984 20314 21040
rect 19522 19236 19578 19272
rect 19522 19216 19524 19236
rect 19524 19216 19576 19236
rect 19576 19216 19578 19236
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 21086 26988 21142 27024
rect 21086 26968 21088 26988
rect 21088 26968 21140 26988
rect 21140 26968 21142 26988
rect 20718 23180 20774 23216
rect 20718 23160 20720 23180
rect 20720 23160 20772 23180
rect 20772 23160 20774 23180
rect 20810 22344 20866 22400
rect 21822 26968 21878 27024
rect 21362 26868 21364 26888
rect 21364 26868 21416 26888
rect 21416 26868 21418 26888
rect 21362 26832 21418 26868
rect 21270 26016 21326 26072
rect 21362 25916 21364 25936
rect 21364 25916 21416 25936
rect 21416 25916 21418 25936
rect 21362 25880 21418 25916
rect 20534 20576 20590 20632
rect 20902 20440 20958 20496
rect 20534 20304 20590 20360
rect 21270 20576 21326 20632
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 22006 26832 22062 26888
rect 22466 30096 22522 30152
rect 22190 26968 22246 27024
rect 21914 24132 21970 24168
rect 21914 24112 21916 24132
rect 21916 24112 21968 24132
rect 21968 24112 21970 24132
rect 23110 32292 23166 32328
rect 23110 32272 23112 32292
rect 23112 32272 23164 32292
rect 23164 32272 23166 32292
rect 24030 32292 24086 32328
rect 24030 32272 24032 32292
rect 24032 32272 24084 32292
rect 24084 32272 24086 32292
rect 23478 29028 23534 29064
rect 23478 29008 23480 29028
rect 23480 29008 23532 29028
rect 23532 29008 23534 29028
rect 22466 25744 22522 25800
rect 23294 24656 23350 24712
rect 23662 26288 23718 26344
rect 22190 23432 22246 23488
rect 21822 23160 21878 23216
rect 21638 22344 21694 22400
rect 21822 22092 21878 22128
rect 21822 22072 21824 22092
rect 21824 22072 21876 22092
rect 21876 22072 21878 22092
rect 22926 22072 22982 22128
rect 23386 23568 23442 23624
rect 22926 19896 22982 19952
rect 23846 23180 23902 23216
rect 23846 23160 23848 23180
rect 23848 23160 23900 23180
rect 23900 23160 23902 23180
rect 24214 23432 24270 23488
rect 24306 23024 24362 23080
rect 24030 22480 24086 22536
rect 23570 21800 23626 21856
rect 23570 20340 23572 20360
rect 23572 20340 23624 20360
rect 23624 20340 23626 20360
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 23570 20304 23626 20340
rect 25502 24692 25504 24712
rect 25504 24692 25556 24712
rect 25556 24692 25558 24712
rect 25502 24656 25558 24692
rect 25042 23568 25098 23624
rect 24398 21292 24400 21312
rect 24400 21292 24452 21312
rect 24452 21292 24454 21312
rect 24398 21256 24454 21292
rect 24674 21256 24730 21312
rect 25410 22480 25466 22536
rect 26514 26288 26570 26344
rect 26514 24656 26570 24712
rect 25318 21004 25374 21040
rect 25318 20984 25320 21004
rect 25320 20984 25372 21004
rect 25372 20984 25374 21004
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 25778 19896 25834 19952
rect 26698 24112 26754 24168
rect 29826 30132 29828 30152
rect 29828 30132 29880 30152
rect 29880 30132 29882 30152
rect 29826 30096 29882 30132
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 31942 52980 31944 53000
rect 31944 52980 31996 53000
rect 31996 52980 31998 53000
rect 31942 52944 31998 52980
rect 35622 57024 35678 57080
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 35898 56908 35954 56944
rect 35898 56888 35900 56908
rect 35900 56888 35952 56908
rect 35952 56888 35954 56908
rect 34978 56344 35034 56400
rect 36082 56208 36138 56264
rect 36450 55800 36506 55856
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34702 52980 34704 53000
rect 34704 52980 34756 53000
rect 34756 52980 34758 53000
rect 34702 52944 34758 52980
rect 50300 57146 50356 57148
rect 50380 57146 50436 57148
rect 50460 57146 50516 57148
rect 50540 57146 50596 57148
rect 50300 57094 50326 57146
rect 50326 57094 50356 57146
rect 50380 57094 50390 57146
rect 50390 57094 50436 57146
rect 50460 57094 50506 57146
rect 50506 57094 50516 57146
rect 50540 57094 50570 57146
rect 50570 57094 50596 57146
rect 50300 57092 50356 57094
rect 50380 57092 50436 57094
rect 50460 57092 50516 57094
rect 50540 57092 50596 57094
rect 50300 56058 50356 56060
rect 50380 56058 50436 56060
rect 50460 56058 50516 56060
rect 50540 56058 50596 56060
rect 50300 56006 50326 56058
rect 50326 56006 50356 56058
rect 50380 56006 50390 56058
rect 50390 56006 50436 56058
rect 50460 56006 50506 56058
rect 50506 56006 50516 56058
rect 50540 56006 50570 56058
rect 50570 56006 50596 56058
rect 50300 56004 50356 56006
rect 50380 56004 50436 56006
rect 50460 56004 50516 56006
rect 50540 56004 50596 56006
rect 55126 58248 55182 58304
rect 50300 54970 50356 54972
rect 50380 54970 50436 54972
rect 50460 54970 50516 54972
rect 50540 54970 50596 54972
rect 50300 54918 50326 54970
rect 50326 54918 50356 54970
rect 50380 54918 50390 54970
rect 50390 54918 50436 54970
rect 50460 54918 50506 54970
rect 50506 54918 50516 54970
rect 50540 54918 50570 54970
rect 50570 54918 50596 54970
rect 50300 54916 50356 54918
rect 50380 54916 50436 54918
rect 50460 54916 50516 54918
rect 50540 54916 50596 54918
rect 50300 53882 50356 53884
rect 50380 53882 50436 53884
rect 50460 53882 50516 53884
rect 50540 53882 50596 53884
rect 50300 53830 50326 53882
rect 50326 53830 50356 53882
rect 50380 53830 50390 53882
rect 50390 53830 50436 53882
rect 50460 53830 50506 53882
rect 50506 53830 50516 53882
rect 50540 53830 50570 53882
rect 50570 53830 50596 53882
rect 50300 53828 50356 53830
rect 50380 53828 50436 53830
rect 50460 53828 50516 53830
rect 50540 53828 50596 53830
rect 50300 52794 50356 52796
rect 50380 52794 50436 52796
rect 50460 52794 50516 52796
rect 50540 52794 50596 52796
rect 50300 52742 50326 52794
rect 50326 52742 50356 52794
rect 50380 52742 50390 52794
rect 50390 52742 50436 52794
rect 50460 52742 50506 52794
rect 50506 52742 50516 52794
rect 50540 52742 50570 52794
rect 50570 52742 50596 52794
rect 50300 52740 50356 52742
rect 50380 52740 50436 52742
rect 50460 52740 50516 52742
rect 50540 52740 50596 52742
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 30470 30132 30472 30152
rect 30472 30132 30524 30152
rect 30524 30132 30526 30152
rect 30470 30096 30526 30132
rect 30286 28056 30342 28112
rect 30470 27920 30526 27976
rect 27802 24656 27858 24712
rect 26422 22888 26478 22944
rect 27066 22480 27122 22536
rect 26698 20848 26754 20904
rect 26974 20984 27030 21040
rect 27894 22480 27950 22536
rect 27986 22072 28042 22128
rect 27342 21800 27398 21856
rect 28630 22616 28686 22672
rect 29090 26832 29146 26888
rect 28814 23180 28870 23216
rect 28814 23160 28816 23180
rect 28816 23160 28868 23180
rect 28868 23160 28870 23180
rect 28722 22072 28778 22128
rect 28814 21256 28870 21312
rect 29458 23024 29514 23080
rect 28722 19216 28778 19272
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 50300 51706 50356 51708
rect 50380 51706 50436 51708
rect 50460 51706 50516 51708
rect 50540 51706 50596 51708
rect 50300 51654 50326 51706
rect 50326 51654 50356 51706
rect 50380 51654 50390 51706
rect 50390 51654 50436 51706
rect 50460 51654 50506 51706
rect 50506 51654 50516 51706
rect 50540 51654 50570 51706
rect 50570 51654 50596 51706
rect 50300 51652 50356 51654
rect 50380 51652 50436 51654
rect 50460 51652 50516 51654
rect 50540 51652 50596 51654
rect 50300 50618 50356 50620
rect 50380 50618 50436 50620
rect 50460 50618 50516 50620
rect 50540 50618 50596 50620
rect 50300 50566 50326 50618
rect 50326 50566 50356 50618
rect 50380 50566 50390 50618
rect 50390 50566 50436 50618
rect 50460 50566 50506 50618
rect 50506 50566 50516 50618
rect 50540 50566 50570 50618
rect 50570 50566 50596 50618
rect 50300 50564 50356 50566
rect 50380 50564 50436 50566
rect 50460 50564 50516 50566
rect 50540 50564 50596 50566
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 50300 49530 50356 49532
rect 50380 49530 50436 49532
rect 50460 49530 50516 49532
rect 50540 49530 50596 49532
rect 50300 49478 50326 49530
rect 50326 49478 50356 49530
rect 50380 49478 50390 49530
rect 50390 49478 50436 49530
rect 50460 49478 50506 49530
rect 50506 49478 50516 49530
rect 50540 49478 50570 49530
rect 50570 49478 50596 49530
rect 50300 49476 50356 49478
rect 50380 49476 50436 49478
rect 50460 49476 50516 49478
rect 50540 49476 50596 49478
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 50300 48442 50356 48444
rect 50380 48442 50436 48444
rect 50460 48442 50516 48444
rect 50540 48442 50596 48444
rect 50300 48390 50326 48442
rect 50326 48390 50356 48442
rect 50380 48390 50390 48442
rect 50390 48390 50436 48442
rect 50460 48390 50506 48442
rect 50506 48390 50516 48442
rect 50540 48390 50570 48442
rect 50570 48390 50596 48442
rect 50300 48388 50356 48390
rect 50380 48388 50436 48390
rect 50460 48388 50516 48390
rect 50540 48388 50596 48390
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 50300 47354 50356 47356
rect 50380 47354 50436 47356
rect 50460 47354 50516 47356
rect 50540 47354 50596 47356
rect 50300 47302 50326 47354
rect 50326 47302 50356 47354
rect 50380 47302 50390 47354
rect 50390 47302 50436 47354
rect 50460 47302 50506 47354
rect 50506 47302 50516 47354
rect 50540 47302 50570 47354
rect 50570 47302 50596 47354
rect 50300 47300 50356 47302
rect 50380 47300 50436 47302
rect 50460 47300 50516 47302
rect 50540 47300 50596 47302
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 50300 46266 50356 46268
rect 50380 46266 50436 46268
rect 50460 46266 50516 46268
rect 50540 46266 50596 46268
rect 50300 46214 50326 46266
rect 50326 46214 50356 46266
rect 50380 46214 50390 46266
rect 50390 46214 50436 46266
rect 50460 46214 50506 46266
rect 50506 46214 50516 46266
rect 50540 46214 50570 46266
rect 50570 46214 50596 46266
rect 50300 46212 50356 46214
rect 50380 46212 50436 46214
rect 50460 46212 50516 46214
rect 50540 46212 50596 46214
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 50300 45178 50356 45180
rect 50380 45178 50436 45180
rect 50460 45178 50516 45180
rect 50540 45178 50596 45180
rect 50300 45126 50326 45178
rect 50326 45126 50356 45178
rect 50380 45126 50390 45178
rect 50390 45126 50436 45178
rect 50460 45126 50506 45178
rect 50506 45126 50516 45178
rect 50540 45126 50570 45178
rect 50570 45126 50596 45178
rect 50300 45124 50356 45126
rect 50380 45124 50436 45126
rect 50460 45124 50516 45126
rect 50540 45124 50596 45126
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 31114 28872 31170 28928
rect 31298 28736 31354 28792
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 50300 33210 50356 33212
rect 50380 33210 50436 33212
rect 50460 33210 50516 33212
rect 50540 33210 50596 33212
rect 50300 33158 50326 33210
rect 50326 33158 50356 33210
rect 50380 33158 50390 33210
rect 50390 33158 50436 33210
rect 50460 33158 50506 33210
rect 50506 33158 50516 33210
rect 50540 33158 50570 33210
rect 50570 33158 50596 33210
rect 50300 33156 50356 33158
rect 50380 33156 50436 33158
rect 50460 33156 50516 33158
rect 50540 33156 50596 33158
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 50300 32122 50356 32124
rect 50380 32122 50436 32124
rect 50460 32122 50516 32124
rect 50540 32122 50596 32124
rect 50300 32070 50326 32122
rect 50326 32070 50356 32122
rect 50380 32070 50390 32122
rect 50390 32070 50436 32122
rect 50460 32070 50506 32122
rect 50506 32070 50516 32122
rect 50540 32070 50570 32122
rect 50570 32070 50596 32122
rect 50300 32068 50356 32070
rect 50380 32068 50436 32070
rect 50460 32068 50516 32070
rect 50540 32068 50596 32070
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 50300 31034 50356 31036
rect 50380 31034 50436 31036
rect 50460 31034 50516 31036
rect 50540 31034 50596 31036
rect 50300 30982 50326 31034
rect 50326 30982 50356 31034
rect 50380 30982 50390 31034
rect 50390 30982 50436 31034
rect 50460 30982 50506 31034
rect 50506 30982 50516 31034
rect 50540 30982 50570 31034
rect 50570 30982 50596 31034
rect 50300 30980 50356 30982
rect 50380 30980 50436 30982
rect 50460 30980 50516 30982
rect 50540 30980 50596 30982
rect 31574 28872 31630 28928
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 50300 29946 50356 29948
rect 50380 29946 50436 29948
rect 50460 29946 50516 29948
rect 50540 29946 50596 29948
rect 50300 29894 50326 29946
rect 50326 29894 50356 29946
rect 50380 29894 50390 29946
rect 50390 29894 50436 29946
rect 50460 29894 50506 29946
rect 50506 29894 50516 29946
rect 50540 29894 50570 29946
rect 50570 29894 50596 29946
rect 50300 29892 50356 29894
rect 50380 29892 50436 29894
rect 50460 29892 50516 29894
rect 50540 29892 50596 29894
rect 33322 28736 33378 28792
rect 30838 22108 30840 22128
rect 30840 22108 30892 22128
rect 30892 22108 30894 22128
rect 30838 22072 30894 22108
rect 31482 24248 31538 24304
rect 31390 23060 31392 23080
rect 31392 23060 31444 23080
rect 31444 23060 31446 23080
rect 31390 23024 31446 23060
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34334 27956 34336 27976
rect 34336 27956 34388 27976
rect 34388 27956 34390 27976
rect 34334 27920 34390 27956
rect 33506 26868 33508 26888
rect 33508 26868 33560 26888
rect 33560 26868 33562 26888
rect 33506 26832 33562 26868
rect 32494 20984 32550 21040
rect 34426 23044 34482 23080
rect 34426 23024 34428 23044
rect 34428 23024 34480 23044
rect 34480 23024 34482 23044
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 50300 28858 50356 28860
rect 50380 28858 50436 28860
rect 50460 28858 50516 28860
rect 50540 28858 50596 28860
rect 50300 28806 50326 28858
rect 50326 28806 50356 28858
rect 50380 28806 50390 28858
rect 50390 28806 50436 28858
rect 50460 28806 50506 28858
rect 50506 28806 50516 28858
rect 50540 28806 50570 28858
rect 50570 28806 50596 28858
rect 50300 28804 50356 28806
rect 50380 28804 50436 28806
rect 50460 28804 50516 28806
rect 50540 28804 50596 28806
rect 36450 28056 36506 28112
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34334 21004 34390 21040
rect 34334 20984 34336 21004
rect 34336 20984 34388 21004
rect 34388 20984 34390 21004
rect 50300 27770 50356 27772
rect 50380 27770 50436 27772
rect 50460 27770 50516 27772
rect 50540 27770 50596 27772
rect 50300 27718 50326 27770
rect 50326 27718 50356 27770
rect 50380 27718 50390 27770
rect 50390 27718 50436 27770
rect 50460 27718 50506 27770
rect 50506 27718 50516 27770
rect 50540 27718 50570 27770
rect 50570 27718 50596 27770
rect 50300 27716 50356 27718
rect 50380 27716 50436 27718
rect 50460 27716 50516 27718
rect 50540 27716 50596 27718
rect 50300 26682 50356 26684
rect 50380 26682 50436 26684
rect 50460 26682 50516 26684
rect 50540 26682 50596 26684
rect 50300 26630 50326 26682
rect 50326 26630 50356 26682
rect 50380 26630 50390 26682
rect 50390 26630 50436 26682
rect 50460 26630 50506 26682
rect 50506 26630 50516 26682
rect 50540 26630 50570 26682
rect 50570 26630 50596 26682
rect 50300 26628 50356 26630
rect 50380 26628 50436 26630
rect 50460 26628 50516 26630
rect 50540 26628 50596 26630
rect 50300 25594 50356 25596
rect 50380 25594 50436 25596
rect 50460 25594 50516 25596
rect 50540 25594 50596 25596
rect 50300 25542 50326 25594
rect 50326 25542 50356 25594
rect 50380 25542 50390 25594
rect 50390 25542 50436 25594
rect 50460 25542 50506 25594
rect 50506 25542 50516 25594
rect 50540 25542 50570 25594
rect 50570 25542 50596 25594
rect 50300 25540 50356 25542
rect 50380 25540 50436 25542
rect 50460 25540 50516 25542
rect 50540 25540 50596 25542
rect 50300 24506 50356 24508
rect 50380 24506 50436 24508
rect 50460 24506 50516 24508
rect 50540 24506 50596 24508
rect 50300 24454 50326 24506
rect 50326 24454 50356 24506
rect 50380 24454 50390 24506
rect 50390 24454 50436 24506
rect 50460 24454 50506 24506
rect 50506 24454 50516 24506
rect 50540 24454 50570 24506
rect 50570 24454 50596 24506
rect 50300 24452 50356 24454
rect 50380 24452 50436 24454
rect 50460 24452 50516 24454
rect 50540 24452 50596 24454
rect 50300 23418 50356 23420
rect 50380 23418 50436 23420
rect 50460 23418 50516 23420
rect 50540 23418 50596 23420
rect 50300 23366 50326 23418
rect 50326 23366 50356 23418
rect 50380 23366 50390 23418
rect 50390 23366 50436 23418
rect 50460 23366 50506 23418
rect 50506 23366 50516 23418
rect 50540 23366 50570 23418
rect 50570 23366 50596 23418
rect 50300 23364 50356 23366
rect 50380 23364 50436 23366
rect 50460 23364 50516 23366
rect 50540 23364 50596 23366
rect 55218 56480 55274 56536
rect 55678 59064 55734 59120
rect 56414 58520 56470 58576
rect 56506 58248 56562 58304
rect 56506 58012 56508 58032
rect 56508 58012 56560 58032
rect 56560 58012 56562 58032
rect 56506 57976 56562 58012
rect 55586 54848 55642 54904
rect 57058 56924 57060 56944
rect 57060 56924 57112 56944
rect 57112 56924 57114 56944
rect 57058 56888 57114 56924
rect 56506 53352 56562 53408
rect 56506 51720 56562 51776
rect 56506 48628 56508 48648
rect 56508 48628 56560 48648
rect 56560 48628 56562 48648
rect 56506 48592 56562 48628
rect 55310 34584 55366 34640
rect 55218 32952 55274 33008
rect 56506 45464 56562 45520
rect 56506 43968 56562 44024
rect 56506 42336 56562 42392
rect 56506 40840 56562 40896
rect 56506 37748 56508 37768
rect 56508 37748 56560 37768
rect 56560 37748 56562 37768
rect 56506 37712 56562 37748
rect 56230 36080 56286 36136
rect 56506 31456 56562 31512
rect 56506 29824 56562 29880
rect 55586 28328 55642 28384
rect 55586 26696 55642 26752
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 50300 22330 50356 22332
rect 50380 22330 50436 22332
rect 50460 22330 50516 22332
rect 50540 22330 50596 22332
rect 50300 22278 50326 22330
rect 50326 22278 50356 22330
rect 50380 22278 50390 22330
rect 50390 22278 50436 22330
rect 50460 22278 50506 22330
rect 50506 22278 50516 22330
rect 50540 22278 50570 22330
rect 50570 22278 50596 22330
rect 50300 22276 50356 22278
rect 50380 22276 50436 22278
rect 50460 22276 50516 22278
rect 50540 22276 50596 22278
rect 36266 22092 36322 22128
rect 36266 22072 36268 22092
rect 36268 22072 36320 22092
rect 36320 22072 36322 22092
rect 50300 21242 50356 21244
rect 50380 21242 50436 21244
rect 50460 21242 50516 21244
rect 50540 21242 50596 21244
rect 50300 21190 50326 21242
rect 50326 21190 50356 21242
rect 50380 21190 50390 21242
rect 50390 21190 50436 21242
rect 50460 21190 50506 21242
rect 50506 21190 50516 21242
rect 50540 21190 50570 21242
rect 50570 21190 50596 21242
rect 50300 21188 50356 21190
rect 50380 21188 50436 21190
rect 50460 21188 50516 21190
rect 50540 21188 50596 21190
rect 50300 20154 50356 20156
rect 50380 20154 50436 20156
rect 50460 20154 50516 20156
rect 50540 20154 50596 20156
rect 50300 20102 50326 20154
rect 50326 20102 50356 20154
rect 50380 20102 50390 20154
rect 50390 20102 50436 20154
rect 50460 20102 50506 20154
rect 50506 20102 50516 20154
rect 50540 20102 50570 20154
rect 50570 20102 50596 20154
rect 50300 20100 50356 20102
rect 50380 20100 50436 20102
rect 50460 20100 50516 20102
rect 50540 20100 50596 20102
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 50300 19066 50356 19068
rect 50380 19066 50436 19068
rect 50460 19066 50516 19068
rect 50540 19066 50596 19068
rect 50300 19014 50326 19066
rect 50326 19014 50356 19066
rect 50380 19014 50390 19066
rect 50390 19014 50436 19066
rect 50460 19014 50506 19066
rect 50506 19014 50516 19066
rect 50540 19014 50570 19066
rect 50570 19014 50596 19066
rect 50300 19012 50356 19014
rect 50380 19012 50436 19014
rect 50460 19012 50516 19014
rect 50540 19012 50596 19014
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 50300 17978 50356 17980
rect 50380 17978 50436 17980
rect 50460 17978 50516 17980
rect 50540 17978 50596 17980
rect 50300 17926 50326 17978
rect 50326 17926 50356 17978
rect 50380 17926 50390 17978
rect 50390 17926 50436 17978
rect 50460 17926 50506 17978
rect 50506 17926 50516 17978
rect 50540 17926 50570 17978
rect 50570 17926 50596 17978
rect 50300 17924 50356 17926
rect 50380 17924 50436 17926
rect 50460 17924 50516 17926
rect 50540 17924 50596 17926
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 50300 16890 50356 16892
rect 50380 16890 50436 16892
rect 50460 16890 50516 16892
rect 50540 16890 50596 16892
rect 50300 16838 50326 16890
rect 50326 16838 50356 16890
rect 50380 16838 50390 16890
rect 50390 16838 50436 16890
rect 50460 16838 50506 16890
rect 50506 16838 50516 16890
rect 50540 16838 50570 16890
rect 50570 16838 50596 16890
rect 50300 16836 50356 16838
rect 50380 16836 50436 16838
rect 50460 16836 50516 16838
rect 50540 16836 50596 16838
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 50300 15802 50356 15804
rect 50380 15802 50436 15804
rect 50460 15802 50516 15804
rect 50540 15802 50596 15804
rect 50300 15750 50326 15802
rect 50326 15750 50356 15802
rect 50380 15750 50390 15802
rect 50390 15750 50436 15802
rect 50460 15750 50506 15802
rect 50506 15750 50516 15802
rect 50540 15750 50570 15802
rect 50570 15750 50596 15802
rect 50300 15748 50356 15750
rect 50380 15748 50436 15750
rect 50460 15748 50516 15750
rect 50540 15748 50596 15750
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 50300 14714 50356 14716
rect 50380 14714 50436 14716
rect 50460 14714 50516 14716
rect 50540 14714 50596 14716
rect 50300 14662 50326 14714
rect 50326 14662 50356 14714
rect 50380 14662 50390 14714
rect 50390 14662 50436 14714
rect 50460 14662 50506 14714
rect 50506 14662 50516 14714
rect 50540 14662 50570 14714
rect 50570 14662 50596 14714
rect 50300 14660 50356 14662
rect 50380 14660 50436 14662
rect 50460 14660 50516 14662
rect 50540 14660 50596 14662
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 50300 13626 50356 13628
rect 50380 13626 50436 13628
rect 50460 13626 50516 13628
rect 50540 13626 50596 13628
rect 50300 13574 50326 13626
rect 50326 13574 50356 13626
rect 50380 13574 50390 13626
rect 50390 13574 50436 13626
rect 50460 13574 50506 13626
rect 50506 13574 50516 13626
rect 50540 13574 50570 13626
rect 50570 13574 50596 13626
rect 50300 13572 50356 13574
rect 50380 13572 50436 13574
rect 50460 13572 50516 13574
rect 50540 13572 50596 13574
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 50300 12538 50356 12540
rect 50380 12538 50436 12540
rect 50460 12538 50516 12540
rect 50540 12538 50596 12540
rect 50300 12486 50326 12538
rect 50326 12486 50356 12538
rect 50380 12486 50390 12538
rect 50390 12486 50436 12538
rect 50460 12486 50506 12538
rect 50506 12486 50516 12538
rect 50540 12486 50570 12538
rect 50570 12486 50596 12538
rect 50300 12484 50356 12486
rect 50380 12484 50436 12486
rect 50460 12484 50516 12486
rect 50540 12484 50596 12486
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 50300 11450 50356 11452
rect 50380 11450 50436 11452
rect 50460 11450 50516 11452
rect 50540 11450 50596 11452
rect 50300 11398 50326 11450
rect 50326 11398 50356 11450
rect 50380 11398 50390 11450
rect 50390 11398 50436 11450
rect 50460 11398 50506 11450
rect 50506 11398 50516 11450
rect 50540 11398 50570 11450
rect 50570 11398 50596 11450
rect 50300 11396 50356 11398
rect 50380 11396 50436 11398
rect 50460 11396 50516 11398
rect 50540 11396 50596 11398
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 50300 10362 50356 10364
rect 50380 10362 50436 10364
rect 50460 10362 50516 10364
rect 50540 10362 50596 10364
rect 50300 10310 50326 10362
rect 50326 10310 50356 10362
rect 50380 10310 50390 10362
rect 50390 10310 50436 10362
rect 50460 10310 50506 10362
rect 50506 10310 50516 10362
rect 50540 10310 50570 10362
rect 50570 10310 50596 10362
rect 50300 10308 50356 10310
rect 50380 10308 50436 10310
rect 50460 10308 50516 10310
rect 50540 10308 50596 10310
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 50300 9274 50356 9276
rect 50380 9274 50436 9276
rect 50460 9274 50516 9276
rect 50540 9274 50596 9276
rect 50300 9222 50326 9274
rect 50326 9222 50356 9274
rect 50380 9222 50390 9274
rect 50390 9222 50436 9274
rect 50460 9222 50506 9274
rect 50506 9222 50516 9274
rect 50540 9222 50570 9274
rect 50570 9222 50596 9274
rect 50300 9220 50356 9222
rect 50380 9220 50436 9222
rect 50460 9220 50516 9222
rect 50540 9220 50596 9222
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 50300 8186 50356 8188
rect 50380 8186 50436 8188
rect 50460 8186 50516 8188
rect 50540 8186 50596 8188
rect 50300 8134 50326 8186
rect 50326 8134 50356 8186
rect 50380 8134 50390 8186
rect 50390 8134 50436 8186
rect 50460 8134 50506 8186
rect 50506 8134 50516 8186
rect 50540 8134 50570 8186
rect 50570 8134 50596 8186
rect 50300 8132 50356 8134
rect 50380 8132 50436 8134
rect 50460 8132 50516 8134
rect 50540 8132 50596 8134
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 50300 7098 50356 7100
rect 50380 7098 50436 7100
rect 50460 7098 50516 7100
rect 50540 7098 50596 7100
rect 50300 7046 50326 7098
rect 50326 7046 50356 7098
rect 50380 7046 50390 7098
rect 50390 7046 50436 7098
rect 50460 7046 50506 7098
rect 50506 7046 50516 7098
rect 50540 7046 50570 7098
rect 50570 7046 50596 7098
rect 50300 7044 50356 7046
rect 50380 7044 50436 7046
rect 50460 7044 50516 7046
rect 50540 7044 50596 7046
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 50300 6010 50356 6012
rect 50380 6010 50436 6012
rect 50460 6010 50516 6012
rect 50540 6010 50596 6012
rect 50300 5958 50326 6010
rect 50326 5958 50356 6010
rect 50380 5958 50390 6010
rect 50390 5958 50436 6010
rect 50460 5958 50506 6010
rect 50506 5958 50516 6010
rect 50540 5958 50570 6010
rect 50570 5958 50596 6010
rect 50300 5956 50356 5958
rect 50380 5956 50436 5958
rect 50460 5956 50516 5958
rect 50540 5956 50596 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 55586 18944 55642 19000
rect 55586 15816 55642 15872
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 50300 4922 50356 4924
rect 50380 4922 50436 4924
rect 50460 4922 50516 4924
rect 50540 4922 50596 4924
rect 50300 4870 50326 4922
rect 50326 4870 50356 4922
rect 50380 4870 50390 4922
rect 50390 4870 50436 4922
rect 50460 4870 50506 4922
rect 50506 4870 50516 4922
rect 50540 4870 50570 4922
rect 50570 4870 50596 4922
rect 50300 4868 50356 4870
rect 50380 4868 50436 4870
rect 50460 4868 50516 4870
rect 50540 4868 50596 4870
rect 50300 3834 50356 3836
rect 50380 3834 50436 3836
rect 50460 3834 50516 3836
rect 50540 3834 50596 3836
rect 50300 3782 50326 3834
rect 50326 3782 50356 3834
rect 50380 3782 50390 3834
rect 50390 3782 50436 3834
rect 50460 3782 50506 3834
rect 50506 3782 50516 3834
rect 50540 3782 50570 3834
rect 50570 3782 50596 3834
rect 50300 3780 50356 3782
rect 50380 3780 50436 3782
rect 50460 3780 50516 3782
rect 50540 3780 50596 3782
rect 50300 2746 50356 2748
rect 50380 2746 50436 2748
rect 50460 2746 50516 2748
rect 50540 2746 50596 2748
rect 50300 2694 50326 2746
rect 50326 2694 50356 2746
rect 50380 2694 50390 2746
rect 50390 2694 50436 2746
rect 50460 2694 50506 2746
rect 50506 2694 50516 2746
rect 50540 2694 50570 2746
rect 50570 2694 50596 2746
rect 50300 2692 50356 2694
rect 50380 2692 50436 2694
rect 50460 2692 50516 2694
rect 50540 2692 50596 2694
rect 2870 448 2926 504
rect 55586 14184 55642 14240
rect 56230 17312 56286 17368
rect 56506 25200 56562 25256
rect 56506 23604 56508 23624
rect 56508 23604 56560 23624
rect 56560 23604 56562 23624
rect 56506 23568 56562 23604
rect 56506 20440 56562 20496
rect 56966 53780 57022 53816
rect 56966 53760 56968 53780
rect 56968 53760 57020 53780
rect 57020 53760 57022 53780
rect 57058 49156 57114 49192
rect 57058 49136 57060 49156
rect 57060 49136 57112 49156
rect 57112 49136 57114 49156
rect 56874 47116 56930 47152
rect 56874 47096 56876 47116
rect 56876 47096 56928 47116
rect 56928 47096 56930 47116
rect 57058 42880 57114 42936
rect 57058 36644 57114 36680
rect 57058 36624 57060 36644
rect 57060 36624 57112 36644
rect 57112 36624 57114 36644
rect 57058 33516 57114 33552
rect 57058 33496 57060 33516
rect 57060 33496 57112 33516
rect 57112 33496 57114 33516
rect 58162 57452 58218 57488
rect 58162 57432 58164 57452
rect 58164 57432 58216 57452
rect 58216 57432 58218 57452
rect 58162 55936 58218 55992
rect 57334 55412 57390 55448
rect 57334 55392 57336 55412
rect 57336 55392 57388 55412
rect 57388 55392 57390 55412
rect 58162 54304 58218 54360
rect 57242 50224 57298 50280
rect 57334 41268 57390 41304
rect 57334 41248 57336 41268
rect 57336 41248 57388 41268
rect 57388 41248 57390 41268
rect 56966 31884 57022 31920
rect 56966 31864 56968 31884
rect 56968 31864 57020 31884
rect 57020 31864 57022 31884
rect 57058 30912 57114 30968
rect 57150 30368 57206 30424
rect 56966 28600 57022 28656
rect 56966 27276 56968 27296
rect 56968 27276 57020 27296
rect 57020 27276 57022 27296
rect 56966 27240 57022 27276
rect 57058 22500 57114 22536
rect 57058 22480 57060 22500
rect 57060 22480 57112 22500
rect 57112 22480 57114 22500
rect 58162 52808 58218 52864
rect 58162 52264 58218 52320
rect 58162 51176 58218 51232
rect 58162 50632 58218 50688
rect 58162 49716 58164 49736
rect 58164 49716 58216 49736
rect 58216 49716 58218 49736
rect 58162 49680 58218 49716
rect 57886 48048 57942 48104
rect 58162 47524 58218 47560
rect 58162 47504 58164 47524
rect 58164 47504 58216 47524
rect 58216 47504 58218 47524
rect 58162 46572 58218 46608
rect 58162 46552 58164 46572
rect 58164 46552 58216 46572
rect 58216 46552 58218 46572
rect 58162 46008 58218 46064
rect 58162 44940 58218 44976
rect 58162 44920 58164 44940
rect 58164 44920 58216 44940
rect 58216 44920 58218 44940
rect 58162 44376 58218 44432
rect 58162 43424 58218 43480
rect 58162 41792 58218 41848
rect 58162 40296 58218 40352
rect 58162 39752 58218 39808
rect 57978 39208 58034 39264
rect 58162 38664 58218 38720
rect 58162 38120 58218 38176
rect 57886 37168 57942 37224
rect 57886 35536 57942 35592
rect 57886 34040 57942 34096
rect 58162 35012 58218 35048
rect 58162 34992 58164 35012
rect 58164 34992 58216 35012
rect 58216 34992 58218 35012
rect 58530 32444 58532 32464
rect 58532 32444 58584 32464
rect 58584 32444 58586 32464
rect 58530 32408 58586 32444
rect 58162 29280 58218 29336
rect 58162 28736 58218 28792
rect 57886 28464 57942 28520
rect 58162 27784 58218 27840
rect 58346 26152 58402 26208
rect 58162 25608 58218 25664
rect 58162 24656 58218 24712
rect 58162 24112 58218 24168
rect 57334 22072 57390 22128
rect 58162 23044 58218 23080
rect 58162 23024 58164 23044
rect 58164 23024 58216 23044
rect 58216 23024 58218 23044
rect 58162 21528 58218 21584
rect 58162 21004 58218 21040
rect 58162 20984 58164 21004
rect 58164 20984 58216 21004
rect 58216 20984 58218 21004
rect 58162 19916 58218 19952
rect 58162 19896 58164 19916
rect 58164 19896 58216 19916
rect 58216 19896 58218 19916
rect 58162 19352 58218 19408
rect 58162 18400 58218 18456
rect 58162 17856 58218 17912
rect 56966 14728 57022 14784
rect 55402 12724 55404 12744
rect 55404 12724 55456 12744
rect 55456 12724 55458 12744
rect 55402 12688 55458 12724
rect 55586 11056 55642 11112
rect 55586 9560 55642 9616
rect 56506 11600 56562 11656
rect 55678 7928 55734 7984
rect 55218 4800 55274 4856
rect 55126 3304 55182 3360
rect 55494 6432 55550 6488
rect 55494 6316 55550 6352
rect 55494 6296 55496 6316
rect 55496 6296 55548 6316
rect 55548 6296 55550 6316
rect 56414 6840 56470 6896
rect 57334 13096 57390 13152
rect 58162 16768 58218 16824
rect 58254 16224 58310 16280
rect 58070 15272 58126 15328
rect 58070 13640 58126 13696
rect 57886 12144 57942 12200
rect 57886 10512 57942 10568
rect 58162 9988 58218 10024
rect 58162 9968 58164 9988
rect 58164 9968 58216 9988
rect 58216 9968 58218 9988
rect 58162 9016 58218 9072
rect 57426 8492 57482 8528
rect 57426 8472 57428 8492
rect 57428 8472 57480 8492
rect 57480 8472 57482 8492
rect 56598 6332 56600 6352
rect 56600 6332 56652 6352
rect 56652 6332 56654 6352
rect 56598 6296 56654 6332
rect 56966 4256 57022 4312
rect 57058 3712 57114 3768
rect 55954 2216 56010 2272
rect 58162 7384 58218 7440
rect 56506 1708 56508 1728
rect 56508 1708 56560 1728
rect 56560 1708 56562 1728
rect 56506 1672 56562 1708
rect 55586 584 55642 640
rect 58162 5888 58218 5944
rect 57886 5344 57942 5400
rect 58162 2760 58218 2816
rect 57886 1128 57942 1184
rect 56322 176 56378 232
<< metal3 >>
rect 56501 59666 56567 59669
rect 59200 59666 60000 59696
rect 56501 59664 60000 59666
rect 56501 59608 56506 59664
rect 56562 59608 60000 59664
rect 56501 59606 60000 59608
rect 56501 59603 56567 59606
rect 59200 59576 60000 59606
rect 0 59530 800 59560
rect 2773 59530 2839 59533
rect 0 59528 2839 59530
rect 0 59472 2778 59528
rect 2834 59472 2839 59528
rect 0 59470 2839 59472
rect 0 59440 800 59470
rect 2773 59467 2839 59470
rect 55673 59122 55739 59125
rect 59200 59122 60000 59152
rect 55673 59120 60000 59122
rect 55673 59064 55678 59120
rect 55734 59064 60000 59120
rect 55673 59062 60000 59064
rect 55673 59059 55739 59062
rect 59200 59032 60000 59062
rect 0 58578 800 58608
rect 1209 58578 1275 58581
rect 0 58576 1275 58578
rect 0 58520 1214 58576
rect 1270 58520 1275 58576
rect 0 58518 1275 58520
rect 0 58488 800 58518
rect 1209 58515 1275 58518
rect 56409 58578 56475 58581
rect 59200 58578 60000 58608
rect 56409 58576 60000 58578
rect 56409 58520 56414 58576
rect 56470 58520 60000 58576
rect 56409 58518 60000 58520
rect 56409 58515 56475 58518
rect 59200 58488 60000 58518
rect 55121 58306 55187 58309
rect 56501 58306 56567 58309
rect 55121 58304 56567 58306
rect 55121 58248 55126 58304
rect 55182 58248 56506 58304
rect 56562 58248 56567 58304
rect 55121 58246 56567 58248
rect 55121 58243 55187 58246
rect 56501 58243 56567 58246
rect 56501 58034 56567 58037
rect 59200 58034 60000 58064
rect 56501 58032 60000 58034
rect 56501 57976 56506 58032
rect 56562 57976 60000 58032
rect 56501 57974 60000 57976
rect 56501 57971 56567 57974
rect 59200 57944 60000 57974
rect 4208 57696 4528 57697
rect 0 57626 800 57656
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 2129 57626 2195 57629
rect 0 57624 2195 57626
rect 0 57568 2134 57624
rect 2190 57568 2195 57624
rect 0 57566 2195 57568
rect 0 57536 800 57566
rect 2129 57563 2195 57566
rect 25589 57626 25655 57629
rect 29269 57626 29335 57629
rect 25589 57624 29335 57626
rect 25589 57568 25594 57624
rect 25650 57568 29274 57624
rect 29330 57568 29335 57624
rect 25589 57566 29335 57568
rect 25589 57563 25655 57566
rect 29269 57563 29335 57566
rect 58157 57490 58223 57493
rect 59200 57490 60000 57520
rect 58157 57488 60000 57490
rect 58157 57432 58162 57488
rect 58218 57432 60000 57488
rect 58157 57430 60000 57432
rect 58157 57427 58223 57430
rect 59200 57400 60000 57430
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 57087 19888 57088
rect 50288 57152 50608 57153
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 57087 50608 57088
rect 28349 57082 28415 57085
rect 29269 57082 29335 57085
rect 28349 57080 29335 57082
rect 28349 57024 28354 57080
rect 28410 57024 29274 57080
rect 29330 57024 29335 57080
rect 28349 57022 29335 57024
rect 28349 57019 28415 57022
rect 29269 57019 29335 57022
rect 31109 57082 31175 57085
rect 35617 57082 35683 57085
rect 31109 57080 35683 57082
rect 31109 57024 31114 57080
rect 31170 57024 35622 57080
rect 35678 57024 35683 57080
rect 31109 57022 35683 57024
rect 31109 57019 31175 57022
rect 35617 57019 35683 57022
rect 29545 56946 29611 56949
rect 35893 56946 35959 56949
rect 29545 56944 35959 56946
rect 29545 56888 29550 56944
rect 29606 56888 35898 56944
rect 35954 56888 35959 56944
rect 29545 56886 35959 56888
rect 29545 56883 29611 56886
rect 35893 56883 35959 56886
rect 57053 56946 57119 56949
rect 59200 56946 60000 56976
rect 57053 56944 60000 56946
rect 57053 56888 57058 56944
rect 57114 56888 60000 56944
rect 57053 56886 60000 56888
rect 57053 56883 57119 56886
rect 59200 56856 60000 56886
rect 29085 56810 29151 56813
rect 29637 56810 29703 56813
rect 29085 56808 29703 56810
rect 29085 56752 29090 56808
rect 29146 56752 29642 56808
rect 29698 56752 29703 56808
rect 29085 56750 29703 56752
rect 29085 56747 29151 56750
rect 29637 56747 29703 56750
rect 0 56674 800 56704
rect 1393 56674 1459 56677
rect 0 56672 1459 56674
rect 0 56616 1398 56672
rect 1454 56616 1459 56672
rect 0 56614 1459 56616
rect 0 56584 800 56614
rect 1393 56611 1459 56614
rect 4208 56608 4528 56609
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 55213 56538 55279 56541
rect 59200 56538 60000 56568
rect 55213 56536 60000 56538
rect 55213 56480 55218 56536
rect 55274 56480 60000 56536
rect 55213 56478 60000 56480
rect 55213 56475 55279 56478
rect 59200 56448 60000 56478
rect 32949 56402 33015 56405
rect 34973 56402 35039 56405
rect 32949 56400 35039 56402
rect 32949 56344 32954 56400
rect 33010 56344 34978 56400
rect 35034 56344 35039 56400
rect 32949 56342 35039 56344
rect 32949 56339 33015 56342
rect 34973 56339 35039 56342
rect 33041 56266 33107 56269
rect 36077 56266 36143 56269
rect 33041 56264 36143 56266
rect 33041 56208 33046 56264
rect 33102 56208 36082 56264
rect 36138 56208 36143 56264
rect 33041 56206 36143 56208
rect 33041 56203 33107 56206
rect 36077 56203 36143 56206
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect 50288 56064 50608 56065
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 55999 50608 56000
rect 58157 55994 58223 55997
rect 59200 55994 60000 56024
rect 58157 55992 60000 55994
rect 58157 55936 58162 55992
rect 58218 55936 60000 55992
rect 58157 55934 60000 55936
rect 58157 55931 58223 55934
rect 59200 55904 60000 55934
rect 0 55858 800 55888
rect 1393 55858 1459 55861
rect 0 55856 1459 55858
rect 0 55800 1398 55856
rect 1454 55800 1459 55856
rect 0 55798 1459 55800
rect 0 55768 800 55798
rect 1393 55795 1459 55798
rect 31937 55858 32003 55861
rect 36445 55858 36511 55861
rect 31937 55856 36511 55858
rect 31937 55800 31942 55856
rect 31998 55800 36450 55856
rect 36506 55800 36511 55856
rect 31937 55798 36511 55800
rect 31937 55795 32003 55798
rect 36445 55795 36511 55798
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 57329 55450 57395 55453
rect 59200 55450 60000 55480
rect 57329 55448 60000 55450
rect 57329 55392 57334 55448
rect 57390 55392 60000 55448
rect 57329 55390 60000 55392
rect 57329 55387 57395 55390
rect 59200 55360 60000 55390
rect 19568 54976 19888 54977
rect 0 54906 800 54936
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 50288 54976 50608 54977
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 54911 50608 54912
rect 1393 54906 1459 54909
rect 0 54904 1459 54906
rect 0 54848 1398 54904
rect 1454 54848 1459 54904
rect 0 54846 1459 54848
rect 0 54816 800 54846
rect 1393 54843 1459 54846
rect 55581 54906 55647 54909
rect 59200 54906 60000 54936
rect 55581 54904 60000 54906
rect 55581 54848 55586 54904
rect 55642 54848 60000 54904
rect 55581 54846 60000 54848
rect 55581 54843 55647 54846
rect 59200 54816 60000 54846
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 54367 35248 54368
rect 58157 54362 58223 54365
rect 59200 54362 60000 54392
rect 58157 54360 60000 54362
rect 58157 54304 58162 54360
rect 58218 54304 60000 54360
rect 58157 54302 60000 54304
rect 58157 54299 58223 54302
rect 59200 54272 60000 54302
rect 0 53954 800 53984
rect 1393 53954 1459 53957
rect 0 53952 1459 53954
rect 0 53896 1398 53952
rect 1454 53896 1459 53952
rect 0 53894 1459 53896
rect 0 53864 800 53894
rect 1393 53891 1459 53894
rect 19568 53888 19888 53889
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 50288 53888 50608 53889
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 53823 50608 53824
rect 56961 53818 57027 53821
rect 59200 53818 60000 53848
rect 56961 53816 60000 53818
rect 56961 53760 56966 53816
rect 57022 53760 60000 53816
rect 56961 53758 60000 53760
rect 56961 53755 57027 53758
rect 59200 53728 60000 53758
rect 56501 53410 56567 53413
rect 59200 53410 60000 53440
rect 56501 53408 60000 53410
rect 56501 53352 56506 53408
rect 56562 53352 60000 53408
rect 56501 53350 60000 53352
rect 56501 53347 56567 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 59200 53320 60000 53350
rect 34928 53279 35248 53280
rect 0 53002 800 53032
rect 1393 53002 1459 53005
rect 0 53000 1459 53002
rect 0 52944 1398 53000
rect 1454 52944 1459 53000
rect 0 52942 1459 52944
rect 0 52912 800 52942
rect 1393 52939 1459 52942
rect 31937 53002 32003 53005
rect 34697 53002 34763 53005
rect 31937 53000 34763 53002
rect 31937 52944 31942 53000
rect 31998 52944 34702 53000
rect 34758 52944 34763 53000
rect 31937 52942 34763 52944
rect 31937 52939 32003 52942
rect 34697 52939 34763 52942
rect 58157 52866 58223 52869
rect 59200 52866 60000 52896
rect 58157 52864 60000 52866
rect 58157 52808 58162 52864
rect 58218 52808 60000 52864
rect 58157 52806 60000 52808
rect 58157 52803 58223 52806
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 50288 52800 50608 52801
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 59200 52776 60000 52806
rect 50288 52735 50608 52736
rect 58157 52322 58223 52325
rect 59200 52322 60000 52352
rect 58157 52320 60000 52322
rect 58157 52264 58162 52320
rect 58218 52264 60000 52320
rect 58157 52262 60000 52264
rect 58157 52259 58223 52262
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 59200 52232 60000 52262
rect 34928 52191 35248 52192
rect 0 52050 800 52080
rect 1393 52050 1459 52053
rect 0 52048 1459 52050
rect 0 51992 1398 52048
rect 1454 51992 1459 52048
rect 0 51990 1459 51992
rect 0 51960 800 51990
rect 1393 51987 1459 51990
rect 56501 51778 56567 51781
rect 59200 51778 60000 51808
rect 56501 51776 60000 51778
rect 56501 51720 56506 51776
rect 56562 51720 60000 51776
rect 56501 51718 60000 51720
rect 56501 51715 56567 51718
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 50288 51712 50608 51713
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 59200 51688 60000 51718
rect 50288 51647 50608 51648
rect 0 51234 800 51264
rect 1393 51234 1459 51237
rect 0 51232 1459 51234
rect 0 51176 1398 51232
rect 1454 51176 1459 51232
rect 0 51174 1459 51176
rect 0 51144 800 51174
rect 1393 51171 1459 51174
rect 58157 51234 58223 51237
rect 59200 51234 60000 51264
rect 58157 51232 60000 51234
rect 58157 51176 58162 51232
rect 58218 51176 60000 51232
rect 58157 51174 60000 51176
rect 58157 51171 58223 51174
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 59200 51144 60000 51174
rect 34928 51103 35248 51104
rect 58157 50690 58223 50693
rect 59200 50690 60000 50720
rect 58157 50688 60000 50690
rect 58157 50632 58162 50688
rect 58218 50632 60000 50688
rect 58157 50630 60000 50632
rect 58157 50627 58223 50630
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 50559 19888 50560
rect 50288 50624 50608 50625
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 59200 50600 60000 50630
rect 50288 50559 50608 50560
rect 0 50282 800 50312
rect 1393 50282 1459 50285
rect 0 50280 1459 50282
rect 0 50224 1398 50280
rect 1454 50224 1459 50280
rect 0 50222 1459 50224
rect 0 50192 800 50222
rect 1393 50219 1459 50222
rect 57237 50282 57303 50285
rect 59200 50282 60000 50312
rect 57237 50280 60000 50282
rect 57237 50224 57242 50280
rect 57298 50224 60000 50280
rect 57237 50222 60000 50224
rect 57237 50219 57303 50222
rect 59200 50192 60000 50222
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 50288 49536 50608 49537
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 49471 50608 49472
rect 0 49330 800 49360
rect 1393 49330 1459 49333
rect 0 49328 1459 49330
rect 0 49272 1398 49328
rect 1454 49272 1459 49328
rect 0 49270 1459 49272
rect 0 49240 800 49270
rect 1393 49267 1459 49270
rect 57053 49194 57119 49197
rect 59200 49194 60000 49224
rect 57053 49192 60000 49194
rect 57053 49136 57058 49192
rect 57114 49136 60000 49192
rect 57053 49134 60000 49136
rect 57053 49131 57119 49134
rect 59200 49104 60000 49134
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 56501 48650 56567 48653
rect 59200 48650 60000 48680
rect 56501 48648 60000 48650
rect 56501 48592 56506 48648
rect 56562 48592 60000 48648
rect 56501 48590 60000 48592
rect 56501 48587 56567 48590
rect 59200 48560 60000 48590
rect 19568 48448 19888 48449
rect 0 48378 800 48408
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 50288 48448 50608 48449
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 48383 50608 48384
rect 1393 48378 1459 48381
rect 0 48376 1459 48378
rect 0 48320 1398 48376
rect 1454 48320 1459 48376
rect 0 48318 1459 48320
rect 0 48288 800 48318
rect 1393 48315 1459 48318
rect 57881 48106 57947 48109
rect 59200 48106 60000 48136
rect 57881 48104 60000 48106
rect 57881 48048 57886 48104
rect 57942 48048 60000 48104
rect 57881 48046 60000 48048
rect 57881 48043 57947 48046
rect 59200 48016 60000 48046
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 0 47562 800 47592
rect 1393 47562 1459 47565
rect 0 47560 1459 47562
rect 0 47504 1398 47560
rect 1454 47504 1459 47560
rect 0 47502 1459 47504
rect 0 47472 800 47502
rect 1393 47499 1459 47502
rect 58157 47562 58223 47565
rect 59200 47562 60000 47592
rect 58157 47560 60000 47562
rect 58157 47504 58162 47560
rect 58218 47504 60000 47560
rect 58157 47502 60000 47504
rect 58157 47499 58223 47502
rect 59200 47472 60000 47502
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 50288 47360 50608 47361
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 47295 50608 47296
rect 56869 47154 56935 47157
rect 59200 47154 60000 47184
rect 56869 47152 60000 47154
rect 56869 47096 56874 47152
rect 56930 47096 60000 47152
rect 56869 47094 60000 47096
rect 56869 47091 56935 47094
rect 59200 47064 60000 47094
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 0 46610 800 46640
rect 1393 46610 1459 46613
rect 0 46608 1459 46610
rect 0 46552 1398 46608
rect 1454 46552 1459 46608
rect 0 46550 1459 46552
rect 0 46520 800 46550
rect 1393 46547 1459 46550
rect 58157 46610 58223 46613
rect 59200 46610 60000 46640
rect 58157 46608 60000 46610
rect 58157 46552 58162 46608
rect 58218 46552 60000 46608
rect 58157 46550 60000 46552
rect 58157 46547 58223 46550
rect 59200 46520 60000 46550
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 50288 46272 50608 46273
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 46207 50608 46208
rect 58157 46066 58223 46069
rect 59200 46066 60000 46096
rect 58157 46064 60000 46066
rect 58157 46008 58162 46064
rect 58218 46008 60000 46064
rect 58157 46006 60000 46008
rect 58157 46003 58223 46006
rect 59200 45976 60000 46006
rect 4208 45728 4528 45729
rect 0 45658 800 45688
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 1393 45658 1459 45661
rect 0 45656 1459 45658
rect 0 45600 1398 45656
rect 1454 45600 1459 45656
rect 0 45598 1459 45600
rect 0 45568 800 45598
rect 1393 45595 1459 45598
rect 56501 45522 56567 45525
rect 59200 45522 60000 45552
rect 56501 45520 60000 45522
rect 56501 45464 56506 45520
rect 56562 45464 60000 45520
rect 56501 45462 60000 45464
rect 56501 45459 56567 45462
rect 59200 45432 60000 45462
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 50288 45184 50608 45185
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 45119 50608 45120
rect 58157 44978 58223 44981
rect 59200 44978 60000 45008
rect 58157 44976 60000 44978
rect 58157 44920 58162 44976
rect 58218 44920 60000 44976
rect 58157 44918 60000 44920
rect 58157 44915 58223 44918
rect 59200 44888 60000 44918
rect 0 44706 800 44736
rect 1393 44706 1459 44709
rect 0 44704 1459 44706
rect 0 44648 1398 44704
rect 1454 44648 1459 44704
rect 0 44646 1459 44648
rect 0 44616 800 44646
rect 1393 44643 1459 44646
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 58157 44434 58223 44437
rect 59200 44434 60000 44464
rect 58157 44432 60000 44434
rect 58157 44376 58162 44432
rect 58218 44376 60000 44432
rect 58157 44374 60000 44376
rect 58157 44371 58223 44374
rect 59200 44344 60000 44374
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 56501 44026 56567 44029
rect 59200 44026 60000 44056
rect 56501 44024 60000 44026
rect 56501 43968 56506 44024
rect 56562 43968 60000 44024
rect 56501 43966 60000 43968
rect 56501 43963 56567 43966
rect 59200 43936 60000 43966
rect 0 43754 800 43784
rect 1393 43754 1459 43757
rect 0 43752 1459 43754
rect 0 43696 1398 43752
rect 1454 43696 1459 43752
rect 0 43694 1459 43696
rect 0 43664 800 43694
rect 1393 43691 1459 43694
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 58157 43482 58223 43485
rect 59200 43482 60000 43512
rect 58157 43480 60000 43482
rect 58157 43424 58162 43480
rect 58218 43424 60000 43480
rect 58157 43422 60000 43424
rect 58157 43419 58223 43422
rect 59200 43392 60000 43422
rect 19568 43008 19888 43009
rect 0 42938 800 42968
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42848 800 42878
rect 1393 42875 1459 42878
rect 57053 42938 57119 42941
rect 59200 42938 60000 42968
rect 57053 42936 60000 42938
rect 57053 42880 57058 42936
rect 57114 42880 60000 42936
rect 57053 42878 60000 42880
rect 57053 42875 57119 42878
rect 59200 42848 60000 42878
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 56501 42394 56567 42397
rect 59200 42394 60000 42424
rect 56501 42392 60000 42394
rect 56501 42336 56506 42392
rect 56562 42336 60000 42392
rect 56501 42334 60000 42336
rect 56501 42331 56567 42334
rect 59200 42304 60000 42334
rect 0 41986 800 42016
rect 1393 41986 1459 41989
rect 0 41984 1459 41986
rect 0 41928 1398 41984
rect 1454 41928 1459 41984
rect 0 41926 1459 41928
rect 0 41896 800 41926
rect 1393 41923 1459 41926
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 58157 41850 58223 41853
rect 59200 41850 60000 41880
rect 58157 41848 60000 41850
rect 58157 41792 58162 41848
rect 58218 41792 60000 41848
rect 58157 41790 60000 41792
rect 58157 41787 58223 41790
rect 59200 41760 60000 41790
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 57329 41306 57395 41309
rect 59200 41306 60000 41336
rect 57329 41304 60000 41306
rect 57329 41248 57334 41304
rect 57390 41248 60000 41304
rect 57329 41246 60000 41248
rect 57329 41243 57395 41246
rect 59200 41216 60000 41246
rect 0 41034 800 41064
rect 1393 41034 1459 41037
rect 0 41032 1459 41034
rect 0 40976 1398 41032
rect 1454 40976 1459 41032
rect 0 40974 1459 40976
rect 0 40944 800 40974
rect 1393 40971 1459 40974
rect 56501 40898 56567 40901
rect 59200 40898 60000 40928
rect 56501 40896 60000 40898
rect 56501 40840 56506 40896
rect 56562 40840 60000 40896
rect 56501 40838 60000 40840
rect 56501 40835 56567 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 59200 40808 60000 40838
rect 50288 40767 50608 40768
rect 58157 40354 58223 40357
rect 59200 40354 60000 40384
rect 58157 40352 60000 40354
rect 58157 40296 58162 40352
rect 58218 40296 60000 40352
rect 58157 40294 60000 40296
rect 58157 40291 58223 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 59200 40264 60000 40294
rect 34928 40223 35248 40224
rect 0 40082 800 40112
rect 1393 40082 1459 40085
rect 0 40080 1459 40082
rect 0 40024 1398 40080
rect 1454 40024 1459 40080
rect 0 40022 1459 40024
rect 0 39992 800 40022
rect 1393 40019 1459 40022
rect 58157 39810 58223 39813
rect 59200 39810 60000 39840
rect 58157 39808 60000 39810
rect 58157 39752 58162 39808
rect 58218 39752 60000 39808
rect 58157 39750 60000 39752
rect 58157 39747 58223 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 59200 39720 60000 39750
rect 50288 39679 50608 39680
rect 57973 39266 58039 39269
rect 59200 39266 60000 39296
rect 57973 39264 60000 39266
rect 57973 39208 57978 39264
rect 58034 39208 60000 39264
rect 57973 39206 60000 39208
rect 57973 39203 58039 39206
rect 4208 39200 4528 39201
rect 0 39130 800 39160
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 59200 39176 60000 39206
rect 34928 39135 35248 39136
rect 1393 39130 1459 39133
rect 0 39128 1459 39130
rect 0 39072 1398 39128
rect 1454 39072 1459 39128
rect 0 39070 1459 39072
rect 0 39040 800 39070
rect 1393 39067 1459 39070
rect 58157 38722 58223 38725
rect 59200 38722 60000 38752
rect 58157 38720 60000 38722
rect 58157 38664 58162 38720
rect 58218 38664 60000 38720
rect 58157 38662 60000 38664
rect 58157 38659 58223 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 59200 38632 60000 38662
rect 50288 38591 50608 38592
rect 0 38314 800 38344
rect 1393 38314 1459 38317
rect 0 38312 1459 38314
rect 0 38256 1398 38312
rect 1454 38256 1459 38312
rect 0 38254 1459 38256
rect 0 38224 800 38254
rect 1393 38251 1459 38254
rect 58157 38178 58223 38181
rect 59200 38178 60000 38208
rect 58157 38176 60000 38178
rect 58157 38120 58162 38176
rect 58218 38120 60000 38176
rect 58157 38118 60000 38120
rect 58157 38115 58223 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 59200 38088 60000 38118
rect 34928 38047 35248 38048
rect 56501 37770 56567 37773
rect 59200 37770 60000 37800
rect 56501 37768 60000 37770
rect 56501 37712 56506 37768
rect 56562 37712 60000 37768
rect 56501 37710 60000 37712
rect 56501 37707 56567 37710
rect 59200 37680 60000 37710
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 0 37362 800 37392
rect 1393 37362 1459 37365
rect 0 37360 1459 37362
rect 0 37304 1398 37360
rect 1454 37304 1459 37360
rect 0 37302 1459 37304
rect 0 37272 800 37302
rect 1393 37299 1459 37302
rect 57881 37226 57947 37229
rect 59200 37226 60000 37256
rect 57881 37224 60000 37226
rect 57881 37168 57886 37224
rect 57942 37168 60000 37224
rect 57881 37166 60000 37168
rect 57881 37163 57947 37166
rect 59200 37136 60000 37166
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 57053 36682 57119 36685
rect 59200 36682 60000 36712
rect 57053 36680 60000 36682
rect 57053 36624 57058 36680
rect 57114 36624 60000 36680
rect 57053 36622 60000 36624
rect 57053 36619 57119 36622
rect 59200 36592 60000 36622
rect 19568 36480 19888 36481
rect 0 36410 800 36440
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 1393 36410 1459 36413
rect 0 36408 1459 36410
rect 0 36352 1398 36408
rect 1454 36352 1459 36408
rect 0 36350 1459 36352
rect 0 36320 800 36350
rect 1393 36347 1459 36350
rect 56225 36138 56291 36141
rect 59200 36138 60000 36168
rect 56225 36136 60000 36138
rect 56225 36080 56230 36136
rect 56286 36080 60000 36136
rect 56225 36078 60000 36080
rect 56225 36075 56291 36078
rect 59200 36048 60000 36078
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 57881 35594 57947 35597
rect 59200 35594 60000 35624
rect 57881 35592 60000 35594
rect 57881 35536 57886 35592
rect 57942 35536 60000 35592
rect 57881 35534 60000 35536
rect 57881 35531 57947 35534
rect 59200 35504 60000 35534
rect 0 35458 800 35488
rect 1393 35458 1459 35461
rect 0 35456 1459 35458
rect 0 35400 1398 35456
rect 1454 35400 1459 35456
rect 0 35398 1459 35400
rect 0 35368 800 35398
rect 1393 35395 1459 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 58157 35050 58223 35053
rect 59200 35050 60000 35080
rect 58157 35048 60000 35050
rect 58157 34992 58162 35048
rect 58218 34992 60000 35048
rect 58157 34990 60000 34992
rect 58157 34987 58223 34990
rect 59200 34960 60000 34990
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 0 34642 800 34672
rect 1393 34642 1459 34645
rect 0 34640 1459 34642
rect 0 34584 1398 34640
rect 1454 34584 1459 34640
rect 0 34582 1459 34584
rect 0 34552 800 34582
rect 1393 34579 1459 34582
rect 55305 34642 55371 34645
rect 59200 34642 60000 34672
rect 55305 34640 60000 34642
rect 55305 34584 55310 34640
rect 55366 34584 60000 34640
rect 55305 34582 60000 34584
rect 55305 34579 55371 34582
rect 59200 34552 60000 34582
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 57881 34098 57947 34101
rect 59200 34098 60000 34128
rect 57881 34096 60000 34098
rect 57881 34040 57886 34096
rect 57942 34040 60000 34096
rect 57881 34038 60000 34040
rect 57881 34035 57947 34038
rect 59200 34008 60000 34038
rect 4208 33760 4528 33761
rect 0 33690 800 33720
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 1393 33690 1459 33693
rect 0 33688 1459 33690
rect 0 33632 1398 33688
rect 1454 33632 1459 33688
rect 0 33630 1459 33632
rect 0 33600 800 33630
rect 1393 33627 1459 33630
rect 57053 33554 57119 33557
rect 59200 33554 60000 33584
rect 57053 33552 60000 33554
rect 57053 33496 57058 33552
rect 57114 33496 60000 33552
rect 57053 33494 60000 33496
rect 57053 33491 57119 33494
rect 59200 33464 60000 33494
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 50288 33216 50608 33217
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 33151 50608 33152
rect 55213 33010 55279 33013
rect 59200 33010 60000 33040
rect 55213 33008 60000 33010
rect 55213 32952 55218 33008
rect 55274 32952 60000 33008
rect 55213 32950 60000 32952
rect 55213 32947 55279 32950
rect 59200 32920 60000 32950
rect 0 32738 800 32768
rect 1393 32738 1459 32741
rect 0 32736 1459 32738
rect 0 32680 1398 32736
rect 1454 32680 1459 32736
rect 0 32678 1459 32680
rect 0 32648 800 32678
rect 1393 32675 1459 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 58525 32466 58591 32469
rect 59200 32466 60000 32496
rect 58525 32464 60000 32466
rect 58525 32408 58530 32464
rect 58586 32408 60000 32464
rect 58525 32406 60000 32408
rect 58525 32403 58591 32406
rect 59200 32376 60000 32406
rect 23105 32330 23171 32333
rect 24025 32330 24091 32333
rect 23105 32328 24091 32330
rect 23105 32272 23110 32328
rect 23166 32272 24030 32328
rect 24086 32272 24091 32328
rect 23105 32270 24091 32272
rect 23105 32267 23171 32270
rect 24025 32267 24091 32270
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 50288 32128 50608 32129
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 32063 50608 32064
rect 56961 31922 57027 31925
rect 59200 31922 60000 31952
rect 56961 31920 60000 31922
rect 56961 31864 56966 31920
rect 57022 31864 60000 31920
rect 56961 31862 60000 31864
rect 56961 31859 57027 31862
rect 59200 31832 60000 31862
rect 0 31786 800 31816
rect 1393 31786 1459 31789
rect 0 31784 1459 31786
rect 0 31728 1398 31784
rect 1454 31728 1459 31784
rect 0 31726 1459 31728
rect 0 31696 800 31726
rect 1393 31723 1459 31726
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 56501 31514 56567 31517
rect 59200 31514 60000 31544
rect 56501 31512 60000 31514
rect 56501 31456 56506 31512
rect 56562 31456 60000 31512
rect 56501 31454 60000 31456
rect 56501 31451 56567 31454
rect 59200 31424 60000 31454
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 50288 31040 50608 31041
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 30975 50608 30976
rect 57053 30970 57119 30973
rect 59200 30970 60000 31000
rect 57053 30968 60000 30970
rect 57053 30912 57058 30968
rect 57114 30912 60000 30968
rect 57053 30910 60000 30912
rect 57053 30907 57119 30910
rect 59200 30880 60000 30910
rect 0 30834 800 30864
rect 1393 30834 1459 30837
rect 0 30832 1459 30834
rect 0 30776 1398 30832
rect 1454 30776 1459 30832
rect 0 30774 1459 30776
rect 0 30744 800 30774
rect 1393 30771 1459 30774
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 57145 30426 57211 30429
rect 59200 30426 60000 30456
rect 57145 30424 60000 30426
rect 57145 30368 57150 30424
rect 57206 30368 60000 30424
rect 57145 30366 60000 30368
rect 57145 30363 57211 30366
rect 59200 30336 60000 30366
rect 19609 30154 19675 30157
rect 22461 30154 22527 30157
rect 19609 30152 22527 30154
rect 19609 30096 19614 30152
rect 19670 30096 22466 30152
rect 22522 30096 22527 30152
rect 19609 30094 22527 30096
rect 19609 30091 19675 30094
rect 22461 30091 22527 30094
rect 29821 30154 29887 30157
rect 30465 30154 30531 30157
rect 29821 30152 30531 30154
rect 29821 30096 29826 30152
rect 29882 30096 30470 30152
rect 30526 30096 30531 30152
rect 29821 30094 30531 30096
rect 29821 30091 29887 30094
rect 30465 30091 30531 30094
rect 0 30018 800 30048
rect 1393 30018 1459 30021
rect 0 30016 1459 30018
rect 0 29960 1398 30016
rect 1454 29960 1459 30016
rect 0 29958 1459 29960
rect 0 29928 800 29958
rect 1393 29955 1459 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 50288 29952 50608 29953
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 29887 50608 29888
rect 56501 29882 56567 29885
rect 59200 29882 60000 29912
rect 56501 29880 60000 29882
rect 56501 29824 56506 29880
rect 56562 29824 60000 29880
rect 56501 29822 60000 29824
rect 56501 29819 56567 29822
rect 59200 29792 60000 29822
rect 4208 29408 4528 29409
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 0 29066 800 29096
rect 1945 29066 2011 29069
rect 0 29064 2011 29066
rect 0 29008 1950 29064
rect 2006 29008 2011 29064
rect 0 29006 2011 29008
rect 0 28976 800 29006
rect 1945 29003 2011 29006
rect 19425 29066 19491 29069
rect 23473 29066 23539 29069
rect 19425 29064 23539 29066
rect 19425 29008 19430 29064
rect 19486 29008 23478 29064
rect 23534 29008 23539 29064
rect 19425 29006 23539 29008
rect 19425 29003 19491 29006
rect 23473 29003 23539 29006
rect 31109 28930 31175 28933
rect 31569 28930 31635 28933
rect 31109 28928 31635 28930
rect 31109 28872 31114 28928
rect 31170 28872 31574 28928
rect 31630 28872 31635 28928
rect 31109 28870 31635 28872
rect 31109 28867 31175 28870
rect 31569 28867 31635 28870
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 50288 28864 50608 28865
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 28799 50608 28800
rect 9673 28794 9739 28797
rect 15837 28794 15903 28797
rect 9673 28792 15903 28794
rect 9673 28736 9678 28792
rect 9734 28736 15842 28792
rect 15898 28736 15903 28792
rect 9673 28734 15903 28736
rect 9673 28731 9739 28734
rect 15837 28731 15903 28734
rect 31293 28794 31359 28797
rect 33317 28794 33383 28797
rect 31293 28792 33383 28794
rect 31293 28736 31298 28792
rect 31354 28736 33322 28792
rect 33378 28736 33383 28792
rect 31293 28734 33383 28736
rect 31293 28731 31359 28734
rect 33317 28731 33383 28734
rect 58157 28794 58223 28797
rect 59200 28794 60000 28824
rect 58157 28792 60000 28794
rect 58157 28736 58162 28792
rect 58218 28736 60000 28792
rect 58157 28734 60000 28736
rect 58157 28731 58223 28734
rect 59200 28704 60000 28734
rect 17861 28658 17927 28661
rect 56961 28658 57027 28661
rect 17861 28656 57027 28658
rect 17861 28600 17866 28656
rect 17922 28600 56966 28656
rect 57022 28600 57027 28656
rect 17861 28598 57027 28600
rect 17861 28595 17927 28598
rect 56961 28595 57027 28598
rect 5073 28522 5139 28525
rect 8201 28522 8267 28525
rect 5073 28520 8267 28522
rect 5073 28464 5078 28520
rect 5134 28464 8206 28520
rect 8262 28464 8267 28520
rect 5073 28462 8267 28464
rect 5073 28459 5139 28462
rect 8201 28459 8267 28462
rect 18045 28522 18111 28525
rect 57881 28522 57947 28525
rect 18045 28520 57947 28522
rect 18045 28464 18050 28520
rect 18106 28464 57886 28520
rect 57942 28464 57947 28520
rect 18045 28462 57947 28464
rect 18045 28459 18111 28462
rect 57881 28459 57947 28462
rect 55581 28386 55647 28389
rect 59200 28386 60000 28416
rect 55581 28384 60000 28386
rect 55581 28328 55586 28384
rect 55642 28328 60000 28384
rect 55581 28326 60000 28328
rect 55581 28323 55647 28326
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 59200 28296 60000 28326
rect 34928 28255 35248 28256
rect 0 28114 800 28144
rect 2037 28114 2103 28117
rect 0 28112 2103 28114
rect 0 28056 2042 28112
rect 2098 28056 2103 28112
rect 0 28054 2103 28056
rect 0 28024 800 28054
rect 2037 28051 2103 28054
rect 30281 28114 30347 28117
rect 36445 28114 36511 28117
rect 30281 28112 36511 28114
rect 30281 28056 30286 28112
rect 30342 28056 36450 28112
rect 36506 28056 36511 28112
rect 30281 28054 36511 28056
rect 30281 28051 30347 28054
rect 36445 28051 36511 28054
rect 17953 27978 18019 27981
rect 18689 27978 18755 27981
rect 19149 27978 19215 27981
rect 17953 27976 19215 27978
rect 17953 27920 17958 27976
rect 18014 27920 18694 27976
rect 18750 27920 19154 27976
rect 19210 27920 19215 27976
rect 17953 27918 19215 27920
rect 17953 27915 18019 27918
rect 18689 27915 18755 27918
rect 19149 27915 19215 27918
rect 30465 27978 30531 27981
rect 34329 27978 34395 27981
rect 30465 27976 34395 27978
rect 30465 27920 30470 27976
rect 30526 27920 34334 27976
rect 34390 27920 34395 27976
rect 30465 27918 34395 27920
rect 30465 27915 30531 27918
rect 34329 27915 34395 27918
rect 14457 27842 14523 27845
rect 18137 27842 18203 27845
rect 14457 27840 18203 27842
rect 14457 27784 14462 27840
rect 14518 27784 18142 27840
rect 18198 27784 18203 27840
rect 14457 27782 18203 27784
rect 14457 27779 14523 27782
rect 18137 27779 18203 27782
rect 58157 27842 58223 27845
rect 59200 27842 60000 27872
rect 58157 27840 60000 27842
rect 58157 27784 58162 27840
rect 58218 27784 60000 27840
rect 58157 27782 60000 27784
rect 58157 27779 58223 27782
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 50288 27776 50608 27777
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 59200 27752 60000 27782
rect 50288 27711 50608 27712
rect 12249 27298 12315 27301
rect 13813 27298 13879 27301
rect 12249 27296 13879 27298
rect 12249 27240 12254 27296
rect 12310 27240 13818 27296
rect 13874 27240 13879 27296
rect 12249 27238 13879 27240
rect 12249 27235 12315 27238
rect 13813 27235 13879 27238
rect 56961 27298 57027 27301
rect 59200 27298 60000 27328
rect 56961 27296 60000 27298
rect 56961 27240 56966 27296
rect 57022 27240 60000 27296
rect 56961 27238 60000 27240
rect 56961 27235 57027 27238
rect 4208 27232 4528 27233
rect 0 27162 800 27192
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 59200 27208 60000 27238
rect 34928 27167 35248 27168
rect 1945 27162 2011 27165
rect 0 27160 2011 27162
rect 0 27104 1950 27160
rect 2006 27104 2011 27160
rect 0 27102 2011 27104
rect 0 27072 800 27102
rect 1945 27099 2011 27102
rect 17033 27162 17099 27165
rect 18781 27162 18847 27165
rect 17033 27160 18847 27162
rect 17033 27104 17038 27160
rect 17094 27104 18786 27160
rect 18842 27104 18847 27160
rect 17033 27102 18847 27104
rect 17033 27099 17099 27102
rect 18781 27099 18847 27102
rect 10133 27026 10199 27029
rect 10685 27026 10751 27029
rect 16113 27026 16179 27029
rect 10133 27024 16179 27026
rect 10133 26968 10138 27024
rect 10194 26968 10690 27024
rect 10746 26968 16118 27024
rect 16174 26968 16179 27024
rect 10133 26966 16179 26968
rect 10133 26963 10199 26966
rect 10685 26963 10751 26966
rect 16113 26963 16179 26966
rect 16573 27026 16639 27029
rect 21081 27026 21147 27029
rect 16573 27024 21147 27026
rect 16573 26968 16578 27024
rect 16634 26968 21086 27024
rect 21142 26968 21147 27024
rect 16573 26966 21147 26968
rect 16573 26963 16639 26966
rect 21081 26963 21147 26966
rect 21817 27026 21883 27029
rect 22185 27026 22251 27029
rect 21817 27024 22251 27026
rect 21817 26968 21822 27024
rect 21878 26968 22190 27024
rect 22246 26968 22251 27024
rect 21817 26966 22251 26968
rect 21817 26963 21883 26966
rect 22185 26963 22251 26966
rect 12709 26890 12775 26893
rect 16941 26890 17007 26893
rect 12709 26888 17007 26890
rect 12709 26832 12714 26888
rect 12770 26832 16946 26888
rect 17002 26832 17007 26888
rect 12709 26830 17007 26832
rect 12709 26827 12775 26830
rect 16941 26827 17007 26830
rect 17585 26890 17651 26893
rect 18413 26890 18479 26893
rect 17585 26888 18479 26890
rect 17585 26832 17590 26888
rect 17646 26832 18418 26888
rect 18474 26832 18479 26888
rect 17585 26830 18479 26832
rect 17585 26827 17651 26830
rect 18413 26827 18479 26830
rect 21357 26890 21423 26893
rect 22001 26890 22067 26893
rect 21357 26888 22067 26890
rect 21357 26832 21362 26888
rect 21418 26832 22006 26888
rect 22062 26832 22067 26888
rect 21357 26830 22067 26832
rect 21357 26827 21423 26830
rect 22001 26827 22067 26830
rect 29085 26890 29151 26893
rect 33501 26890 33567 26893
rect 29085 26888 33567 26890
rect 29085 26832 29090 26888
rect 29146 26832 33506 26888
rect 33562 26832 33567 26888
rect 29085 26830 33567 26832
rect 29085 26827 29151 26830
rect 33501 26827 33567 26830
rect 14181 26754 14247 26757
rect 17953 26754 18019 26757
rect 14181 26752 18019 26754
rect 14181 26696 14186 26752
rect 14242 26696 17958 26752
rect 18014 26696 18019 26752
rect 14181 26694 18019 26696
rect 14181 26691 14247 26694
rect 17953 26691 18019 26694
rect 55581 26754 55647 26757
rect 59200 26754 60000 26784
rect 55581 26752 60000 26754
rect 55581 26696 55586 26752
rect 55642 26696 60000 26752
rect 55581 26694 60000 26696
rect 55581 26691 55647 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 50288 26688 50608 26689
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 59200 26664 60000 26694
rect 50288 26623 50608 26624
rect 10777 26482 10843 26485
rect 11973 26482 12039 26485
rect 10777 26480 12039 26482
rect 10777 26424 10782 26480
rect 10838 26424 11978 26480
rect 12034 26424 12039 26480
rect 10777 26422 12039 26424
rect 10777 26419 10843 26422
rect 11973 26419 12039 26422
rect 16481 26482 16547 26485
rect 17861 26482 17927 26485
rect 16481 26480 17927 26482
rect 16481 26424 16486 26480
rect 16542 26424 17866 26480
rect 17922 26424 17927 26480
rect 16481 26422 17927 26424
rect 16481 26419 16547 26422
rect 17861 26419 17927 26422
rect 23657 26346 23723 26349
rect 26509 26346 26575 26349
rect 23657 26344 26575 26346
rect 23657 26288 23662 26344
rect 23718 26288 26514 26344
rect 26570 26288 26575 26344
rect 23657 26286 26575 26288
rect 23657 26283 23723 26286
rect 26509 26283 26575 26286
rect 0 26210 800 26240
rect 1393 26210 1459 26213
rect 0 26208 1459 26210
rect 0 26152 1398 26208
rect 1454 26152 1459 26208
rect 0 26150 1459 26152
rect 0 26120 800 26150
rect 1393 26147 1459 26150
rect 58341 26210 58407 26213
rect 59200 26210 60000 26240
rect 58341 26208 60000 26210
rect 58341 26152 58346 26208
rect 58402 26152 60000 26208
rect 58341 26150 60000 26152
rect 58341 26147 58407 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 59200 26120 60000 26150
rect 34928 26079 35248 26080
rect 13997 26074 14063 26077
rect 16665 26074 16731 26077
rect 13997 26072 16731 26074
rect 13997 26016 14002 26072
rect 14058 26016 16670 26072
rect 16726 26016 16731 26072
rect 13997 26014 16731 26016
rect 13997 26011 14063 26014
rect 16665 26011 16731 26014
rect 18505 26074 18571 26077
rect 21265 26074 21331 26077
rect 18505 26072 21331 26074
rect 18505 26016 18510 26072
rect 18566 26016 21270 26072
rect 21326 26016 21331 26072
rect 18505 26014 21331 26016
rect 18505 26011 18571 26014
rect 21265 26011 21331 26014
rect 18413 25938 18479 25941
rect 21357 25938 21423 25941
rect 18413 25936 21423 25938
rect 18413 25880 18418 25936
rect 18474 25880 21362 25936
rect 21418 25880 21423 25936
rect 18413 25878 21423 25880
rect 18413 25875 18479 25878
rect 21357 25875 21423 25878
rect 15101 25802 15167 25805
rect 19057 25802 19123 25805
rect 22461 25802 22527 25805
rect 15101 25800 19123 25802
rect 15101 25744 15106 25800
rect 15162 25744 19062 25800
rect 19118 25744 19123 25800
rect 15101 25742 19123 25744
rect 15101 25739 15167 25742
rect 19057 25739 19123 25742
rect 19382 25800 22527 25802
rect 19382 25744 22466 25800
rect 22522 25744 22527 25800
rect 19382 25742 22527 25744
rect 15561 25666 15627 25669
rect 18137 25666 18203 25669
rect 15561 25664 18203 25666
rect 15561 25608 15566 25664
rect 15622 25608 18142 25664
rect 18198 25608 18203 25664
rect 15561 25606 18203 25608
rect 15561 25603 15627 25606
rect 18137 25603 18203 25606
rect 18965 25666 19031 25669
rect 19382 25666 19442 25742
rect 22461 25739 22527 25742
rect 18965 25664 19442 25666
rect 18965 25608 18970 25664
rect 19026 25608 19442 25664
rect 18965 25606 19442 25608
rect 58157 25666 58223 25669
rect 59200 25666 60000 25696
rect 58157 25664 60000 25666
rect 58157 25608 58162 25664
rect 58218 25608 60000 25664
rect 58157 25606 60000 25608
rect 18965 25603 19031 25606
rect 58157 25603 58223 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 50288 25600 50608 25601
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 59200 25576 60000 25606
rect 50288 25535 50608 25536
rect 0 25394 800 25424
rect 3141 25394 3207 25397
rect 0 25392 3207 25394
rect 0 25336 3146 25392
rect 3202 25336 3207 25392
rect 0 25334 3207 25336
rect 0 25304 800 25334
rect 3141 25331 3207 25334
rect 56501 25258 56567 25261
rect 59200 25258 60000 25288
rect 56501 25256 60000 25258
rect 56501 25200 56506 25256
rect 56562 25200 60000 25256
rect 56501 25198 60000 25200
rect 56501 25195 56567 25198
rect 59200 25168 60000 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 23289 24714 23355 24717
rect 25497 24714 25563 24717
rect 26509 24714 26575 24717
rect 27797 24714 27863 24717
rect 23289 24712 27863 24714
rect 23289 24656 23294 24712
rect 23350 24656 25502 24712
rect 25558 24656 26514 24712
rect 26570 24656 27802 24712
rect 27858 24656 27863 24712
rect 23289 24654 27863 24656
rect 23289 24651 23355 24654
rect 25497 24651 25563 24654
rect 26509 24651 26575 24654
rect 27797 24651 27863 24654
rect 58157 24714 58223 24717
rect 59200 24714 60000 24744
rect 58157 24712 60000 24714
rect 58157 24656 58162 24712
rect 58218 24656 60000 24712
rect 58157 24654 60000 24656
rect 58157 24651 58223 24654
rect 59200 24624 60000 24654
rect 19568 24512 19888 24513
rect 0 24442 800 24472
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 50288 24512 50608 24513
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 24447 50608 24448
rect 1945 24442 2011 24445
rect 0 24440 2011 24442
rect 0 24384 1950 24440
rect 2006 24384 2011 24440
rect 0 24382 2011 24384
rect 0 24352 800 24382
rect 1945 24379 2011 24382
rect 10133 24442 10199 24445
rect 10777 24442 10843 24445
rect 11329 24442 11395 24445
rect 10133 24440 11395 24442
rect 10133 24384 10138 24440
rect 10194 24384 10782 24440
rect 10838 24384 11334 24440
rect 11390 24384 11395 24440
rect 10133 24382 11395 24384
rect 10133 24379 10199 24382
rect 10777 24379 10843 24382
rect 11329 24379 11395 24382
rect 7465 24306 7531 24309
rect 31477 24306 31543 24309
rect 7465 24304 31543 24306
rect 7465 24248 7470 24304
rect 7526 24248 31482 24304
rect 31538 24248 31543 24304
rect 7465 24246 31543 24248
rect 7465 24243 7531 24246
rect 31477 24243 31543 24246
rect 9581 24170 9647 24173
rect 12433 24170 12499 24173
rect 9581 24168 12499 24170
rect 9581 24112 9586 24168
rect 9642 24112 12438 24168
rect 12494 24112 12499 24168
rect 9581 24110 12499 24112
rect 9581 24107 9647 24110
rect 12433 24107 12499 24110
rect 21909 24170 21975 24173
rect 26693 24170 26759 24173
rect 21909 24168 26759 24170
rect 21909 24112 21914 24168
rect 21970 24112 26698 24168
rect 26754 24112 26759 24168
rect 21909 24110 26759 24112
rect 21909 24107 21975 24110
rect 26693 24107 26759 24110
rect 58157 24170 58223 24173
rect 59200 24170 60000 24200
rect 58157 24168 60000 24170
rect 58157 24112 58162 24168
rect 58218 24112 60000 24168
rect 58157 24110 60000 24112
rect 58157 24107 58223 24110
rect 59200 24080 60000 24110
rect 10777 24034 10843 24037
rect 17953 24034 18019 24037
rect 10777 24032 18019 24034
rect 10777 23976 10782 24032
rect 10838 23976 17958 24032
rect 18014 23976 18019 24032
rect 10777 23974 18019 23976
rect 10777 23971 10843 23974
rect 17953 23971 18019 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 11973 23762 12039 23765
rect 18689 23762 18755 23765
rect 11973 23760 18755 23762
rect 11973 23704 11978 23760
rect 12034 23704 18694 23760
rect 18750 23704 18755 23760
rect 11973 23702 18755 23704
rect 11973 23699 12039 23702
rect 18689 23699 18755 23702
rect 23381 23626 23447 23629
rect 25037 23626 25103 23629
rect 23381 23624 25103 23626
rect 23381 23568 23386 23624
rect 23442 23568 25042 23624
rect 25098 23568 25103 23624
rect 23381 23566 25103 23568
rect 23381 23563 23447 23566
rect 25037 23563 25103 23566
rect 56501 23626 56567 23629
rect 59200 23626 60000 23656
rect 56501 23624 60000 23626
rect 56501 23568 56506 23624
rect 56562 23568 60000 23624
rect 56501 23566 60000 23568
rect 56501 23563 56567 23566
rect 59200 23536 60000 23566
rect 0 23490 800 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 800 23430
rect 1577 23427 1643 23430
rect 22185 23490 22251 23493
rect 24209 23490 24275 23493
rect 22185 23488 24275 23490
rect 22185 23432 22190 23488
rect 22246 23432 24214 23488
rect 24270 23432 24275 23488
rect 22185 23430 24275 23432
rect 22185 23427 22251 23430
rect 24209 23427 24275 23430
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 50288 23424 50608 23425
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 23359 50608 23360
rect 20713 23218 20779 23221
rect 21817 23218 21883 23221
rect 23841 23218 23907 23221
rect 28809 23218 28875 23221
rect 20713 23216 22386 23218
rect 20713 23160 20718 23216
rect 20774 23160 21822 23216
rect 21878 23160 22386 23216
rect 20713 23158 22386 23160
rect 20713 23155 20779 23158
rect 21817 23155 21883 23158
rect 22326 23082 22386 23158
rect 23841 23216 28875 23218
rect 23841 23160 23846 23216
rect 23902 23160 28814 23216
rect 28870 23160 28875 23216
rect 23841 23158 28875 23160
rect 23841 23155 23907 23158
rect 28809 23155 28875 23158
rect 24301 23082 24367 23085
rect 29453 23082 29519 23085
rect 22326 23080 29519 23082
rect 22326 23024 24306 23080
rect 24362 23024 29458 23080
rect 29514 23024 29519 23080
rect 22326 23022 29519 23024
rect 24301 23019 24367 23022
rect 29453 23019 29519 23022
rect 31385 23082 31451 23085
rect 34421 23082 34487 23085
rect 31385 23080 34487 23082
rect 31385 23024 31390 23080
rect 31446 23024 34426 23080
rect 34482 23024 34487 23080
rect 31385 23022 34487 23024
rect 31385 23019 31451 23022
rect 34421 23019 34487 23022
rect 58157 23082 58223 23085
rect 59200 23082 60000 23112
rect 58157 23080 60000 23082
rect 58157 23024 58162 23080
rect 58218 23024 60000 23080
rect 58157 23022 60000 23024
rect 58157 23019 58223 23022
rect 59200 22992 60000 23022
rect 20069 22946 20135 22949
rect 26417 22946 26483 22949
rect 20069 22944 26483 22946
rect 20069 22888 20074 22944
rect 20130 22888 26422 22944
rect 26478 22888 26483 22944
rect 20069 22886 26483 22888
rect 20069 22883 20135 22886
rect 26417 22883 26483 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 19333 22674 19399 22677
rect 28625 22674 28691 22677
rect 19333 22672 28691 22674
rect 19333 22616 19338 22672
rect 19394 22616 28630 22672
rect 28686 22616 28691 22672
rect 19333 22614 28691 22616
rect 19333 22611 19399 22614
rect 28625 22611 28691 22614
rect 0 22538 800 22568
rect 1945 22538 2011 22541
rect 0 22536 2011 22538
rect 0 22480 1950 22536
rect 2006 22480 2011 22536
rect 0 22478 2011 22480
rect 0 22448 800 22478
rect 1945 22475 2011 22478
rect 19793 22538 19859 22541
rect 24025 22538 24091 22541
rect 25405 22538 25471 22541
rect 27061 22538 27127 22541
rect 27889 22538 27955 22541
rect 19793 22536 27955 22538
rect 19793 22480 19798 22536
rect 19854 22480 24030 22536
rect 24086 22480 25410 22536
rect 25466 22480 27066 22536
rect 27122 22480 27894 22536
rect 27950 22480 27955 22536
rect 19793 22478 27955 22480
rect 19793 22475 19859 22478
rect 24025 22475 24091 22478
rect 25405 22475 25471 22478
rect 27061 22475 27127 22478
rect 27889 22475 27955 22478
rect 57053 22538 57119 22541
rect 59200 22538 60000 22568
rect 57053 22536 60000 22538
rect 57053 22480 57058 22536
rect 57114 22480 60000 22536
rect 57053 22478 60000 22480
rect 57053 22475 57119 22478
rect 59200 22448 60000 22478
rect 20805 22402 20871 22405
rect 21633 22402 21699 22405
rect 20805 22400 21699 22402
rect 20805 22344 20810 22400
rect 20866 22344 21638 22400
rect 21694 22344 21699 22400
rect 20805 22342 21699 22344
rect 20805 22339 20871 22342
rect 21633 22339 21699 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 50288 22336 50608 22337
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 22271 50608 22272
rect 15561 22130 15627 22133
rect 16481 22130 16547 22133
rect 18229 22130 18295 22133
rect 15561 22128 18295 22130
rect 15561 22072 15566 22128
rect 15622 22072 16486 22128
rect 16542 22072 18234 22128
rect 18290 22072 18295 22128
rect 15561 22070 18295 22072
rect 15561 22067 15627 22070
rect 16481 22067 16547 22070
rect 18229 22067 18295 22070
rect 19333 22130 19399 22133
rect 21817 22130 21883 22133
rect 19333 22128 21883 22130
rect 19333 22072 19338 22128
rect 19394 22072 21822 22128
rect 21878 22072 21883 22128
rect 19333 22070 21883 22072
rect 19333 22067 19399 22070
rect 21817 22067 21883 22070
rect 22921 22130 22987 22133
rect 27981 22130 28047 22133
rect 28717 22130 28783 22133
rect 22921 22128 28783 22130
rect 22921 22072 22926 22128
rect 22982 22072 27986 22128
rect 28042 22072 28722 22128
rect 28778 22072 28783 22128
rect 22921 22070 28783 22072
rect 22921 22067 22987 22070
rect 27981 22067 28047 22070
rect 28717 22067 28783 22070
rect 30833 22130 30899 22133
rect 36261 22130 36327 22133
rect 30833 22128 36327 22130
rect 30833 22072 30838 22128
rect 30894 22072 36266 22128
rect 36322 22072 36327 22128
rect 30833 22070 36327 22072
rect 30833 22067 30899 22070
rect 36261 22067 36327 22070
rect 57329 22130 57395 22133
rect 59200 22130 60000 22160
rect 57329 22128 60000 22130
rect 57329 22072 57334 22128
rect 57390 22072 60000 22128
rect 57329 22070 60000 22072
rect 57329 22067 57395 22070
rect 59200 22040 60000 22070
rect 13261 21858 13327 21861
rect 18137 21858 18203 21861
rect 13261 21856 18203 21858
rect 13261 21800 13266 21856
rect 13322 21800 18142 21856
rect 18198 21800 18203 21856
rect 13261 21798 18203 21800
rect 13261 21795 13327 21798
rect 18137 21795 18203 21798
rect 23565 21858 23631 21861
rect 27337 21858 27403 21861
rect 23565 21856 27403 21858
rect 23565 21800 23570 21856
rect 23626 21800 27342 21856
rect 27398 21800 27403 21856
rect 23565 21798 27403 21800
rect 23565 21795 23631 21798
rect 27337 21795 27403 21798
rect 4208 21792 4528 21793
rect 0 21722 800 21752
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 21727 35248 21728
rect 1945 21722 2011 21725
rect 0 21720 2011 21722
rect 0 21664 1950 21720
rect 2006 21664 2011 21720
rect 0 21662 2011 21664
rect 0 21632 800 21662
rect 1945 21659 2011 21662
rect 58157 21586 58223 21589
rect 59200 21586 60000 21616
rect 58157 21584 60000 21586
rect 58157 21528 58162 21584
rect 58218 21528 60000 21584
rect 58157 21526 60000 21528
rect 58157 21523 58223 21526
rect 59200 21496 60000 21526
rect 20069 21314 20135 21317
rect 24393 21314 24459 21317
rect 24669 21314 24735 21317
rect 28809 21314 28875 21317
rect 20069 21312 20178 21314
rect 20069 21256 20074 21312
rect 20130 21256 20178 21312
rect 20069 21251 20178 21256
rect 24393 21312 28875 21314
rect 24393 21256 24398 21312
rect 24454 21256 24674 21312
rect 24730 21256 28814 21312
rect 28870 21256 28875 21312
rect 24393 21254 28875 21256
rect 24393 21251 24459 21254
rect 24669 21251 24735 21254
rect 28809 21251 28875 21254
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 17677 21042 17743 21045
rect 19241 21042 19307 21045
rect 17677 21040 19307 21042
rect 17677 20984 17682 21040
rect 17738 20984 19246 21040
rect 19302 20984 19307 21040
rect 17677 20982 19307 20984
rect 20118 21042 20178 21251
rect 50288 21248 50608 21249
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 21183 50608 21184
rect 20253 21042 20319 21045
rect 20118 21040 20319 21042
rect 20118 20984 20258 21040
rect 20314 20984 20319 21040
rect 20118 20982 20319 20984
rect 17677 20979 17743 20982
rect 19241 20979 19307 20982
rect 20253 20979 20319 20982
rect 25313 21042 25379 21045
rect 26969 21042 27035 21045
rect 25313 21040 27035 21042
rect 25313 20984 25318 21040
rect 25374 20984 26974 21040
rect 27030 20984 27035 21040
rect 25313 20982 27035 20984
rect 25313 20979 25379 20982
rect 26969 20979 27035 20982
rect 32489 21042 32555 21045
rect 34329 21042 34395 21045
rect 32489 21040 34395 21042
rect 32489 20984 32494 21040
rect 32550 20984 34334 21040
rect 34390 20984 34395 21040
rect 32489 20982 34395 20984
rect 32489 20979 32555 20982
rect 34329 20979 34395 20982
rect 58157 21042 58223 21045
rect 59200 21042 60000 21072
rect 58157 21040 60000 21042
rect 58157 20984 58162 21040
rect 58218 20984 60000 21040
rect 58157 20982 60000 20984
rect 58157 20979 58223 20982
rect 59200 20952 60000 20982
rect 19793 20906 19859 20909
rect 26693 20906 26759 20909
rect 19793 20904 26759 20906
rect 19793 20848 19798 20904
rect 19854 20848 26698 20904
rect 26754 20848 26759 20904
rect 19793 20846 26759 20848
rect 19793 20843 19859 20846
rect 26693 20843 26759 20846
rect 0 20770 800 20800
rect 1945 20770 2011 20773
rect 0 20768 2011 20770
rect 0 20712 1950 20768
rect 2006 20712 2011 20768
rect 0 20710 2011 20712
rect 0 20680 800 20710
rect 1945 20707 2011 20710
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 20529 20634 20595 20637
rect 21265 20634 21331 20637
rect 20529 20632 21331 20634
rect 20529 20576 20534 20632
rect 20590 20576 21270 20632
rect 21326 20576 21331 20632
rect 20529 20574 21331 20576
rect 20529 20571 20595 20574
rect 21265 20571 21331 20574
rect 19609 20498 19675 20501
rect 20897 20498 20963 20501
rect 19609 20496 20963 20498
rect 19609 20440 19614 20496
rect 19670 20440 20902 20496
rect 20958 20440 20963 20496
rect 19609 20438 20963 20440
rect 19609 20435 19675 20438
rect 20897 20435 20963 20438
rect 56501 20498 56567 20501
rect 59200 20498 60000 20528
rect 56501 20496 60000 20498
rect 56501 20440 56506 20496
rect 56562 20440 60000 20496
rect 56501 20438 60000 20440
rect 56501 20435 56567 20438
rect 59200 20408 60000 20438
rect 20529 20362 20595 20365
rect 23565 20362 23631 20365
rect 20529 20360 23631 20362
rect 20529 20304 20534 20360
rect 20590 20304 23570 20360
rect 23626 20304 23631 20360
rect 20529 20302 23631 20304
rect 20529 20299 20595 20302
rect 23565 20299 23631 20302
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 50288 20160 50608 20161
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 20095 50608 20096
rect 22921 19954 22987 19957
rect 25773 19954 25839 19957
rect 22921 19952 25839 19954
rect 22921 19896 22926 19952
rect 22982 19896 25778 19952
rect 25834 19896 25839 19952
rect 22921 19894 25839 19896
rect 22921 19891 22987 19894
rect 25773 19891 25839 19894
rect 58157 19954 58223 19957
rect 59200 19954 60000 19984
rect 58157 19952 60000 19954
rect 58157 19896 58162 19952
rect 58218 19896 60000 19952
rect 58157 19894 60000 19896
rect 58157 19891 58223 19894
rect 59200 19864 60000 19894
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 58157 19410 58223 19413
rect 59200 19410 60000 19440
rect 58157 19408 60000 19410
rect 58157 19352 58162 19408
rect 58218 19352 60000 19408
rect 58157 19350 60000 19352
rect 58157 19347 58223 19350
rect 59200 19320 60000 19350
rect 15101 19274 15167 19277
rect 16113 19274 16179 19277
rect 15101 19272 16179 19274
rect 15101 19216 15106 19272
rect 15162 19216 16118 19272
rect 16174 19216 16179 19272
rect 15101 19214 16179 19216
rect 15101 19211 15167 19214
rect 16113 19211 16179 19214
rect 19517 19274 19583 19277
rect 28717 19274 28783 19277
rect 19517 19272 28783 19274
rect 19517 19216 19522 19272
rect 19578 19216 28722 19272
rect 28778 19216 28783 19272
rect 19517 19214 28783 19216
rect 19517 19211 19583 19214
rect 28717 19211 28783 19214
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 50288 19072 50608 19073
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 19007 50608 19008
rect 55581 19002 55647 19005
rect 59200 19002 60000 19032
rect 55581 19000 60000 19002
rect 55581 18944 55586 19000
rect 55642 18944 60000 19000
rect 55581 18942 60000 18944
rect 55581 18939 55647 18942
rect 59200 18912 60000 18942
rect 0 18866 800 18896
rect 2037 18866 2103 18869
rect 0 18864 2103 18866
rect 0 18808 2042 18864
rect 2098 18808 2103 18864
rect 0 18806 2103 18808
rect 0 18776 800 18806
rect 2037 18803 2103 18806
rect 12249 18730 12315 18733
rect 17125 18730 17191 18733
rect 12249 18728 17191 18730
rect 12249 18672 12254 18728
rect 12310 18672 17130 18728
rect 17186 18672 17191 18728
rect 12249 18670 17191 18672
rect 12249 18667 12315 18670
rect 17125 18667 17191 18670
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 58157 18458 58223 18461
rect 59200 18458 60000 18488
rect 58157 18456 60000 18458
rect 58157 18400 58162 18456
rect 58218 18400 60000 18456
rect 58157 18398 60000 18400
rect 58157 18395 58223 18398
rect 59200 18368 60000 18398
rect 12433 18186 12499 18189
rect 18045 18186 18111 18189
rect 12433 18184 18111 18186
rect 12433 18128 12438 18184
rect 12494 18128 18050 18184
rect 18106 18128 18111 18184
rect 12433 18126 18111 18128
rect 12433 18123 12499 18126
rect 18045 18123 18111 18126
rect 19568 17984 19888 17985
rect 0 17914 800 17944
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 50288 17984 50608 17985
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 17919 50608 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 800 17854
rect 1945 17851 2011 17854
rect 58157 17914 58223 17917
rect 59200 17914 60000 17944
rect 58157 17912 60000 17914
rect 58157 17856 58162 17912
rect 58218 17856 60000 17912
rect 58157 17854 60000 17856
rect 58157 17851 58223 17854
rect 59200 17824 60000 17854
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 56225 17370 56291 17373
rect 59200 17370 60000 17400
rect 56225 17368 60000 17370
rect 56225 17312 56230 17368
rect 56286 17312 60000 17368
rect 56225 17310 60000 17312
rect 56225 17307 56291 17310
rect 59200 17280 60000 17310
rect 0 17098 800 17128
rect 2037 17098 2103 17101
rect 0 17096 2103 17098
rect 0 17040 2042 17096
rect 2098 17040 2103 17096
rect 0 17038 2103 17040
rect 0 17008 800 17038
rect 2037 17035 2103 17038
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 50288 16896 50608 16897
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 16831 50608 16832
rect 58157 16826 58223 16829
rect 59200 16826 60000 16856
rect 58157 16824 60000 16826
rect 58157 16768 58162 16824
rect 58218 16768 60000 16824
rect 58157 16766 60000 16768
rect 58157 16763 58223 16766
rect 59200 16736 60000 16766
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 16287 35248 16288
rect 58249 16282 58315 16285
rect 59200 16282 60000 16312
rect 58249 16280 60000 16282
rect 58249 16224 58254 16280
rect 58310 16224 60000 16280
rect 58249 16222 60000 16224
rect 58249 16219 58315 16222
rect 59200 16192 60000 16222
rect 0 16146 800 16176
rect 2037 16146 2103 16149
rect 0 16144 2103 16146
rect 0 16088 2042 16144
rect 2098 16088 2103 16144
rect 0 16086 2103 16088
rect 0 16056 800 16086
rect 2037 16083 2103 16086
rect 55581 15874 55647 15877
rect 59200 15874 60000 15904
rect 55581 15872 60000 15874
rect 55581 15816 55586 15872
rect 55642 15816 60000 15872
rect 55581 15814 60000 15816
rect 55581 15811 55647 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 50288 15808 50608 15809
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 59200 15784 60000 15814
rect 50288 15743 50608 15744
rect 58065 15330 58131 15333
rect 59200 15330 60000 15360
rect 58065 15328 60000 15330
rect 58065 15272 58070 15328
rect 58126 15272 60000 15328
rect 58065 15270 60000 15272
rect 58065 15267 58131 15270
rect 4208 15264 4528 15265
rect 0 15194 800 15224
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 59200 15240 60000 15270
rect 34928 15199 35248 15200
rect 1945 15194 2011 15197
rect 0 15192 2011 15194
rect 0 15136 1950 15192
rect 2006 15136 2011 15192
rect 0 15134 2011 15136
rect 0 15104 800 15134
rect 1945 15131 2011 15134
rect 56961 14786 57027 14789
rect 59200 14786 60000 14816
rect 56961 14784 60000 14786
rect 56961 14728 56966 14784
rect 57022 14728 60000 14784
rect 56961 14726 60000 14728
rect 56961 14723 57027 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 50288 14720 50608 14721
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 59200 14696 60000 14726
rect 50288 14655 50608 14656
rect 0 14242 800 14272
rect 1945 14242 2011 14245
rect 0 14240 2011 14242
rect 0 14184 1950 14240
rect 2006 14184 2011 14240
rect 0 14182 2011 14184
rect 0 14152 800 14182
rect 1945 14179 2011 14182
rect 55581 14242 55647 14245
rect 59200 14242 60000 14272
rect 55581 14240 60000 14242
rect 55581 14184 55586 14240
rect 55642 14184 60000 14240
rect 55581 14182 60000 14184
rect 55581 14179 55647 14182
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 59200 14152 60000 14182
rect 34928 14111 35248 14112
rect 58065 13698 58131 13701
rect 59200 13698 60000 13728
rect 58065 13696 60000 13698
rect 58065 13640 58070 13696
rect 58126 13640 60000 13696
rect 58065 13638 60000 13640
rect 58065 13635 58131 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 50288 13632 50608 13633
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 59200 13608 60000 13638
rect 50288 13567 50608 13568
rect 0 13290 800 13320
rect 2037 13290 2103 13293
rect 0 13288 2103 13290
rect 0 13232 2042 13288
rect 2098 13232 2103 13288
rect 0 13230 2103 13232
rect 0 13200 800 13230
rect 2037 13227 2103 13230
rect 57329 13154 57395 13157
rect 59200 13154 60000 13184
rect 57329 13152 60000 13154
rect 57329 13096 57334 13152
rect 57390 13096 60000 13152
rect 57329 13094 60000 13096
rect 57329 13091 57395 13094
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 59200 13064 60000 13094
rect 34928 13023 35248 13024
rect 55397 12746 55463 12749
rect 59200 12746 60000 12776
rect 55397 12744 60000 12746
rect 55397 12688 55402 12744
rect 55458 12688 60000 12744
rect 55397 12686 60000 12688
rect 55397 12683 55463 12686
rect 59200 12656 60000 12686
rect 19568 12544 19888 12545
rect 0 12474 800 12504
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 50288 12544 50608 12545
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 12479 50608 12480
rect 1945 12474 2011 12477
rect 0 12472 2011 12474
rect 0 12416 1950 12472
rect 2006 12416 2011 12472
rect 0 12414 2011 12416
rect 0 12384 800 12414
rect 1945 12411 2011 12414
rect 57881 12202 57947 12205
rect 59200 12202 60000 12232
rect 57881 12200 60000 12202
rect 57881 12144 57886 12200
rect 57942 12144 60000 12200
rect 57881 12142 60000 12144
rect 57881 12139 57947 12142
rect 59200 12112 60000 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 56501 11658 56567 11661
rect 59200 11658 60000 11688
rect 56501 11656 60000 11658
rect 56501 11600 56506 11656
rect 56562 11600 60000 11656
rect 56501 11598 60000 11600
rect 56501 11595 56567 11598
rect 59200 11568 60000 11598
rect 0 11522 800 11552
rect 1945 11522 2011 11525
rect 0 11520 2011 11522
rect 0 11464 1950 11520
rect 2006 11464 2011 11520
rect 0 11462 2011 11464
rect 0 11432 800 11462
rect 1945 11459 2011 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 50288 11456 50608 11457
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 11391 50608 11392
rect 55581 11114 55647 11117
rect 59200 11114 60000 11144
rect 55581 11112 60000 11114
rect 55581 11056 55586 11112
rect 55642 11056 60000 11112
rect 55581 11054 60000 11056
rect 55581 11051 55647 11054
rect 59200 11024 60000 11054
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 10847 35248 10848
rect 0 10570 800 10600
rect 2037 10570 2103 10573
rect 0 10568 2103 10570
rect 0 10512 2042 10568
rect 2098 10512 2103 10568
rect 0 10510 2103 10512
rect 0 10480 800 10510
rect 2037 10507 2103 10510
rect 57881 10570 57947 10573
rect 59200 10570 60000 10600
rect 57881 10568 60000 10570
rect 57881 10512 57886 10568
rect 57942 10512 60000 10568
rect 57881 10510 60000 10512
rect 57881 10507 57947 10510
rect 59200 10480 60000 10510
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 50288 10368 50608 10369
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 10303 50608 10304
rect 58157 10026 58223 10029
rect 59200 10026 60000 10056
rect 58157 10024 60000 10026
rect 58157 9968 58162 10024
rect 58218 9968 60000 10024
rect 58157 9966 60000 9968
rect 58157 9963 58223 9966
rect 59200 9936 60000 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 0 9618 800 9648
rect 2037 9618 2103 9621
rect 0 9616 2103 9618
rect 0 9560 2042 9616
rect 2098 9560 2103 9616
rect 0 9558 2103 9560
rect 0 9528 800 9558
rect 2037 9555 2103 9558
rect 55581 9618 55647 9621
rect 59200 9618 60000 9648
rect 55581 9616 60000 9618
rect 55581 9560 55586 9616
rect 55642 9560 60000 9616
rect 55581 9558 60000 9560
rect 55581 9555 55647 9558
rect 59200 9528 60000 9558
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 50288 9280 50608 9281
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 9215 50608 9216
rect 58157 9074 58223 9077
rect 59200 9074 60000 9104
rect 58157 9072 60000 9074
rect 58157 9016 58162 9072
rect 58218 9016 60000 9072
rect 58157 9014 60000 9016
rect 58157 9011 58223 9014
rect 59200 8984 60000 9014
rect 0 8802 800 8832
rect 1945 8802 2011 8805
rect 0 8800 2011 8802
rect 0 8744 1950 8800
rect 2006 8744 2011 8800
rect 0 8742 2011 8744
rect 0 8712 800 8742
rect 1945 8739 2011 8742
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 57421 8530 57487 8533
rect 59200 8530 60000 8560
rect 57421 8528 60000 8530
rect 57421 8472 57426 8528
rect 57482 8472 60000 8528
rect 57421 8470 60000 8472
rect 57421 8467 57487 8470
rect 59200 8440 60000 8470
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 50288 8192 50608 8193
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 8127 50608 8128
rect 55673 7986 55739 7989
rect 59200 7986 60000 8016
rect 55673 7984 60000 7986
rect 55673 7928 55678 7984
rect 55734 7928 60000 7984
rect 55673 7926 60000 7928
rect 55673 7923 55739 7926
rect 59200 7896 60000 7926
rect 0 7850 800 7880
rect 2037 7850 2103 7853
rect 0 7848 2103 7850
rect 0 7792 2042 7848
rect 2098 7792 2103 7848
rect 0 7790 2103 7792
rect 0 7760 800 7790
rect 2037 7787 2103 7790
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 58157 7442 58223 7445
rect 59200 7442 60000 7472
rect 58157 7440 60000 7442
rect 58157 7384 58162 7440
rect 58218 7384 60000 7440
rect 58157 7382 60000 7384
rect 58157 7379 58223 7382
rect 59200 7352 60000 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 50288 7104 50608 7105
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 7039 50608 7040
rect 0 6898 800 6928
rect 2037 6898 2103 6901
rect 0 6896 2103 6898
rect 0 6840 2042 6896
rect 2098 6840 2103 6896
rect 0 6838 2103 6840
rect 0 6808 800 6838
rect 2037 6835 2103 6838
rect 56409 6898 56475 6901
rect 59200 6898 60000 6928
rect 56409 6896 60000 6898
rect 56409 6840 56414 6896
rect 56470 6840 60000 6896
rect 56409 6838 60000 6840
rect 56409 6835 56475 6838
rect 59200 6808 60000 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 55489 6490 55555 6493
rect 59200 6490 60000 6520
rect 55489 6488 60000 6490
rect 55489 6432 55494 6488
rect 55550 6432 60000 6488
rect 55489 6430 60000 6432
rect 55489 6427 55555 6430
rect 59200 6400 60000 6430
rect 55489 6354 55555 6357
rect 56593 6354 56659 6357
rect 55489 6352 56659 6354
rect 55489 6296 55494 6352
rect 55550 6296 56598 6352
rect 56654 6296 56659 6352
rect 55489 6294 56659 6296
rect 55489 6291 55555 6294
rect 56593 6291 56659 6294
rect 19568 6016 19888 6017
rect 0 5946 800 5976
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 50288 6016 50608 6017
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 5951 50608 5952
rect 1945 5946 2011 5949
rect 0 5944 2011 5946
rect 0 5888 1950 5944
rect 2006 5888 2011 5944
rect 0 5886 2011 5888
rect 0 5856 800 5886
rect 1945 5883 2011 5886
rect 58157 5946 58223 5949
rect 59200 5946 60000 5976
rect 58157 5944 60000 5946
rect 58157 5888 58162 5944
rect 58218 5888 60000 5944
rect 58157 5886 60000 5888
rect 58157 5883 58223 5886
rect 59200 5856 60000 5886
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 57881 5402 57947 5405
rect 59200 5402 60000 5432
rect 57881 5400 60000 5402
rect 57881 5344 57886 5400
rect 57942 5344 60000 5400
rect 57881 5342 60000 5344
rect 57881 5339 57947 5342
rect 59200 5312 60000 5342
rect 0 4994 800 5024
rect 1945 4994 2011 4997
rect 0 4992 2011 4994
rect 0 4936 1950 4992
rect 2006 4936 2011 4992
rect 0 4934 2011 4936
rect 0 4904 800 4934
rect 1945 4931 2011 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 50288 4928 50608 4929
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 4863 50608 4864
rect 55213 4858 55279 4861
rect 59200 4858 60000 4888
rect 55213 4856 60000 4858
rect 55213 4800 55218 4856
rect 55274 4800 60000 4856
rect 55213 4798 60000 4800
rect 55213 4795 55279 4798
rect 59200 4768 60000 4798
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 56961 4314 57027 4317
rect 59200 4314 60000 4344
rect 56961 4312 60000 4314
rect 56961 4256 56966 4312
rect 57022 4256 60000 4312
rect 56961 4254 60000 4256
rect 56961 4251 57027 4254
rect 59200 4224 60000 4254
rect 0 4178 800 4208
rect 2037 4178 2103 4181
rect 0 4176 2103 4178
rect 0 4120 2042 4176
rect 2098 4120 2103 4176
rect 0 4118 2103 4120
rect 0 4088 800 4118
rect 2037 4115 2103 4118
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 50288 3840 50608 3841
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 3775 50608 3776
rect 57053 3770 57119 3773
rect 59200 3770 60000 3800
rect 57053 3768 60000 3770
rect 57053 3712 57058 3768
rect 57114 3712 60000 3768
rect 57053 3710 60000 3712
rect 57053 3707 57119 3710
rect 59200 3680 60000 3710
rect 55121 3362 55187 3365
rect 59200 3362 60000 3392
rect 55121 3360 60000 3362
rect 55121 3304 55126 3360
rect 55182 3304 60000 3360
rect 55121 3302 60000 3304
rect 55121 3299 55187 3302
rect 4208 3296 4528 3297
rect 0 3226 800 3256
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 59200 3272 60000 3302
rect 34928 3231 35248 3232
rect 3049 3226 3115 3229
rect 0 3224 3115 3226
rect 0 3168 3054 3224
rect 3110 3168 3115 3224
rect 0 3166 3115 3168
rect 0 3136 800 3166
rect 3049 3163 3115 3166
rect 58157 2818 58223 2821
rect 59200 2818 60000 2848
rect 58157 2816 60000 2818
rect 58157 2760 58162 2816
rect 58218 2760 60000 2816
rect 58157 2758 60000 2760
rect 58157 2755 58223 2758
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 50288 2752 50608 2753
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 59200 2728 60000 2758
rect 50288 2687 50608 2688
rect 0 2274 800 2304
rect 1945 2274 2011 2277
rect 0 2272 2011 2274
rect 0 2216 1950 2272
rect 2006 2216 2011 2272
rect 0 2214 2011 2216
rect 0 2184 800 2214
rect 1945 2211 2011 2214
rect 55949 2274 56015 2277
rect 59200 2274 60000 2304
rect 55949 2272 60000 2274
rect 55949 2216 55954 2272
rect 56010 2216 60000 2272
rect 55949 2214 60000 2216
rect 55949 2211 56015 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 59200 2184 60000 2214
rect 34928 2143 35248 2144
rect 56501 1730 56567 1733
rect 59200 1730 60000 1760
rect 56501 1728 60000 1730
rect 56501 1672 56506 1728
rect 56562 1672 60000 1728
rect 56501 1670 60000 1672
rect 56501 1667 56567 1670
rect 59200 1640 60000 1670
rect 0 1322 800 1352
rect 2773 1322 2839 1325
rect 0 1320 2839 1322
rect 0 1264 2778 1320
rect 2834 1264 2839 1320
rect 0 1262 2839 1264
rect 0 1232 800 1262
rect 2773 1259 2839 1262
rect 57881 1186 57947 1189
rect 59200 1186 60000 1216
rect 57881 1184 60000 1186
rect 57881 1128 57886 1184
rect 57942 1128 60000 1184
rect 57881 1126 60000 1128
rect 57881 1123 57947 1126
rect 59200 1096 60000 1126
rect 55581 642 55647 645
rect 59200 642 60000 672
rect 55581 640 60000 642
rect 55581 584 55586 640
rect 55642 584 60000 640
rect 55581 582 60000 584
rect 55581 579 55647 582
rect 59200 552 60000 582
rect 0 506 800 536
rect 2865 506 2931 509
rect 0 504 2931 506
rect 0 448 2870 504
rect 2926 448 2931 504
rect 0 446 2931 448
rect 0 416 800 446
rect 2865 443 2931 446
rect 56317 234 56383 237
rect 59200 234 60000 264
rect 56317 232 60000 234
rect 56317 176 56322 232
rect 56378 176 60000 232
rect 56317 174 60000 176
rect 56317 171 56383 174
rect 59200 144 60000 174
<< via3 >>
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 50296 57148 50360 57152
rect 50296 57092 50300 57148
rect 50300 57092 50356 57148
rect 50356 57092 50360 57148
rect 50296 57088 50360 57092
rect 50376 57148 50440 57152
rect 50376 57092 50380 57148
rect 50380 57092 50436 57148
rect 50436 57092 50440 57148
rect 50376 57088 50440 57092
rect 50456 57148 50520 57152
rect 50456 57092 50460 57148
rect 50460 57092 50516 57148
rect 50516 57092 50520 57148
rect 50456 57088 50520 57092
rect 50536 57148 50600 57152
rect 50536 57092 50540 57148
rect 50540 57092 50596 57148
rect 50596 57092 50600 57148
rect 50536 57088 50600 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 50296 56060 50360 56064
rect 50296 56004 50300 56060
rect 50300 56004 50356 56060
rect 50356 56004 50360 56060
rect 50296 56000 50360 56004
rect 50376 56060 50440 56064
rect 50376 56004 50380 56060
rect 50380 56004 50436 56060
rect 50436 56004 50440 56060
rect 50376 56000 50440 56004
rect 50456 56060 50520 56064
rect 50456 56004 50460 56060
rect 50460 56004 50516 56060
rect 50516 56004 50520 56060
rect 50456 56000 50520 56004
rect 50536 56060 50600 56064
rect 50536 56004 50540 56060
rect 50540 56004 50596 56060
rect 50596 56004 50600 56060
rect 50536 56000 50600 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 50296 54972 50360 54976
rect 50296 54916 50300 54972
rect 50300 54916 50356 54972
rect 50356 54916 50360 54972
rect 50296 54912 50360 54916
rect 50376 54972 50440 54976
rect 50376 54916 50380 54972
rect 50380 54916 50436 54972
rect 50436 54916 50440 54972
rect 50376 54912 50440 54916
rect 50456 54972 50520 54976
rect 50456 54916 50460 54972
rect 50460 54916 50516 54972
rect 50516 54916 50520 54972
rect 50456 54912 50520 54916
rect 50536 54972 50600 54976
rect 50536 54916 50540 54972
rect 50540 54916 50596 54972
rect 50596 54916 50600 54972
rect 50536 54912 50600 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 50296 53884 50360 53888
rect 50296 53828 50300 53884
rect 50300 53828 50356 53884
rect 50356 53828 50360 53884
rect 50296 53824 50360 53828
rect 50376 53884 50440 53888
rect 50376 53828 50380 53884
rect 50380 53828 50436 53884
rect 50436 53828 50440 53884
rect 50376 53824 50440 53828
rect 50456 53884 50520 53888
rect 50456 53828 50460 53884
rect 50460 53828 50516 53884
rect 50516 53828 50520 53884
rect 50456 53824 50520 53828
rect 50536 53884 50600 53888
rect 50536 53828 50540 53884
rect 50540 53828 50596 53884
rect 50596 53828 50600 53884
rect 50536 53824 50600 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 50296 52796 50360 52800
rect 50296 52740 50300 52796
rect 50300 52740 50356 52796
rect 50356 52740 50360 52796
rect 50296 52736 50360 52740
rect 50376 52796 50440 52800
rect 50376 52740 50380 52796
rect 50380 52740 50436 52796
rect 50436 52740 50440 52796
rect 50376 52736 50440 52740
rect 50456 52796 50520 52800
rect 50456 52740 50460 52796
rect 50460 52740 50516 52796
rect 50516 52740 50520 52796
rect 50456 52736 50520 52740
rect 50536 52796 50600 52800
rect 50536 52740 50540 52796
rect 50540 52740 50596 52796
rect 50596 52740 50600 52796
rect 50536 52736 50600 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 50296 51708 50360 51712
rect 50296 51652 50300 51708
rect 50300 51652 50356 51708
rect 50356 51652 50360 51708
rect 50296 51648 50360 51652
rect 50376 51708 50440 51712
rect 50376 51652 50380 51708
rect 50380 51652 50436 51708
rect 50436 51652 50440 51708
rect 50376 51648 50440 51652
rect 50456 51708 50520 51712
rect 50456 51652 50460 51708
rect 50460 51652 50516 51708
rect 50516 51652 50520 51708
rect 50456 51648 50520 51652
rect 50536 51708 50600 51712
rect 50536 51652 50540 51708
rect 50540 51652 50596 51708
rect 50596 51652 50600 51708
rect 50536 51648 50600 51652
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 50296 50620 50360 50624
rect 50296 50564 50300 50620
rect 50300 50564 50356 50620
rect 50356 50564 50360 50620
rect 50296 50560 50360 50564
rect 50376 50620 50440 50624
rect 50376 50564 50380 50620
rect 50380 50564 50436 50620
rect 50436 50564 50440 50620
rect 50376 50560 50440 50564
rect 50456 50620 50520 50624
rect 50456 50564 50460 50620
rect 50460 50564 50516 50620
rect 50516 50564 50520 50620
rect 50456 50560 50520 50564
rect 50536 50620 50600 50624
rect 50536 50564 50540 50620
rect 50540 50564 50596 50620
rect 50596 50564 50600 50620
rect 50536 50560 50600 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 50296 49532 50360 49536
rect 50296 49476 50300 49532
rect 50300 49476 50356 49532
rect 50356 49476 50360 49532
rect 50296 49472 50360 49476
rect 50376 49532 50440 49536
rect 50376 49476 50380 49532
rect 50380 49476 50436 49532
rect 50436 49476 50440 49532
rect 50376 49472 50440 49476
rect 50456 49532 50520 49536
rect 50456 49476 50460 49532
rect 50460 49476 50516 49532
rect 50516 49476 50520 49532
rect 50456 49472 50520 49476
rect 50536 49532 50600 49536
rect 50536 49476 50540 49532
rect 50540 49476 50596 49532
rect 50596 49476 50600 49532
rect 50536 49472 50600 49476
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 50296 48444 50360 48448
rect 50296 48388 50300 48444
rect 50300 48388 50356 48444
rect 50356 48388 50360 48444
rect 50296 48384 50360 48388
rect 50376 48444 50440 48448
rect 50376 48388 50380 48444
rect 50380 48388 50436 48444
rect 50436 48388 50440 48444
rect 50376 48384 50440 48388
rect 50456 48444 50520 48448
rect 50456 48388 50460 48444
rect 50460 48388 50516 48444
rect 50516 48388 50520 48444
rect 50456 48384 50520 48388
rect 50536 48444 50600 48448
rect 50536 48388 50540 48444
rect 50540 48388 50596 48444
rect 50596 48388 50600 48444
rect 50536 48384 50600 48388
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 50296 47356 50360 47360
rect 50296 47300 50300 47356
rect 50300 47300 50356 47356
rect 50356 47300 50360 47356
rect 50296 47296 50360 47300
rect 50376 47356 50440 47360
rect 50376 47300 50380 47356
rect 50380 47300 50436 47356
rect 50436 47300 50440 47356
rect 50376 47296 50440 47300
rect 50456 47356 50520 47360
rect 50456 47300 50460 47356
rect 50460 47300 50516 47356
rect 50516 47300 50520 47356
rect 50456 47296 50520 47300
rect 50536 47356 50600 47360
rect 50536 47300 50540 47356
rect 50540 47300 50596 47356
rect 50596 47300 50600 47356
rect 50536 47296 50600 47300
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 50296 46268 50360 46272
rect 50296 46212 50300 46268
rect 50300 46212 50356 46268
rect 50356 46212 50360 46268
rect 50296 46208 50360 46212
rect 50376 46268 50440 46272
rect 50376 46212 50380 46268
rect 50380 46212 50436 46268
rect 50436 46212 50440 46268
rect 50376 46208 50440 46212
rect 50456 46268 50520 46272
rect 50456 46212 50460 46268
rect 50460 46212 50516 46268
rect 50516 46212 50520 46268
rect 50456 46208 50520 46212
rect 50536 46268 50600 46272
rect 50536 46212 50540 46268
rect 50540 46212 50596 46268
rect 50596 46212 50600 46268
rect 50536 46208 50600 46212
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 50296 45180 50360 45184
rect 50296 45124 50300 45180
rect 50300 45124 50356 45180
rect 50356 45124 50360 45180
rect 50296 45120 50360 45124
rect 50376 45180 50440 45184
rect 50376 45124 50380 45180
rect 50380 45124 50436 45180
rect 50436 45124 50440 45180
rect 50376 45120 50440 45124
rect 50456 45180 50520 45184
rect 50456 45124 50460 45180
rect 50460 45124 50516 45180
rect 50516 45124 50520 45180
rect 50456 45120 50520 45124
rect 50536 45180 50600 45184
rect 50536 45124 50540 45180
rect 50540 45124 50596 45180
rect 50596 45124 50600 45180
rect 50536 45120 50600 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 50296 33212 50360 33216
rect 50296 33156 50300 33212
rect 50300 33156 50356 33212
rect 50356 33156 50360 33212
rect 50296 33152 50360 33156
rect 50376 33212 50440 33216
rect 50376 33156 50380 33212
rect 50380 33156 50436 33212
rect 50436 33156 50440 33212
rect 50376 33152 50440 33156
rect 50456 33212 50520 33216
rect 50456 33156 50460 33212
rect 50460 33156 50516 33212
rect 50516 33156 50520 33212
rect 50456 33152 50520 33156
rect 50536 33212 50600 33216
rect 50536 33156 50540 33212
rect 50540 33156 50596 33212
rect 50596 33156 50600 33212
rect 50536 33152 50600 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 50296 32124 50360 32128
rect 50296 32068 50300 32124
rect 50300 32068 50356 32124
rect 50356 32068 50360 32124
rect 50296 32064 50360 32068
rect 50376 32124 50440 32128
rect 50376 32068 50380 32124
rect 50380 32068 50436 32124
rect 50436 32068 50440 32124
rect 50376 32064 50440 32068
rect 50456 32124 50520 32128
rect 50456 32068 50460 32124
rect 50460 32068 50516 32124
rect 50516 32068 50520 32124
rect 50456 32064 50520 32068
rect 50536 32124 50600 32128
rect 50536 32068 50540 32124
rect 50540 32068 50596 32124
rect 50596 32068 50600 32124
rect 50536 32064 50600 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 50296 31036 50360 31040
rect 50296 30980 50300 31036
rect 50300 30980 50356 31036
rect 50356 30980 50360 31036
rect 50296 30976 50360 30980
rect 50376 31036 50440 31040
rect 50376 30980 50380 31036
rect 50380 30980 50436 31036
rect 50436 30980 50440 31036
rect 50376 30976 50440 30980
rect 50456 31036 50520 31040
rect 50456 30980 50460 31036
rect 50460 30980 50516 31036
rect 50516 30980 50520 31036
rect 50456 30976 50520 30980
rect 50536 31036 50600 31040
rect 50536 30980 50540 31036
rect 50540 30980 50596 31036
rect 50596 30980 50600 31036
rect 50536 30976 50600 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 50296 29948 50360 29952
rect 50296 29892 50300 29948
rect 50300 29892 50356 29948
rect 50356 29892 50360 29948
rect 50296 29888 50360 29892
rect 50376 29948 50440 29952
rect 50376 29892 50380 29948
rect 50380 29892 50436 29948
rect 50436 29892 50440 29948
rect 50376 29888 50440 29892
rect 50456 29948 50520 29952
rect 50456 29892 50460 29948
rect 50460 29892 50516 29948
rect 50516 29892 50520 29948
rect 50456 29888 50520 29892
rect 50536 29948 50600 29952
rect 50536 29892 50540 29948
rect 50540 29892 50596 29948
rect 50596 29892 50600 29948
rect 50536 29888 50600 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 50296 28860 50360 28864
rect 50296 28804 50300 28860
rect 50300 28804 50356 28860
rect 50356 28804 50360 28860
rect 50296 28800 50360 28804
rect 50376 28860 50440 28864
rect 50376 28804 50380 28860
rect 50380 28804 50436 28860
rect 50436 28804 50440 28860
rect 50376 28800 50440 28804
rect 50456 28860 50520 28864
rect 50456 28804 50460 28860
rect 50460 28804 50516 28860
rect 50516 28804 50520 28860
rect 50456 28800 50520 28804
rect 50536 28860 50600 28864
rect 50536 28804 50540 28860
rect 50540 28804 50596 28860
rect 50596 28804 50600 28860
rect 50536 28800 50600 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 50296 27772 50360 27776
rect 50296 27716 50300 27772
rect 50300 27716 50356 27772
rect 50356 27716 50360 27772
rect 50296 27712 50360 27716
rect 50376 27772 50440 27776
rect 50376 27716 50380 27772
rect 50380 27716 50436 27772
rect 50436 27716 50440 27772
rect 50376 27712 50440 27716
rect 50456 27772 50520 27776
rect 50456 27716 50460 27772
rect 50460 27716 50516 27772
rect 50516 27716 50520 27772
rect 50456 27712 50520 27716
rect 50536 27772 50600 27776
rect 50536 27716 50540 27772
rect 50540 27716 50596 27772
rect 50596 27716 50600 27772
rect 50536 27712 50600 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 50296 26684 50360 26688
rect 50296 26628 50300 26684
rect 50300 26628 50356 26684
rect 50356 26628 50360 26684
rect 50296 26624 50360 26628
rect 50376 26684 50440 26688
rect 50376 26628 50380 26684
rect 50380 26628 50436 26684
rect 50436 26628 50440 26684
rect 50376 26624 50440 26628
rect 50456 26684 50520 26688
rect 50456 26628 50460 26684
rect 50460 26628 50516 26684
rect 50516 26628 50520 26684
rect 50456 26624 50520 26628
rect 50536 26684 50600 26688
rect 50536 26628 50540 26684
rect 50540 26628 50596 26684
rect 50596 26628 50600 26684
rect 50536 26624 50600 26628
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 50296 25596 50360 25600
rect 50296 25540 50300 25596
rect 50300 25540 50356 25596
rect 50356 25540 50360 25596
rect 50296 25536 50360 25540
rect 50376 25596 50440 25600
rect 50376 25540 50380 25596
rect 50380 25540 50436 25596
rect 50436 25540 50440 25596
rect 50376 25536 50440 25540
rect 50456 25596 50520 25600
rect 50456 25540 50460 25596
rect 50460 25540 50516 25596
rect 50516 25540 50520 25596
rect 50456 25536 50520 25540
rect 50536 25596 50600 25600
rect 50536 25540 50540 25596
rect 50540 25540 50596 25596
rect 50596 25540 50600 25596
rect 50536 25536 50600 25540
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 50296 24508 50360 24512
rect 50296 24452 50300 24508
rect 50300 24452 50356 24508
rect 50356 24452 50360 24508
rect 50296 24448 50360 24452
rect 50376 24508 50440 24512
rect 50376 24452 50380 24508
rect 50380 24452 50436 24508
rect 50436 24452 50440 24508
rect 50376 24448 50440 24452
rect 50456 24508 50520 24512
rect 50456 24452 50460 24508
rect 50460 24452 50516 24508
rect 50516 24452 50520 24508
rect 50456 24448 50520 24452
rect 50536 24508 50600 24512
rect 50536 24452 50540 24508
rect 50540 24452 50596 24508
rect 50596 24452 50600 24508
rect 50536 24448 50600 24452
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 50296 23420 50360 23424
rect 50296 23364 50300 23420
rect 50300 23364 50356 23420
rect 50356 23364 50360 23420
rect 50296 23360 50360 23364
rect 50376 23420 50440 23424
rect 50376 23364 50380 23420
rect 50380 23364 50436 23420
rect 50436 23364 50440 23420
rect 50376 23360 50440 23364
rect 50456 23420 50520 23424
rect 50456 23364 50460 23420
rect 50460 23364 50516 23420
rect 50516 23364 50520 23420
rect 50456 23360 50520 23364
rect 50536 23420 50600 23424
rect 50536 23364 50540 23420
rect 50540 23364 50596 23420
rect 50596 23364 50600 23420
rect 50536 23360 50600 23364
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 50296 22332 50360 22336
rect 50296 22276 50300 22332
rect 50300 22276 50356 22332
rect 50356 22276 50360 22332
rect 50296 22272 50360 22276
rect 50376 22332 50440 22336
rect 50376 22276 50380 22332
rect 50380 22276 50436 22332
rect 50436 22276 50440 22332
rect 50376 22272 50440 22276
rect 50456 22332 50520 22336
rect 50456 22276 50460 22332
rect 50460 22276 50516 22332
rect 50516 22276 50520 22332
rect 50456 22272 50520 22276
rect 50536 22332 50600 22336
rect 50536 22276 50540 22332
rect 50540 22276 50596 22332
rect 50596 22276 50600 22332
rect 50536 22272 50600 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 50296 21244 50360 21248
rect 50296 21188 50300 21244
rect 50300 21188 50356 21244
rect 50356 21188 50360 21244
rect 50296 21184 50360 21188
rect 50376 21244 50440 21248
rect 50376 21188 50380 21244
rect 50380 21188 50436 21244
rect 50436 21188 50440 21244
rect 50376 21184 50440 21188
rect 50456 21244 50520 21248
rect 50456 21188 50460 21244
rect 50460 21188 50516 21244
rect 50516 21188 50520 21244
rect 50456 21184 50520 21188
rect 50536 21244 50600 21248
rect 50536 21188 50540 21244
rect 50540 21188 50596 21244
rect 50596 21188 50600 21244
rect 50536 21184 50600 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 50296 20156 50360 20160
rect 50296 20100 50300 20156
rect 50300 20100 50356 20156
rect 50356 20100 50360 20156
rect 50296 20096 50360 20100
rect 50376 20156 50440 20160
rect 50376 20100 50380 20156
rect 50380 20100 50436 20156
rect 50436 20100 50440 20156
rect 50376 20096 50440 20100
rect 50456 20156 50520 20160
rect 50456 20100 50460 20156
rect 50460 20100 50516 20156
rect 50516 20100 50520 20156
rect 50456 20096 50520 20100
rect 50536 20156 50600 20160
rect 50536 20100 50540 20156
rect 50540 20100 50596 20156
rect 50596 20100 50600 20156
rect 50536 20096 50600 20100
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 50296 19068 50360 19072
rect 50296 19012 50300 19068
rect 50300 19012 50356 19068
rect 50356 19012 50360 19068
rect 50296 19008 50360 19012
rect 50376 19068 50440 19072
rect 50376 19012 50380 19068
rect 50380 19012 50436 19068
rect 50436 19012 50440 19068
rect 50376 19008 50440 19012
rect 50456 19068 50520 19072
rect 50456 19012 50460 19068
rect 50460 19012 50516 19068
rect 50516 19012 50520 19068
rect 50456 19008 50520 19012
rect 50536 19068 50600 19072
rect 50536 19012 50540 19068
rect 50540 19012 50596 19068
rect 50596 19012 50600 19068
rect 50536 19008 50600 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 50296 17980 50360 17984
rect 50296 17924 50300 17980
rect 50300 17924 50356 17980
rect 50356 17924 50360 17980
rect 50296 17920 50360 17924
rect 50376 17980 50440 17984
rect 50376 17924 50380 17980
rect 50380 17924 50436 17980
rect 50436 17924 50440 17980
rect 50376 17920 50440 17924
rect 50456 17980 50520 17984
rect 50456 17924 50460 17980
rect 50460 17924 50516 17980
rect 50516 17924 50520 17980
rect 50456 17920 50520 17924
rect 50536 17980 50600 17984
rect 50536 17924 50540 17980
rect 50540 17924 50596 17980
rect 50596 17924 50600 17980
rect 50536 17920 50600 17924
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 50296 16892 50360 16896
rect 50296 16836 50300 16892
rect 50300 16836 50356 16892
rect 50356 16836 50360 16892
rect 50296 16832 50360 16836
rect 50376 16892 50440 16896
rect 50376 16836 50380 16892
rect 50380 16836 50436 16892
rect 50436 16836 50440 16892
rect 50376 16832 50440 16836
rect 50456 16892 50520 16896
rect 50456 16836 50460 16892
rect 50460 16836 50516 16892
rect 50516 16836 50520 16892
rect 50456 16832 50520 16836
rect 50536 16892 50600 16896
rect 50536 16836 50540 16892
rect 50540 16836 50596 16892
rect 50596 16836 50600 16892
rect 50536 16832 50600 16836
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 50296 15804 50360 15808
rect 50296 15748 50300 15804
rect 50300 15748 50356 15804
rect 50356 15748 50360 15804
rect 50296 15744 50360 15748
rect 50376 15804 50440 15808
rect 50376 15748 50380 15804
rect 50380 15748 50436 15804
rect 50436 15748 50440 15804
rect 50376 15744 50440 15748
rect 50456 15804 50520 15808
rect 50456 15748 50460 15804
rect 50460 15748 50516 15804
rect 50516 15748 50520 15804
rect 50456 15744 50520 15748
rect 50536 15804 50600 15808
rect 50536 15748 50540 15804
rect 50540 15748 50596 15804
rect 50596 15748 50600 15804
rect 50536 15744 50600 15748
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 50296 14716 50360 14720
rect 50296 14660 50300 14716
rect 50300 14660 50356 14716
rect 50356 14660 50360 14716
rect 50296 14656 50360 14660
rect 50376 14716 50440 14720
rect 50376 14660 50380 14716
rect 50380 14660 50436 14716
rect 50436 14660 50440 14716
rect 50376 14656 50440 14660
rect 50456 14716 50520 14720
rect 50456 14660 50460 14716
rect 50460 14660 50516 14716
rect 50516 14660 50520 14716
rect 50456 14656 50520 14660
rect 50536 14716 50600 14720
rect 50536 14660 50540 14716
rect 50540 14660 50596 14716
rect 50596 14660 50600 14716
rect 50536 14656 50600 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 50296 13628 50360 13632
rect 50296 13572 50300 13628
rect 50300 13572 50356 13628
rect 50356 13572 50360 13628
rect 50296 13568 50360 13572
rect 50376 13628 50440 13632
rect 50376 13572 50380 13628
rect 50380 13572 50436 13628
rect 50436 13572 50440 13628
rect 50376 13568 50440 13572
rect 50456 13628 50520 13632
rect 50456 13572 50460 13628
rect 50460 13572 50516 13628
rect 50516 13572 50520 13628
rect 50456 13568 50520 13572
rect 50536 13628 50600 13632
rect 50536 13572 50540 13628
rect 50540 13572 50596 13628
rect 50596 13572 50600 13628
rect 50536 13568 50600 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 50296 12540 50360 12544
rect 50296 12484 50300 12540
rect 50300 12484 50356 12540
rect 50356 12484 50360 12540
rect 50296 12480 50360 12484
rect 50376 12540 50440 12544
rect 50376 12484 50380 12540
rect 50380 12484 50436 12540
rect 50436 12484 50440 12540
rect 50376 12480 50440 12484
rect 50456 12540 50520 12544
rect 50456 12484 50460 12540
rect 50460 12484 50516 12540
rect 50516 12484 50520 12540
rect 50456 12480 50520 12484
rect 50536 12540 50600 12544
rect 50536 12484 50540 12540
rect 50540 12484 50596 12540
rect 50596 12484 50600 12540
rect 50536 12480 50600 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 50296 11452 50360 11456
rect 50296 11396 50300 11452
rect 50300 11396 50356 11452
rect 50356 11396 50360 11452
rect 50296 11392 50360 11396
rect 50376 11452 50440 11456
rect 50376 11396 50380 11452
rect 50380 11396 50436 11452
rect 50436 11396 50440 11452
rect 50376 11392 50440 11396
rect 50456 11452 50520 11456
rect 50456 11396 50460 11452
rect 50460 11396 50516 11452
rect 50516 11396 50520 11452
rect 50456 11392 50520 11396
rect 50536 11452 50600 11456
rect 50536 11396 50540 11452
rect 50540 11396 50596 11452
rect 50596 11396 50600 11452
rect 50536 11392 50600 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 50296 10364 50360 10368
rect 50296 10308 50300 10364
rect 50300 10308 50356 10364
rect 50356 10308 50360 10364
rect 50296 10304 50360 10308
rect 50376 10364 50440 10368
rect 50376 10308 50380 10364
rect 50380 10308 50436 10364
rect 50436 10308 50440 10364
rect 50376 10304 50440 10308
rect 50456 10364 50520 10368
rect 50456 10308 50460 10364
rect 50460 10308 50516 10364
rect 50516 10308 50520 10364
rect 50456 10304 50520 10308
rect 50536 10364 50600 10368
rect 50536 10308 50540 10364
rect 50540 10308 50596 10364
rect 50596 10308 50600 10364
rect 50536 10304 50600 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 50296 9276 50360 9280
rect 50296 9220 50300 9276
rect 50300 9220 50356 9276
rect 50356 9220 50360 9276
rect 50296 9216 50360 9220
rect 50376 9276 50440 9280
rect 50376 9220 50380 9276
rect 50380 9220 50436 9276
rect 50436 9220 50440 9276
rect 50376 9216 50440 9220
rect 50456 9276 50520 9280
rect 50456 9220 50460 9276
rect 50460 9220 50516 9276
rect 50516 9220 50520 9276
rect 50456 9216 50520 9220
rect 50536 9276 50600 9280
rect 50536 9220 50540 9276
rect 50540 9220 50596 9276
rect 50596 9220 50600 9276
rect 50536 9216 50600 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 50296 8188 50360 8192
rect 50296 8132 50300 8188
rect 50300 8132 50356 8188
rect 50356 8132 50360 8188
rect 50296 8128 50360 8132
rect 50376 8188 50440 8192
rect 50376 8132 50380 8188
rect 50380 8132 50436 8188
rect 50436 8132 50440 8188
rect 50376 8128 50440 8132
rect 50456 8188 50520 8192
rect 50456 8132 50460 8188
rect 50460 8132 50516 8188
rect 50516 8132 50520 8188
rect 50456 8128 50520 8132
rect 50536 8188 50600 8192
rect 50536 8132 50540 8188
rect 50540 8132 50596 8188
rect 50596 8132 50600 8188
rect 50536 8128 50600 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 50296 7100 50360 7104
rect 50296 7044 50300 7100
rect 50300 7044 50356 7100
rect 50356 7044 50360 7100
rect 50296 7040 50360 7044
rect 50376 7100 50440 7104
rect 50376 7044 50380 7100
rect 50380 7044 50436 7100
rect 50436 7044 50440 7100
rect 50376 7040 50440 7044
rect 50456 7100 50520 7104
rect 50456 7044 50460 7100
rect 50460 7044 50516 7100
rect 50516 7044 50520 7100
rect 50456 7040 50520 7044
rect 50536 7100 50600 7104
rect 50536 7044 50540 7100
rect 50540 7044 50596 7100
rect 50596 7044 50600 7100
rect 50536 7040 50600 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 50296 6012 50360 6016
rect 50296 5956 50300 6012
rect 50300 5956 50356 6012
rect 50356 5956 50360 6012
rect 50296 5952 50360 5956
rect 50376 6012 50440 6016
rect 50376 5956 50380 6012
rect 50380 5956 50436 6012
rect 50436 5956 50440 6012
rect 50376 5952 50440 5956
rect 50456 6012 50520 6016
rect 50456 5956 50460 6012
rect 50460 5956 50516 6012
rect 50516 5956 50520 6012
rect 50456 5952 50520 5956
rect 50536 6012 50600 6016
rect 50536 5956 50540 6012
rect 50540 5956 50596 6012
rect 50596 5956 50600 6012
rect 50536 5952 50600 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 50296 4924 50360 4928
rect 50296 4868 50300 4924
rect 50300 4868 50356 4924
rect 50356 4868 50360 4924
rect 50296 4864 50360 4868
rect 50376 4924 50440 4928
rect 50376 4868 50380 4924
rect 50380 4868 50436 4924
rect 50436 4868 50440 4924
rect 50376 4864 50440 4868
rect 50456 4924 50520 4928
rect 50456 4868 50460 4924
rect 50460 4868 50516 4924
rect 50516 4868 50520 4924
rect 50456 4864 50520 4868
rect 50536 4924 50600 4928
rect 50536 4868 50540 4924
rect 50540 4868 50596 4924
rect 50596 4868 50600 4924
rect 50536 4864 50600 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 50296 3836 50360 3840
rect 50296 3780 50300 3836
rect 50300 3780 50356 3836
rect 50356 3780 50360 3836
rect 50296 3776 50360 3780
rect 50376 3836 50440 3840
rect 50376 3780 50380 3836
rect 50380 3780 50436 3836
rect 50436 3780 50440 3836
rect 50376 3776 50440 3780
rect 50456 3836 50520 3840
rect 50456 3780 50460 3836
rect 50460 3780 50516 3836
rect 50516 3780 50520 3836
rect 50456 3776 50520 3780
rect 50536 3836 50600 3840
rect 50536 3780 50540 3836
rect 50540 3780 50596 3836
rect 50596 3780 50600 3836
rect 50536 3776 50600 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 50296 2748 50360 2752
rect 50296 2692 50300 2748
rect 50300 2692 50356 2748
rect 50356 2692 50360 2748
rect 50296 2688 50360 2692
rect 50376 2748 50440 2752
rect 50376 2692 50380 2748
rect 50380 2692 50436 2748
rect 50436 2692 50440 2748
rect 50376 2688 50440 2692
rect 50456 2748 50520 2752
rect 50456 2692 50460 2748
rect 50460 2692 50516 2748
rect 50516 2692 50520 2748
rect 50456 2688 50520 2692
rect 50536 2748 50600 2752
rect 50536 2692 50540 2748
rect 50540 2692 50596 2748
rect 50596 2692 50600 2748
rect 50536 2688 50600 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
<< metal4 >>
rect 4208 57696 4528 57712
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5472 4528 6496
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4868 2176 5188 57664
rect 5528 2176 5848 57664
rect 6188 2176 6508 57664
rect 19568 57152 19888 57712
rect 34928 57696 35248 57712
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 50624 19888 51648
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 4208 2128 4528 2144
rect 19568 2128 19888 2688
rect 20228 2176 20548 57664
rect 20888 2176 21208 57664
rect 21548 2176 21868 57664
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5472 35248 6496
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 4384 35248 5408
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 35588 2176 35908 57664
rect 36248 2176 36568 57664
rect 36908 2176 37228 57664
rect 50288 57152 50608 57712
rect 50288 57088 50296 57152
rect 50360 57088 50376 57152
rect 50440 57088 50456 57152
rect 50520 57088 50536 57152
rect 50600 57088 50608 57152
rect 50288 56064 50608 57088
rect 50288 56000 50296 56064
rect 50360 56000 50376 56064
rect 50440 56000 50456 56064
rect 50520 56000 50536 56064
rect 50600 56000 50608 56064
rect 50288 54976 50608 56000
rect 50288 54912 50296 54976
rect 50360 54912 50376 54976
rect 50440 54912 50456 54976
rect 50520 54912 50536 54976
rect 50600 54912 50608 54976
rect 50288 53888 50608 54912
rect 50288 53824 50296 53888
rect 50360 53824 50376 53888
rect 50440 53824 50456 53888
rect 50520 53824 50536 53888
rect 50600 53824 50608 53888
rect 50288 52800 50608 53824
rect 50288 52736 50296 52800
rect 50360 52736 50376 52800
rect 50440 52736 50456 52800
rect 50520 52736 50536 52800
rect 50600 52736 50608 52800
rect 50288 51712 50608 52736
rect 50288 51648 50296 51712
rect 50360 51648 50376 51712
rect 50440 51648 50456 51712
rect 50520 51648 50536 51712
rect 50600 51648 50608 51712
rect 50288 50624 50608 51648
rect 50288 50560 50296 50624
rect 50360 50560 50376 50624
rect 50440 50560 50456 50624
rect 50520 50560 50536 50624
rect 50600 50560 50608 50624
rect 50288 49536 50608 50560
rect 50288 49472 50296 49536
rect 50360 49472 50376 49536
rect 50440 49472 50456 49536
rect 50520 49472 50536 49536
rect 50600 49472 50608 49536
rect 50288 48448 50608 49472
rect 50288 48384 50296 48448
rect 50360 48384 50376 48448
rect 50440 48384 50456 48448
rect 50520 48384 50536 48448
rect 50600 48384 50608 48448
rect 50288 47360 50608 48384
rect 50288 47296 50296 47360
rect 50360 47296 50376 47360
rect 50440 47296 50456 47360
rect 50520 47296 50536 47360
rect 50600 47296 50608 47360
rect 50288 46272 50608 47296
rect 50288 46208 50296 46272
rect 50360 46208 50376 46272
rect 50440 46208 50456 46272
rect 50520 46208 50536 46272
rect 50600 46208 50608 46272
rect 50288 45184 50608 46208
rect 50288 45120 50296 45184
rect 50360 45120 50376 45184
rect 50440 45120 50456 45184
rect 50520 45120 50536 45184
rect 50600 45120 50608 45184
rect 50288 44096 50608 45120
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33216 50608 34240
rect 50288 33152 50296 33216
rect 50360 33152 50376 33216
rect 50440 33152 50456 33216
rect 50520 33152 50536 33216
rect 50600 33152 50608 33216
rect 50288 32128 50608 33152
rect 50288 32064 50296 32128
rect 50360 32064 50376 32128
rect 50440 32064 50456 32128
rect 50520 32064 50536 32128
rect 50600 32064 50608 32128
rect 50288 31040 50608 32064
rect 50288 30976 50296 31040
rect 50360 30976 50376 31040
rect 50440 30976 50456 31040
rect 50520 30976 50536 31040
rect 50600 30976 50608 31040
rect 50288 29952 50608 30976
rect 50288 29888 50296 29952
rect 50360 29888 50376 29952
rect 50440 29888 50456 29952
rect 50520 29888 50536 29952
rect 50600 29888 50608 29952
rect 50288 28864 50608 29888
rect 50288 28800 50296 28864
rect 50360 28800 50376 28864
rect 50440 28800 50456 28864
rect 50520 28800 50536 28864
rect 50600 28800 50608 28864
rect 50288 27776 50608 28800
rect 50288 27712 50296 27776
rect 50360 27712 50376 27776
rect 50440 27712 50456 27776
rect 50520 27712 50536 27776
rect 50600 27712 50608 27776
rect 50288 26688 50608 27712
rect 50288 26624 50296 26688
rect 50360 26624 50376 26688
rect 50440 26624 50456 26688
rect 50520 26624 50536 26688
rect 50600 26624 50608 26688
rect 50288 25600 50608 26624
rect 50288 25536 50296 25600
rect 50360 25536 50376 25600
rect 50440 25536 50456 25600
rect 50520 25536 50536 25600
rect 50600 25536 50608 25600
rect 50288 24512 50608 25536
rect 50288 24448 50296 24512
rect 50360 24448 50376 24512
rect 50440 24448 50456 24512
rect 50520 24448 50536 24512
rect 50600 24448 50608 24512
rect 50288 23424 50608 24448
rect 50288 23360 50296 23424
rect 50360 23360 50376 23424
rect 50440 23360 50456 23424
rect 50520 23360 50536 23424
rect 50600 23360 50608 23424
rect 50288 22336 50608 23360
rect 50288 22272 50296 22336
rect 50360 22272 50376 22336
rect 50440 22272 50456 22336
rect 50520 22272 50536 22336
rect 50600 22272 50608 22336
rect 50288 21248 50608 22272
rect 50288 21184 50296 21248
rect 50360 21184 50376 21248
rect 50440 21184 50456 21248
rect 50520 21184 50536 21248
rect 50600 21184 50608 21248
rect 50288 20160 50608 21184
rect 50288 20096 50296 20160
rect 50360 20096 50376 20160
rect 50440 20096 50456 20160
rect 50520 20096 50536 20160
rect 50600 20096 50608 20160
rect 50288 19072 50608 20096
rect 50288 19008 50296 19072
rect 50360 19008 50376 19072
rect 50440 19008 50456 19072
rect 50520 19008 50536 19072
rect 50600 19008 50608 19072
rect 50288 17984 50608 19008
rect 50288 17920 50296 17984
rect 50360 17920 50376 17984
rect 50440 17920 50456 17984
rect 50520 17920 50536 17984
rect 50600 17920 50608 17984
rect 50288 16896 50608 17920
rect 50288 16832 50296 16896
rect 50360 16832 50376 16896
rect 50440 16832 50456 16896
rect 50520 16832 50536 16896
rect 50600 16832 50608 16896
rect 50288 15808 50608 16832
rect 50288 15744 50296 15808
rect 50360 15744 50376 15808
rect 50440 15744 50456 15808
rect 50520 15744 50536 15808
rect 50600 15744 50608 15808
rect 50288 14720 50608 15744
rect 50288 14656 50296 14720
rect 50360 14656 50376 14720
rect 50440 14656 50456 14720
rect 50520 14656 50536 14720
rect 50600 14656 50608 14720
rect 50288 13632 50608 14656
rect 50288 13568 50296 13632
rect 50360 13568 50376 13632
rect 50440 13568 50456 13632
rect 50520 13568 50536 13632
rect 50600 13568 50608 13632
rect 50288 12544 50608 13568
rect 50288 12480 50296 12544
rect 50360 12480 50376 12544
rect 50440 12480 50456 12544
rect 50520 12480 50536 12544
rect 50600 12480 50608 12544
rect 50288 11456 50608 12480
rect 50288 11392 50296 11456
rect 50360 11392 50376 11456
rect 50440 11392 50456 11456
rect 50520 11392 50536 11456
rect 50600 11392 50608 11456
rect 50288 10368 50608 11392
rect 50288 10304 50296 10368
rect 50360 10304 50376 10368
rect 50440 10304 50456 10368
rect 50520 10304 50536 10368
rect 50600 10304 50608 10368
rect 50288 9280 50608 10304
rect 50288 9216 50296 9280
rect 50360 9216 50376 9280
rect 50440 9216 50456 9280
rect 50520 9216 50536 9280
rect 50600 9216 50608 9280
rect 50288 8192 50608 9216
rect 50288 8128 50296 8192
rect 50360 8128 50376 8192
rect 50440 8128 50456 8192
rect 50520 8128 50536 8192
rect 50600 8128 50608 8192
rect 50288 7104 50608 8128
rect 50288 7040 50296 7104
rect 50360 7040 50376 7104
rect 50440 7040 50456 7104
rect 50520 7040 50536 7104
rect 50600 7040 50608 7104
rect 50288 6016 50608 7040
rect 50288 5952 50296 6016
rect 50360 5952 50376 6016
rect 50440 5952 50456 6016
rect 50520 5952 50536 6016
rect 50600 5952 50608 6016
rect 50288 4928 50608 5952
rect 50288 4864 50296 4928
rect 50360 4864 50376 4928
rect 50440 4864 50456 4928
rect 50520 4864 50536 4928
rect 50600 4864 50608 4928
rect 50288 3840 50608 4864
rect 50288 3776 50296 3840
rect 50360 3776 50376 3840
rect 50440 3776 50456 3840
rect 50520 3776 50536 3840
rect 50600 3776 50608 3840
rect 50288 2752 50608 3776
rect 50288 2688 50296 2752
rect 50360 2688 50376 2752
rect 50440 2688 50456 2752
rect 50520 2688 50536 2752
rect 50600 2688 50608 2752
rect 34928 2128 35248 2144
rect 50288 2128 50608 2688
rect 50948 2176 51268 57664
rect 51608 2176 51928 57664
rect 52268 2176 52588 57664
use sky130_fd_sc_hd__decap_4  FILLER_1_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1564 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1621523292
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1621523292
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1621523292
transform 1 0 2300 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output300 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output289
timestamp 1621523292
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output314
timestamp 1621523292
transform 1 0 2852 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1621523292
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1621523292
transform 1 0 3220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1621523292
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4508 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1621523292
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1621523292
transform 1 0 4232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1621523292
transform 1 0 4232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4508 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_49
timestamp 1621523292
transform 1 0 5612 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1621523292
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46
timestamp 1621523292
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1621523292
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1621523292
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1621523292
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1621523292
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1621523292
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1621523292
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1621523292
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1621523292
transform 1 0 7820 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1621523292
transform 1 0 8464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66
timestamp 1621523292
transform 1 0 7176 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72
timestamp 1621523292
transform 1 0 7728 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76
timestamp 1621523292
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1621523292
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1621523292
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1621523292
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1621523292
transform 1 0 9660 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1621523292
transform 1 0 10580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_88
timestamp 1621523292
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1621523292
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96
timestamp 1621523292
transform 1 0 9936 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102
timestamp 1621523292
transform 1 0 10488 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_106
timestamp 1621523292
transform 1 0 10856 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1621523292
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106
timestamp 1621523292
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1621523292
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_114
timestamp 1621523292
transform 1 0 11592 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1621523292
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1621523292
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_131
timestamp 1621523292
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_124
timestamp 1621523292
transform 1 0 12512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1621523292
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1621523292
transform 1 0 12236 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1621523292
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1621523292
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1621523292
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1621523292
transform 1 0 13524 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1621523292
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_138
timestamp 1621523292
transform 1 0 13800 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1621523292
transform 1 0 14352 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1621523292
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1621523292
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1621523292
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1621523292
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_160
timestamp 1621523292
transform 1 0 15824 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_153
timestamp 1621523292
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1621523292
transform 1 0 15548 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1621523292
transform 1 0 17020 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_167
timestamp 1621523292
transform 1 0 16468 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1621523292
transform 1 0 16192 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1621523292
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1621523292
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1621523292
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1621523292
transform 1 0 17572 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1621523292
transform 1 0 18216 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1621523292
transform 1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1621523292
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1621523292
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_189
timestamp 1621523292
transform 1 0 18492 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_196
timestamp 1621523292
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1621523292
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1621523292
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1621523292
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1621523292
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1621523292
transform 1 0 20884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_202
timestamp 1621523292
transform 1 0 19688 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1621523292
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_211
timestamp 1621523292
transform 1 0 20516 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1621523292
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1621523292
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_220
timestamp 1621523292
transform 1 0 21344 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_226
timestamp 1621523292
transform 1 0 21896 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1621523292
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1621523292
transform 1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1621523292
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1621523292
transform 1 0 23184 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1621523292
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1621523292
transform 1 0 22908 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1621523292
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_229
timestamp 1621523292
transform 1 0 22172 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1621523292
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1621523292
transform 1 0 23552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1621523292
transform 1 0 24380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_247
timestamp 1621523292
transform 1 0 23828 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1621523292
transform 1 0 24656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_260
timestamp 1621523292
transform 1 0 25024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1621523292
transform 1 0 25208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_241
timestamp 1621523292
transform 1 0 23276 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_253
timestamp 1621523292
transform 1 0 24380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1621523292
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1621523292
transform 1 0 26220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1621523292
transform 1 0 27140 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1621523292
transform 1 0 25852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_276
timestamp 1621523292
transform 1 0 26496 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_282
timestamp 1621523292
transform 1 0 27048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_265
timestamp 1621523292
transform 1 0 25484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_277
timestamp 1621523292
transform 1 0 26588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_292
timestamp 1621523292
transform 1 0 27968 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_286
timestamp 1621523292
transform 1 0 27416 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1621523292
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1621523292
transform 1 0 27416 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1621523292
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1621523292
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1621523292
transform 1 0 28336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_300
timestamp 1621523292
transform 1 0 28704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_295
timestamp 1621523292
transform 1 0 28244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output256
timestamp 1621523292
transform 1 0 28336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1621523292
transform 1 0 28704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1621523292
transform 1 0 28060 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1621523292
transform 1 0 28980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 29072 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1621523292
transform 1 0 29624 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_312
timestamp 1621523292
transform 1 0 29808 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _2225_
timestamp 1621523292
transform 1 0 29992 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1714_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 29348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_322
timestamp 1621523292
transform 1 0 30728 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1621523292
transform 1 0 30544 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_318
timestamp 1621523292
transform 1 0 30360 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1621523292
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2226_
timestamp 1621523292
transform 1 0 30912 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1671_
timestamp 1621523292
transform 1 0 31096 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_333
timestamp 1621523292
transform 1 0 31740 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_329
timestamp 1621523292
transform 1 0 31372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1621523292
transform 1 0 31648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output278
timestamp 1621523292
transform 1 0 31832 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output267
timestamp 1621523292
transform 1 0 32016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1621523292
transform 1 0 32660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_338
timestamp 1621523292
transform 1 0 32200 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_340
timestamp 1621523292
transform 1 0 32384 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1621523292
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1621523292
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1621523292
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2227_
timestamp 1621523292
transform 1 0 33028 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1664_
timestamp 1621523292
transform 1 0 34132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2228_
timestamp 1621523292
transform 1 0 33580 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2229_
timestamp 1621523292
transform 1 0 34684 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2230_
timestamp 1621523292
transform 1 0 34776 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_361
timestamp 1621523292
transform 1 0 34316 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1621523292
transform 1 0 33764 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_362
timestamp 1621523292
transform 1 0 34408 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_374
timestamp 1621523292
transform 1 0 35512 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1621523292
transform 1 0 35880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1621523292
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output283
timestamp 1621523292
transform 1 0 35880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1621523292
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_382
timestamp 1621523292
transform 1 0 36248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output285
timestamp 1621523292
transform 1 0 36616 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2231_
timestamp 1621523292
transform 1 0 36248 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_390
timestamp 1621523292
transform 1 0 36984 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_390
timestamp 1621523292
transform 1 0 36984 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2232_
timestamp 1621523292
transform 1 0 37352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2233_
timestamp 1621523292
transform 1 0 38272 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1621523292
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1621523292
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1621523292
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_407
timestamp 1621523292
transform 1 0 38548 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_398
timestamp 1621523292
transform 1 0 37720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_400
timestamp 1621523292
transform 1 0 37904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_412
timestamp 1621523292
transform 1 0 39008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_415
timestamp 1621523292
transform 1 0 39284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _2235_
timestamp 1621523292
transform 1 0 39468 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2234_
timestamp 1621523292
transform 1 0 39376 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1621523292
transform 1 0 40112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_425
timestamp 1621523292
transform 1 0 40204 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2236_
timestamp 1621523292
transform 1 0 40480 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_436
timestamp 1621523292
transform 1 0 41216 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_436
timestamp 1621523292
transform 1 0 41216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_433
timestamp 1621523292
transform 1 0 40940 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1621523292
transform 1 0 41124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2237_
timestamp 1621523292
transform 1 0 41584 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2238_
timestamp 1621523292
transform 1 0 42688 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1621523292
transform 1 0 43056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output259
timestamp 1621523292
transform 1 0 41584 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output260
timestamp 1621523292
transform 1 0 42320 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_448
timestamp 1621523292
transform 1 0 42320 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1621523292
transform 1 0 41952 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1621523292
transform 1 0 42688 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1621523292
transform 1 0 43148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2239_
timestamp 1621523292
transform 1 0 43516 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2240_
timestamp 1621523292
transform 1 0 44252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1621523292
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output262
timestamp 1621523292
transform 1 0 44620 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_460
timestamp 1621523292
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_465
timestamp 1621523292
transform 1 0 43884 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1621523292
transform 1 0 44988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_469
timestamp 1621523292
transform 1 0 44252 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_477
timestamp 1621523292
transform 1 0 44988 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_485
timestamp 1621523292
transform 1 0 45724 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1621523292
transform 1 0 46092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output264
timestamp 1621523292
transform 1 0 46092 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output263
timestamp 1621523292
transform 1 0 45356 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2241_
timestamp 1621523292
transform 1 0 45356 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_497
timestamp 1621523292
transform 1 0 46828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_493
timestamp 1621523292
transform 1 0 46460 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1621523292
transform 1 0 46552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1621523292
transform 1 0 46460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2243_
timestamp 1621523292
transform 1 0 46920 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2242_
timestamp 1621523292
transform 1 0 46920 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_506
timestamp 1621523292
transform 1 0 47656 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_506
timestamp 1621523292
transform 1 0 47656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2244_
timestamp 1621523292
transform 1 0 48024 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_514
timestamp 1621523292
transform 1 0 48392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_512
timestamp 1621523292
transform 1 0 48208 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_518
timestamp 1621523292
transform 1 0 48760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1621523292
transform 1 0 48300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2245_
timestamp 1621523292
transform 1 0 48760 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_523
timestamp 1621523292
transform 1 0 49220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1621523292
transform 1 0 49128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2246_
timestamp 1621523292
transform 1 0 49588 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2247_
timestamp 1621523292
transform 1 0 50784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output265
timestamp 1621523292
transform 1 0 50692 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output269
timestamp 1621523292
transform 1 0 49864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_535
timestamp 1621523292
transform 1 0 50324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_543
timestamp 1621523292
transform 1 0 51060 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_526
timestamp 1621523292
transform 1 0 49496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_534
timestamp 1621523292
transform 1 0 50232 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _2248_
timestamp 1621523292
transform 1 0 52256 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2249_
timestamp 1621523292
transform 1 0 52164 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1621523292
transform 1 0 51796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_552
timestamp 1621523292
transform 1 0 51888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_564
timestamp 1621523292
transform 1 0 52992 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_548
timestamp 1621523292
transform 1 0 51520 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_554
timestamp 1621523292
transform 1 0 52072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_563
timestamp 1621523292
transform 1 0 52900 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1621523292
transform 1 0 53636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_569
timestamp 1621523292
transform 1 0 53452 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_576
timestamp 1621523292
transform 1 0 54096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output254
timestamp 1621523292
transform 1 0 53728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1621523292
transform 1 0 53544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2251_
timestamp 1621523292
transform 1 0 54004 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_583
timestamp 1621523292
transform 1 0 54740 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_581
timestamp 1621523292
transform 1 0 54556 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1621523292
transform 1 0 54464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output215
timestamp 1621523292
transform 1 0 55292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2252_
timestamp 1621523292
transform 1 0 55108 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2253_
timestamp 1621523292
transform 1 0 56212 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2255_
timestamp 1621523292
transform 1 0 56028 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1621523292
transform 1 0 57132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1621523292
transform 1 0 55660 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_605
timestamp 1621523292
transform 1 0 56764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_610
timestamp 1621523292
transform 1 0 57224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_595
timestamp 1621523292
transform 1 0 55844 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_607
timestamp 1621523292
transform 1 0 56948 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _2256_
timestamp 1621523292
transform 1 0 57500 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1621523292
transform -1 0 58880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1621523292
transform -1 0 58880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output177
timestamp 1621523292
transform 1 0 57868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_616
timestamp 1621523292
transform 1 0 57776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1621523292
transform 1 0 58236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1621523292
transform 1 0 58236 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1621523292
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1621523292
transform 1 0 2852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output311
timestamp 1621523292
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1621523292
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_11
timestamp 1621523292
transform 1 0 2116 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1621523292
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_22
timestamp 1621523292
transform 1 0 3128 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1621523292
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1621523292
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1621523292
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1621523292
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1621523292
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1621523292
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1621523292
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1621523292
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_2  _2192_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_99
timestamp 1621523292
transform 1 0 10212 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1621523292
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1715_
timestamp 1621523292
transform 1 0 12328 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1621523292
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_125
timestamp 1621523292
transform 1 0 12604 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1621523292
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_137
timestamp 1621523292
transform 1 0 13708 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1621523292
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1621523292
transform 1 0 15456 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1621523292
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1621523292
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1621523292
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1621523292
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1621523292
transform 1 0 19596 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_213
timestamp 1621523292
transform 1 0 20700 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1621523292
transform 1 0 21804 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_237
timestamp 1621523292
transform 1 0 22908 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1621523292
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_249
timestamp 1621523292
transform 1 0 24012 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1621523292
transform 1 0 24840 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_270
timestamp 1621523292
transform 1 0 25944 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_282
timestamp 1621523292
transform 1 0 27048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_294
timestamp 1621523292
transform 1 0 28152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1672_
timestamp 1621523292
transform 1 0 30452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2106_
timestamp 1621523292
transform 1 0 31096 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1621523292
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1621523292
transform 1 0 29532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1621523292
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1621523292
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1621523292
transform 1 0 30728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1668_
timestamp 1621523292
transform 1 0 32108 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output281
timestamp 1621523292
transform 1 0 32752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_329
timestamp 1621523292
transform 1 0 31372 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1621523292
transform 1 0 32384 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_348
timestamp 1621523292
transform 1 0 33120 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1665_
timestamp 1621523292
transform 1 0 34592 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1621523292
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output282
timestamp 1621523292
transform 1 0 33672 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1621523292
transform 1 0 34040 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_367
timestamp 1621523292
transform 1 0 34868 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1657_
timestamp 1621523292
transform 1 0 36708 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output284
timestamp 1621523292
transform 1 0 35696 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1621523292
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_380
timestamp 1621523292
transform 1 0 36064 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_386
timestamp 1621523292
transform 1 0 36616 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_390
timestamp 1621523292
transform 1 0 36984 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output257
timestamp 1621523292
transform 1 0 39192 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output286
timestamp 1621523292
transform 1 0 37352 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output287
timestamp 1621523292
transform 1 0 38272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_398
timestamp 1621523292
transform 1 0 37720 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_408
timestamp 1621523292
transform 1 0 38640 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1621523292
transform 1 0 40480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output258
timestamp 1621523292
transform 1 0 40940 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_418
timestamp 1621523292
transform 1 0 39560 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_426
timestamp 1621523292
transform 1 0 40296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1621523292
transform 1 0 40572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1655_
timestamp 1621523292
transform 1 0 42228 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output261
timestamp 1621523292
transform 1 0 42872 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_437
timestamp 1621523292
transform 1 0 41308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_445
timestamp 1621523292
transform 1 0 42044 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_450
timestamp 1621523292
transform 1 0 42504 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_458
timestamp 1621523292
transform 1 0 43240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1651_
timestamp 1621523292
transform 1 0 43700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1652_
timestamp 1621523292
transform 1 0 44528 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_462
timestamp 1621523292
transform 1 0 43608 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_466
timestamp 1621523292
transform 1 0 43976 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_475
timestamp 1621523292
transform 1 0 44804 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1621523292
transform 1 0 46828 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1650_
timestamp 1621523292
transform 1 0 46184 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1621523292
transform 1 0 45724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_483
timestamp 1621523292
transform 1 0 45540 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_486
timestamp 1621523292
transform 1 0 45816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_493
timestamp 1621523292
transform 1 0 46460 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_500
timestamp 1621523292
transform 1 0 47104 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output266
timestamp 1621523292
transform 1 0 47472 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output268
timestamp 1621523292
transform 1 0 48392 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_508
timestamp 1621523292
transform 1 0 47840 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_518
timestamp 1621523292
transform 1 0 48760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1644_
timestamp 1621523292
transform 1 0 49588 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1621523292
transform 1 0 50968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output270
timestamp 1621523292
transform 1 0 50232 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_526
timestamp 1621523292
transform 1 0 49496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_530
timestamp 1621523292
transform 1 0 49864 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_538
timestamp 1621523292
transform 1 0 50600 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_543
timestamp 1621523292
transform 1 0 51060 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2250_
timestamp 1621523292
transform 1 0 53084 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output271
timestamp 1621523292
transform 1 0 51428 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output272
timestamp 1621523292
transform 1 0 52164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1621523292
transform 1 0 51796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_559
timestamp 1621523292
transform 1 0 52532 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output273
timestamp 1621523292
transform 1 0 54188 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_573
timestamp 1621523292
transform 1 0 53820 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_581
timestamp 1621523292
transform 1 0 54556 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_589
timestamp 1621523292
transform 1 0 55292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1586_
timestamp 1621523292
transform 1 0 56672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2294_
timestamp 1621523292
transform 1 0 57316 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1621523292
transform 1 0 56212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output226
timestamp 1621523292
transform 1 0 55476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_595
timestamp 1621523292
transform 1 0 55844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_600
timestamp 1621523292
transform 1 0 56304 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_607
timestamp 1621523292
transform 1 0 56948 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1621523292
transform -1 0 58880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_619
timestamp 1621523292
transform 1 0 58052 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1621523292
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output315
timestamp 1621523292
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1621523292
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_11
timestamp 1621523292
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_23
timestamp 1621523292
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_35
timestamp 1621523292
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1621523292
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1621523292
transform 1 0 5428 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1621523292
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1621523292
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1621523292
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1621523292
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1621523292
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1621523292
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1621523292
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1621523292
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1621523292
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1621523292
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1621523292
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1621523292
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1621523292
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1621523292
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1621523292
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1621523292
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1621523292
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1621523292
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_220
timestamp 1621523292
transform 1 0 21344 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_229
timestamp 1621523292
transform 1 0 22172 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_241
timestamp 1621523292
transform 1 0 23276 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1621523292
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_265
timestamp 1621523292
transform 1 0 25484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_277
timestamp 1621523292
transform 1 0 26588 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1621523292
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_286
timestamp 1621523292
transform 1 0 27416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_298
timestamp 1621523292
transform 1 0 28520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2105_
timestamp 1621523292
transform 1 0 30084 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_310
timestamp 1621523292
transform 1 0 29624 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_314
timestamp 1621523292
transform 1 0 29992 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1621523292
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1667_
timestamp 1621523292
transform 1 0 33028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2107_
timestamp 1621523292
transform 1 0 31924 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1621523292
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_330
timestamp 1621523292
transform 1 0 31464 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_334
timestamp 1621523292
transform 1 0 31832 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_338
timestamp 1621523292
transform 1 0 32200 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_343
timestamp 1621523292
transform 1 0 32660 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1666_
timestamp 1621523292
transform 1 0 33948 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2109_
timestamp 1621523292
transform 1 0 34592 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2110_
timestamp 1621523292
transform 1 0 35236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_350
timestamp 1621523292
transform 1 0 33304 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_356
timestamp 1621523292
transform 1 0 33856 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_360
timestamp 1621523292
transform 1 0 34224 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_367
timestamp 1621523292
transform 1 0 34868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1662_
timestamp 1621523292
transform 1 0 37168 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1663_
timestamp 1621523292
transform 1 0 36064 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_374
timestamp 1621523292
transform 1 0 35512 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_383
timestamp 1621523292
transform 1 0 36340 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1621523292
transform 1 0 37076 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1660_
timestamp 1621523292
transform 1 0 38640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1621523292
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1621523292
transform 1 0 37444 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_400
timestamp 1621523292
transform 1 0 37904 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_411
timestamp 1621523292
transform 1 0 38916 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1658_
timestamp 1621523292
transform 1 0 39744 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1659_
timestamp 1621523292
transform 1 0 40388 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2116_
timestamp 1621523292
transform 1 0 41032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_419
timestamp 1621523292
transform 1 0 39652 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_423
timestamp 1621523292
transform 1 0 40020 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_430
timestamp 1621523292
transform 1 0 40664 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1656_
timestamp 1621523292
transform 1 0 41860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1621523292
transform 1 0 43056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_437
timestamp 1621523292
transform 1 0 41308 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_446
timestamp 1621523292
transform 1 0 42136 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_454
timestamp 1621523292
transform 1 0 42872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_457
timestamp 1621523292
transform 1 0 43148 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1621523292
transform 1 0 44252 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1654_
timestamp 1621523292
transform 1 0 43516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2120_
timestamp 1621523292
transform 1 0 44896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_464
timestamp 1621523292
transform 1 0 43792 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_468
timestamp 1621523292
transform 1 0 44160 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_472
timestamp 1621523292
transform 1 0 44528 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_479
timestamp 1621523292
transform 1 0 45172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1621523292
transform 1 0 46736 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2121_
timestamp 1621523292
transform 1 0 45540 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_486
timestamp 1621523292
transform 1 0 45816 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_494
timestamp 1621523292
transform 1 0 46552 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_499
timestamp 1621523292
transform 1 0 47012 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1645_
timestamp 1621523292
transform 1 0 47656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1646_
timestamp 1621523292
transform 1 0 48944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1621523292
transform 1 0 48300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_505
timestamp 1621523292
transform 1 0 47564 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_509
timestamp 1621523292
transform 1 0 47932 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_514
timestamp 1621523292
transform 1 0 48392 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_523
timestamp 1621523292
transform 1 0 49220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1638_
timestamp 1621523292
transform 1 0 49588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1639_
timestamp 1621523292
transform 1 0 50324 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1643_
timestamp 1621523292
transform 1 0 50968 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_531
timestamp 1621523292
transform 1 0 49956 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_538
timestamp 1621523292
transform 1 0 50600 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_545
timestamp 1621523292
transform 1 0 51244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1633_
timestamp 1621523292
transform 1 0 52900 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1634_
timestamp 1621523292
transform 1 0 52256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1640_
timestamp 1621523292
transform 1 0 51612 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_552
timestamp 1621523292
transform 1 0 51888 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_559
timestamp 1621523292
transform 1 0 52532 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_566
timestamp 1621523292
transform 1 0 53176 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1621523292
transform 1 0 53544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output274
timestamp 1621523292
transform 1 0 54004 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output275
timestamp 1621523292
transform 1 0 54832 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1621523292
transform 1 0 53636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_579
timestamp 1621523292
transform 1 0 54372 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_583
timestamp 1621523292
transform 1 0 54740 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_588
timestamp 1621523292
transform 1 0 55200 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1587_
timestamp 1621523292
transform 1 0 55568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2254_
timestamp 1621523292
transform 1 0 56212 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_595
timestamp 1621523292
transform 1 0 55844 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_607
timestamp 1621523292
transform 1 0 56948 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1621523292
transform -1 0 58880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output188
timestamp 1621523292
transform 1 0 57868 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_615
timestamp 1621523292
transform 1 0 57684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1621523292
transform 1 0 58236 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1621523292
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1621523292
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1621523292
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1621523292
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1621523292
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1621523292
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1621523292
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1621523292
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1621523292
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1621523292
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1621523292
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1621523292
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1621523292
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1621523292
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1621523292
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1621523292
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1621523292
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1621523292
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1621523292
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1621523292
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1621523292
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1621523292
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1621523292
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1621523292
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_213
timestamp 1621523292
transform 1 0 20700 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1621523292
transform 1 0 21804 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1621523292
transform 1 0 22908 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1621523292
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_249
timestamp 1621523292
transform 1 0 24012 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1621523292
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_270
timestamp 1621523292
transform 1 0 25944 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_282
timestamp 1621523292
transform 1 0 27048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_294
timestamp 1621523292
transform 1 0 28152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1621523292
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_306
timestamp 1621523292
transform 1 0 29256 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_315
timestamp 1621523292
transform 1 0 30084 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_327
timestamp 1621523292
transform 1 0 31188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2108_
timestamp 1621523292
transform 1 0 32752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_339
timestamp 1621523292
transform 1 0 32292 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_343
timestamp 1621523292
transform 1 0 32660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_347
timestamp 1621523292
transform 1 0 33028 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1621523292
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_359
timestamp 1621523292
transform 1 0 34132 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2111_
timestamp 1621523292
transform 1 0 35880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2112_
timestamp 1621523292
transform 1 0 36800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_372
timestamp 1621523292
transform 1 0 35328 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_381
timestamp 1621523292
transform 1 0 36156 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_387
timestamp 1621523292
transform 1 0 36708 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_391
timestamp 1621523292
transform 1 0 37076 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1621523292
transform 1 0 37720 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2113_
timestamp 1621523292
transform 1 0 38364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2114_
timestamp 1621523292
transform 1 0 39008 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_397
timestamp 1621523292
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_401
timestamp 1621523292
transform 1 0 37996 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_408
timestamp 1621523292
transform 1 0 38640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2115_
timestamp 1621523292
transform 1 0 39652 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1621523292
transform 1 0 40480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_415
timestamp 1621523292
transform 1 0 39284 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_422
timestamp 1621523292
transform 1 0 39928 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_429
timestamp 1621523292
transform 1 0 40572 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2117_
timestamp 1621523292
transform 1 0 41308 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2118_
timestamp 1621523292
transform 1 0 42136 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2119_
timestamp 1621523292
transform 1 0 43240 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_440
timestamp 1621523292
transform 1 0 41584 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_449
timestamp 1621523292
transform 1 0 42412 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_457
timestamp 1621523292
transform 1 0 43148 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_461
timestamp 1621523292
transform 1 0 43516 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_473
timestamp 1621523292
transform 1 0 44620 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2122_
timestamp 1621523292
transform 1 0 46184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2123_
timestamp 1621523292
transform 1 0 46828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1621523292
transform 1 0 45724 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_486
timestamp 1621523292
transform 1 0 45816 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_493
timestamp 1621523292
transform 1 0 46460 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_500
timestamp 1621523292
transform 1 0 47104 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1621523292
transform 1 0 48760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2124_
timestamp 1621523292
transform 1 0 47840 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_511
timestamp 1621523292
transform 1 0 48116 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_517
timestamp 1621523292
transform 1 0 48668 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_521
timestamp 1621523292
transform 1 0 49036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2125_
timestamp 1621523292
transform 1 0 49404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2126_
timestamp 1621523292
transform 1 0 50048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1621523292
transform 1 0 50968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1621523292
transform 1 0 49680 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_535
timestamp 1621523292
transform 1 0 50324 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_541
timestamp 1621523292
transform 1 0 50876 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_543
timestamp 1621523292
transform 1 0 51060 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1635_
timestamp 1621523292
transform 1 0 52992 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1637_
timestamp 1621523292
transform 1 0 52348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1642_
timestamp 1621523292
transform 1 0 51704 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_549
timestamp 1621523292
transform 1 0 51612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_553
timestamp 1621523292
transform 1 0 51980 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_560
timestamp 1621523292
transform 1 0 52624 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_567
timestamp 1621523292
transform 1 0 53268 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2257_
timestamp 1621523292
transform 1 0 55108 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output277
timestamp 1621523292
transform 1 0 54372 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output280
timestamp 1621523292
transform 1 0 53636 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_575
timestamp 1621523292
transform 1 0 54004 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_583
timestamp 1621523292
transform 1 0 54740 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1621523292
transform 1 0 56212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output199
timestamp 1621523292
transform 1 0 56764 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_595
timestamp 1621523292
transform 1 0 55844 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_600
timestamp 1621523292
transform 1 0 56304 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_604
timestamp 1621523292
transform 1 0 56672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_609
timestamp 1621523292
transform 1 0 57132 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2295_
timestamp 1621523292
transform 1 0 57500 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1621523292
transform -1 0 58880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1621523292
transform 1 0 58236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1621523292
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output316
timestamp 1621523292
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1621523292
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_11
timestamp 1621523292
transform 1 0 2116 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_23
timestamp 1621523292
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_35
timestamp 1621523292
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1621523292
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1621523292
transform 1 0 5428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1621523292
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1621523292
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1621523292
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1621523292
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1621523292
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1621523292
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1621523292
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1621523292
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1621523292
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1621523292
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1621523292
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1621523292
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1621523292
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1621523292
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1621523292
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1621523292
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1621523292
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1621523292
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_220
timestamp 1621523292
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_229
timestamp 1621523292
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_241
timestamp 1621523292
transform 1 0 23276 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_253
timestamp 1621523292
transform 1 0 24380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_265
timestamp 1621523292
transform 1 0 25484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_277
timestamp 1621523292
transform 1 0 26588 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1621523292
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_286
timestamp 1621523292
transform 1 0 27416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_298
timestamp 1621523292
transform 1 0 28520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_310
timestamp 1621523292
transform 1 0 29624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_322
timestamp 1621523292
transform 1 0 30728 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1621523292
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_334
timestamp 1621523292
transform 1 0 31832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1621523292
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_355
timestamp 1621523292
transform 1 0 33764 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1621523292
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1621523292
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_391
timestamp 1621523292
transform 1 0 37076 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1621523292
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_400
timestamp 1621523292
transform 1 0 37904 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_412
timestamp 1621523292
transform 1 0 39008 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_424
timestamp 1621523292
transform 1 0 40112 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_436
timestamp 1621523292
transform 1 0 41216 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1621523292
transform 1 0 43056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_448
timestamp 1621523292
transform 1 0 42320 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_457
timestamp 1621523292
transform 1 0 43148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_469
timestamp 1621523292
transform 1 0 44252 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_481
timestamp 1621523292
transform 1 0 45356 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_493
timestamp 1621523292
transform 1 0 46460 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1621523292
transform 1 0 48300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1621523292
transform 1 0 47564 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_514
timestamp 1621523292
transform 1 0 48392 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2127_
timestamp 1621523292
transform 1 0 50416 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1621523292
transform 1 0 49772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_526
timestamp 1621523292
transform 1 0 49496 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_532
timestamp 1621523292
transform 1 0 50048 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_539
timestamp 1621523292
transform 1 0 50692 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1621523292
transform 1 0 52900 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2128_
timestamp 1621523292
transform 1 0 51428 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2129_
timestamp 1621523292
transform 1 0 52256 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_550
timestamp 1621523292
transform 1 0 51704 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_559
timestamp 1621523292
transform 1 0 52532 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_566
timestamp 1621523292
transform 1 0 53176 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1607_
timestamp 1621523292
transform 1 0 54648 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1632_
timestamp 1621523292
transform 1 0 54004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1621523292
transform 1 0 53544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_571
timestamp 1621523292
transform 1 0 53636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_578
timestamp 1621523292
transform 1 0 54280 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_586
timestamp 1621523292
transform 1 0 55016 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output237
timestamp 1621523292
transform 1 0 56764 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output276
timestamp 1621523292
transform 1 0 55752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_598
timestamp 1621523292
transform 1 0 56120 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_604
timestamp 1621523292
transform 1 0 56672 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_609
timestamp 1621523292
transform 1 0 57132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2296_
timestamp 1621523292
transform 1 0 57500 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1621523292
transform -1 0 58880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1621523292
transform 1 0 58236 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1621523292
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1621523292
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output317
timestamp 1621523292
transform 1 0 1748 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1621523292
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_11
timestamp 1621523292
transform 1 0 2116 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1621523292
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1621523292
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1621523292
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_23
timestamp 1621523292
transform 1 0 3220 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1621523292
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1621523292
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1621523292
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1621523292
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1621523292
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1621523292
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1621523292
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1621523292
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1621523292
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1621523292
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1621523292
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1621523292
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1621523292
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1621523292
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1621523292
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1621523292
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1621523292
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1621523292
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1621523292
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1621523292
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1621523292
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1621523292
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1621523292
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1621523292
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1621523292
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1621523292
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1621523292
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1621523292
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1621523292
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1621523292
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1621523292
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1621523292
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1621523292
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1621523292
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1621523292
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1621523292
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1621523292
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1621523292
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1621523292
transform 1 0 20700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1621523292
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1621523292
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1621523292
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_237
timestamp 1621523292
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_220
timestamp 1621523292
transform 1 0 21344 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1621523292
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1621523292
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_249
timestamp 1621523292
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1621523292
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_241
timestamp 1621523292
transform 1 0 23276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1621523292
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_270
timestamp 1621523292
transform 1 0 25944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1621523292
transform 1 0 27048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1621523292
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1621523292
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1621523292
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_294
timestamp 1621523292
transform 1 0 28152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1621523292
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_298
timestamp 1621523292
transform 1 0 28520 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1621523292
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_306
timestamp 1621523292
transform 1 0 29256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_315
timestamp 1621523292
transform 1 0 30084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_327
timestamp 1621523292
transform 1 0 31188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_310
timestamp 1621523292
transform 1 0 29624 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_322
timestamp 1621523292
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1621523292
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_339
timestamp 1621523292
transform 1 0 32292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_334
timestamp 1621523292
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_343
timestamp 1621523292
transform 1 0 32660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1621523292
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_351
timestamp 1621523292
transform 1 0 33396 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_363
timestamp 1621523292
transform 1 0 34500 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_355
timestamp 1621523292
transform 1 0 33764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1621523292
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_372
timestamp 1621523292
transform 1 0 35328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_384
timestamp 1621523292
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1621523292
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_391
timestamp 1621523292
transform 1 0 37076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1621523292
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_396
timestamp 1621523292
transform 1 0 37536 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_408
timestamp 1621523292
transform 1 0 38640 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_400
timestamp 1621523292
transform 1 0 37904 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_412
timestamp 1621523292
transform 1 0 39008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1621523292
transform 1 0 40480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_420
timestamp 1621523292
transform 1 0 39744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_429
timestamp 1621523292
transform 1 0 40572 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_424
timestamp 1621523292
transform 1 0 40112 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_436
timestamp 1621523292
transform 1 0 41216 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1621523292
transform 1 0 43056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_441
timestamp 1621523292
transform 1 0 41676 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_453
timestamp 1621523292
transform 1 0 42780 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_448
timestamp 1621523292
transform 1 0 42320 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_457
timestamp 1621523292
transform 1 0 43148 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_465
timestamp 1621523292
transform 1 0 43884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_477
timestamp 1621523292
transform 1 0 44988 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_469
timestamp 1621523292
transform 1 0 44252 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1621523292
transform 1 0 45724 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_486
timestamp 1621523292
transform 1 0 45816 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_498
timestamp 1621523292
transform 1 0 46920 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_481
timestamp 1621523292
transform 1 0 45356 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_493
timestamp 1621523292
transform 1 0 46460 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1621523292
transform 1 0 48300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_510
timestamp 1621523292
transform 1 0 48024 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_522
timestamp 1621523292
transform 1 0 49128 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1621523292
transform 1 0 47564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_514
timestamp 1621523292
transform 1 0 48392 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1621523292
transform 1 0 50968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_534
timestamp 1621523292
transform 1 0 50232 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_543
timestamp 1621523292
transform 1 0 51060 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_526
timestamp 1621523292
transform 1 0 49496 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_538
timestamp 1621523292
transform 1 0 50600 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_546
timestamp 1621523292
transform 1 0 51336 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1621523292
transform 1 0 51612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2146_
timestamp 1621523292
transform 1 0 51612 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_552
timestamp 1621523292
transform 1 0 51888 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_552
timestamp 1621523292
transform 1 0 51888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_559
timestamp 1621523292
transform 1 0 52532 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_559
timestamp 1621523292
transform 1 0 52532 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2145_
timestamp 1621523292
transform 1 0 52256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2136_
timestamp 1621523292
transform 1 0 52256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2138_
timestamp 1621523292
transform 1 0 52900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2130_
timestamp 1621523292
transform 1 0 52900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_566
timestamp 1621523292
transform 1 0 53176 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_566
timestamp 1621523292
transform 1 0 53176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_571
timestamp 1621523292
transform 1 0 53636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1621523292
transform 1 0 53544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1621523292
transform 1 0 53544 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_573
timestamp 1621523292
transform 1 0 53820 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2131_
timestamp 1621523292
transform 1 0 54004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1631_
timestamp 1621523292
transform 1 0 54188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_582
timestamp 1621523292
transform 1 0 54648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_578
timestamp 1621523292
transform 1 0 54280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_580
timestamp 1621523292
transform 1 0 54464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_586
timestamp 1621523292
transform 1 0 55016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_587
timestamp 1621523292
transform 1 0 55108 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1636_
timestamp 1621523292
transform 1 0 54740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1630_
timestamp 1621523292
transform 1 0 54832 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_593
timestamp 1621523292
transform 1 0 55660 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_595
timestamp 1621523292
transform 1 0 55844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output279
timestamp 1621523292
transform 1 0 55476 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output247
timestamp 1621523292
transform 1 0 56028 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1585_
timestamp 1621523292
transform 1 0 55384 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_601
timestamp 1621523292
transform 1 0 56396 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_600
timestamp 1621523292
transform 1 0 56304 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1621523292
transform 1 0 56212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2259_
timestamp 1621523292
transform 1 0 56764 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2258_
timestamp 1621523292
transform 1 0 56672 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1621523292
transform -1 0 58880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1621523292
transform -1 0 58880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output208
timestamp 1621523292
transform 1 0 57868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output246
timestamp 1621523292
transform 1 0 57868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_612
timestamp 1621523292
transform 1 0 57408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_616
timestamp 1621523292
transform 1 0 57776 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1621523292
transform 1 0 58236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_613
timestamp 1621523292
transform 1 0 57500 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1621523292
transform 1 0 58236 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1621523292
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output318
timestamp 1621523292
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1621523292
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_11
timestamp 1621523292
transform 1 0 2116 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1621523292
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_23
timestamp 1621523292
transform 1 0 3220 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1621523292
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1621523292
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1621523292
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1621523292
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1621523292
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1621523292
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1621523292
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1621523292
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1621523292
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1621523292
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1621523292
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1621523292
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1621523292
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1621523292
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1621523292
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1621523292
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1621523292
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1621523292
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1621523292
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_213
timestamp 1621523292
transform 1 0 20700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_225
timestamp 1621523292
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_237
timestamp 1621523292
transform 1 0 22908 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1621523292
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1621523292
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_258
timestamp 1621523292
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_270
timestamp 1621523292
transform 1 0 25944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1621523292
transform 1 0 27048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_294
timestamp 1621523292
transform 1 0 28152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1621523292
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1621523292
transform 1 0 29256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_315
timestamp 1621523292
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_327
timestamp 1621523292
transform 1 0 31188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_339
timestamp 1621523292
transform 1 0 32292 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1621523292
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_351
timestamp 1621523292
transform 1 0 33396 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_363
timestamp 1621523292
transform 1 0 34500 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1621523292
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1621523292
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_396
timestamp 1621523292
transform 1 0 37536 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_408
timestamp 1621523292
transform 1 0 38640 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1621523292
transform 1 0 40480 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_420
timestamp 1621523292
transform 1 0 39744 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_429
timestamp 1621523292
transform 1 0 40572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_441
timestamp 1621523292
transform 1 0 41676 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_453
timestamp 1621523292
transform 1 0 42780 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_465
timestamp 1621523292
transform 1 0 43884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_477
timestamp 1621523292
transform 1 0 44988 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1621523292
transform 1 0 45724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_486
timestamp 1621523292
transform 1 0 45816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_498
timestamp 1621523292
transform 1 0 46920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_510
timestamp 1621523292
transform 1 0 48024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_522
timestamp 1621523292
transform 1 0 49128 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1621523292
transform 1 0 50968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_534
timestamp 1621523292
transform 1 0 50232 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_543
timestamp 1621523292
transform 1 0 51060 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _2140_
timestamp 1621523292
transform 1 0 52992 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2148_
timestamp 1621523292
transform 1 0 52348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1621523292
transform 1 0 51704 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_549
timestamp 1621523292
transform 1 0 51612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_553
timestamp 1621523292
transform 1 0 51980 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_560
timestamp 1621523292
transform 1 0 52624 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_567
timestamp 1621523292
transform 1 0 53268 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1713_
timestamp 1621523292
transform 1 0 54924 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2132_
timestamp 1621523292
transform 1 0 54280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2137_
timestamp 1621523292
transform 1 0 53636 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_574
timestamp 1621523292
transform 1 0 53912 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_581
timestamp 1621523292
transform 1 0 54556 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_588
timestamp 1621523292
transform 1 0 55200 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1629_
timestamp 1621523292
transform 1 0 55568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2260_
timestamp 1621523292
transform 1 0 56764 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1621523292
transform 1 0 56212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_595
timestamp 1621523292
transform 1 0 55844 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_600
timestamp 1621523292
transform 1 0 56304 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_604
timestamp 1621523292
transform 1 0 56672 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1621523292
transform -1 0 58880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output209
timestamp 1621523292
transform 1 0 57868 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_613
timestamp 1621523292
transform 1 0 57500 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_621
timestamp 1621523292
transform 1 0 58236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1621523292
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1621523292
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1621523292
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1621523292
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1621523292
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1621523292
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1621523292
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1621523292
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1621523292
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1621523292
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1621523292
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1621523292
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1621523292
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1621523292
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1621523292
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1621523292
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1621523292
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1621523292
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1621523292
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1621523292
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1621523292
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1621523292
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1621523292
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1621523292
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1621523292
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1621523292
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1621523292
transform 1 0 23276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1621523292
transform 1 0 24380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_265
timestamp 1621523292
transform 1 0 25484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_277
timestamp 1621523292
transform 1 0 26588 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1621523292
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_286
timestamp 1621523292
transform 1 0 27416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_298
timestamp 1621523292
transform 1 0 28520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_310
timestamp 1621523292
transform 1 0 29624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_322
timestamp 1621523292
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1621523292
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_334
timestamp 1621523292
transform 1 0 31832 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1621523292
transform 1 0 32660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1621523292
transform 1 0 33764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1621523292
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1621523292
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1621523292
transform 1 0 37076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1621523292
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_400
timestamp 1621523292
transform 1 0 37904 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_412
timestamp 1621523292
transform 1 0 39008 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_424
timestamp 1621523292
transform 1 0 40112 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_436
timestamp 1621523292
transform 1 0 41216 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1621523292
transform 1 0 43056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_448
timestamp 1621523292
transform 1 0 42320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_457
timestamp 1621523292
transform 1 0 43148 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_469
timestamp 1621523292
transform 1 0 44252 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_481
timestamp 1621523292
transform 1 0 45356 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_493
timestamp 1621523292
transform 1 0 46460 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1621523292
transform 1 0 48300 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1621523292
transform 1 0 47564 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_514
timestamp 1621523292
transform 1 0 48392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_526
timestamp 1621523292
transform 1 0 49496 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_538
timestamp 1621523292
transform 1 0 50600 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1621523292
transform 1 0 52900 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_550
timestamp 1621523292
transform 1 0 51704 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_562
timestamp 1621523292
transform 1 0 52808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_566
timestamp 1621523292
transform 1 0 53176 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2133_
timestamp 1621523292
transform 1 0 55108 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2135_
timestamp 1621523292
transform 1 0 54464 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1621523292
transform 1 0 53544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_571
timestamp 1621523292
transform 1 0 53636 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_579
timestamp 1621523292
transform 1 0 54372 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_583
timestamp 1621523292
transform 1 0 54740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1584_
timestamp 1621523292
transform 1 0 55752 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2298_
timestamp 1621523292
transform 1 0 56396 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_590
timestamp 1621523292
transform 1 0 55384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_597
timestamp 1621523292
transform 1 0 56028 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_609
timestamp 1621523292
transform 1 0 57132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2297_
timestamp 1621523292
transform 1 0 57500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1621523292
transform -1 0 58880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1621523292
transform 1 0 58236 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1621523292
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output319
timestamp 1621523292
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1621523292
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_11
timestamp 1621523292
transform 1 0 2116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1621523292
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_23
timestamp 1621523292
transform 1 0 3220 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1621523292
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1621523292
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1621523292
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1621523292
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1621523292
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1621523292
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1621523292
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1621523292
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1621523292
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1621523292
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1621523292
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1621523292
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1621523292
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1621523292
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1621523292
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1621523292
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1621523292
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1621523292
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1621523292
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_213
timestamp 1621523292
transform 1 0 20700 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_225
timestamp 1621523292
transform 1 0 21804 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1621523292
transform 1 0 22908 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1621523292
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_249
timestamp 1621523292
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1621523292
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_270
timestamp 1621523292
transform 1 0 25944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_282
timestamp 1621523292
transform 1 0 27048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_294
timestamp 1621523292
transform 1 0 28152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1621523292
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_306
timestamp 1621523292
transform 1 0 29256 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1621523292
transform 1 0 30084 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_327
timestamp 1621523292
transform 1 0 31188 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_339
timestamp 1621523292
transform 1 0 32292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1621523292
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_351
timestamp 1621523292
transform 1 0 33396 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_363
timestamp 1621523292
transform 1 0 34500 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1621523292
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_384
timestamp 1621523292
transform 1 0 36432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_396
timestamp 1621523292
transform 1 0 37536 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_408
timestamp 1621523292
transform 1 0 38640 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1621523292
transform 1 0 40480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_420
timestamp 1621523292
transform 1 0 39744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_429
timestamp 1621523292
transform 1 0 40572 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_441
timestamp 1621523292
transform 1 0 41676 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_453
timestamp 1621523292
transform 1 0 42780 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_465
timestamp 1621523292
transform 1 0 43884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_477
timestamp 1621523292
transform 1 0 44988 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1621523292
transform 1 0 45724 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_486
timestamp 1621523292
transform 1 0 45816 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_498
timestamp 1621523292
transform 1 0 46920 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_510
timestamp 1621523292
transform 1 0 48024 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_522
timestamp 1621523292
transform 1 0 49128 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1621523292
transform 1 0 50968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_534
timestamp 1621523292
transform 1 0 50232 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_543
timestamp 1621523292
transform 1 0 51060 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_555
timestamp 1621523292
transform 1 0 52164 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_567
timestamp 1621523292
transform 1 0 53268 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2139_
timestamp 1621523292
transform 1 0 54924 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2147_
timestamp 1621523292
transform 1 0 54280 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1621523292
transform 1 0 53636 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_574
timestamp 1621523292
transform 1 0 53912 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_581
timestamp 1621523292
transform 1 0 54556 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_588
timestamp 1621523292
transform 1 0 55200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2134_
timestamp 1621523292
transform 1 0 55568 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2261_
timestamp 1621523292
transform 1 0 57132 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1621523292
transform 1 0 56212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_595
timestamp 1621523292
transform 1 0 55844 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_600
timestamp 1621523292
transform 1 0 56304 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_608
timestamp 1621523292
transform 1 0 57040 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1621523292
transform -1 0 58880 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_617
timestamp 1621523292
transform 1 0 57868 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1621523292
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1621523292
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1621523292
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1621523292
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1621523292
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1621523292
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1621523292
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1621523292
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1621523292
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1621523292
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1621523292
transform 1 0 9752 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_106
timestamp 1621523292
transform 1 0 10856 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1621523292
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1621523292
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1621523292
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1621523292
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1621523292
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1621523292
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1621523292
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1621523292
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1621523292
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1621523292
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1621523292
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1621523292
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1621523292
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_229
timestamp 1621523292
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_241
timestamp 1621523292
transform 1 0 23276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1621523292
transform 1 0 24380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_265
timestamp 1621523292
transform 1 0 25484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_277
timestamp 1621523292
transform 1 0 26588 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1621523292
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1621523292
transform 1 0 27416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1621523292
transform 1 0 28520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1621523292
transform 1 0 29624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1621523292
transform 1 0 30728 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1621523292
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_334
timestamp 1621523292
transform 1 0 31832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_343
timestamp 1621523292
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1621523292
transform 1 0 33764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1621523292
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1621523292
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_391
timestamp 1621523292
transform 1 0 37076 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1621523292
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_400
timestamp 1621523292
transform 1 0 37904 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_412
timestamp 1621523292
transform 1 0 39008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_424
timestamp 1621523292
transform 1 0 40112 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_436
timestamp 1621523292
transform 1 0 41216 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1621523292
transform 1 0 43056 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_448
timestamp 1621523292
transform 1 0 42320 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_457
timestamp 1621523292
transform 1 0 43148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_469
timestamp 1621523292
transform 1 0 44252 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_481
timestamp 1621523292
transform 1 0 45356 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_493
timestamp 1621523292
transform 1 0 46460 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1621523292
transform 1 0 48300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1621523292
transform 1 0 47564 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_514
timestamp 1621523292
transform 1 0 48392 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_526
timestamp 1621523292
transform 1 0 49496 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_538
timestamp 1621523292
transform 1 0 50600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_550
timestamp 1621523292
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_562
timestamp 1621523292
transform 1 0 52808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1628_
timestamp 1621523292
transform 1 0 55292 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2149_
timestamp 1621523292
transform 1 0 54648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1621523292
transform 1 0 53544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_571
timestamp 1621523292
transform 1 0 53636 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_579
timestamp 1621523292
transform 1 0 54372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_585
timestamp 1621523292
transform 1 0 54924 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1626_
timestamp 1621523292
transform 1 0 55936 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output248
timestamp 1621523292
transform 1 0 57132 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_592
timestamp 1621523292
transform 1 0 55568 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_599
timestamp 1621523292
transform 1 0 56212 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_607
timestamp 1621523292
transform 1 0 56948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1621523292
transform -1 0 58880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output210
timestamp 1621523292
transform 1 0 57868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_613
timestamp 1621523292
transform 1 0 57500 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_621
timestamp 1621523292
transform 1 0 58236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1621523292
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output320
timestamp 1621523292
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1621523292
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_11
timestamp 1621523292
transform 1 0 2116 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1621523292
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_23
timestamp 1621523292
transform 1 0 3220 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1621523292
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1621523292
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1621523292
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1621523292
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1621523292
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1621523292
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1621523292
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1621523292
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1621523292
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1621523292
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1621523292
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1621523292
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1621523292
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1621523292
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1621523292
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1621523292
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1621523292
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1621523292
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1621523292
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1621523292
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_225
timestamp 1621523292
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_237
timestamp 1621523292
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1621523292
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_249
timestamp 1621523292
transform 1 0 24012 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1621523292
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1621523292
transform 1 0 25944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1621523292
transform 1 0 27048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1621523292
transform 1 0 28152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1621523292
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_306
timestamp 1621523292
transform 1 0 29256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_315
timestamp 1621523292
transform 1 0 30084 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_327
timestamp 1621523292
transform 1 0 31188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_339
timestamp 1621523292
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1621523292
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1621523292
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1621523292
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1621523292
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1621523292
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_396
timestamp 1621523292
transform 1 0 37536 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_408
timestamp 1621523292
transform 1 0 38640 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1621523292
transform 1 0 40480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_420
timestamp 1621523292
transform 1 0 39744 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_429
timestamp 1621523292
transform 1 0 40572 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_441
timestamp 1621523292
transform 1 0 41676 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_453
timestamp 1621523292
transform 1 0 42780 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_465
timestamp 1621523292
transform 1 0 43884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1621523292
transform 1 0 44988 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1621523292
transform 1 0 45724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_486
timestamp 1621523292
transform 1 0 45816 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_498
timestamp 1621523292
transform 1 0 46920 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_510
timestamp 1621523292
transform 1 0 48024 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_522
timestamp 1621523292
transform 1 0 49128 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1621523292
transform 1 0 50968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_534
timestamp 1621523292
transform 1 0 50232 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_543
timestamp 1621523292
transform 1 0 51060 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_555
timestamp 1621523292
transform 1 0 52164 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_567
timestamp 1621523292
transform 1 0 53268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2150_
timestamp 1621523292
transform 1 0 54924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_579
timestamp 1621523292
transform 1 0 54372 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_588
timestamp 1621523292
transform 1 0 55200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1627_
timestamp 1621523292
transform 1 0 56856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2142_
timestamp 1621523292
transform 1 0 55568 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1621523292
transform 1 0 56212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_595
timestamp 1621523292
transform 1 0 55844 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_600
timestamp 1621523292
transform 1 0 56304 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_609
timestamp 1621523292
transform 1 0 57132 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2299_
timestamp 1621523292
transform 1 0 57500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1621523292
transform -1 0 58880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1621523292
transform 1 0 58236 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1621523292
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1621523292
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output290
timestamp 1621523292
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1621523292
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_11
timestamp 1621523292
transform 1 0 2116 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1621523292
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1621523292
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1621523292
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_23
timestamp 1621523292
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_35
timestamp 1621523292
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1621523292
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1621523292
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1621523292
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1621523292
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1621523292
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1621523292
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1621523292
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1621523292
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1621523292
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1621523292
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1621523292
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1621523292
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1621523292
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1621523292
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1621523292
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1621523292
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1621523292
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1621523292
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1621523292
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1621523292
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1621523292
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1621523292
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1621523292
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1621523292
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1621523292
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1621523292
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1621523292
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1621523292
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1621523292
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1621523292
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1621523292
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1621523292
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1621523292
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1621523292
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1621523292
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1621523292
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1621523292
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1621523292
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1621523292
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1621523292
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1621523292
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1621523292
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1621523292
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1621523292
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1621523292
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1621523292
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1621523292
transform 1 0 23276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1621523292
transform 1 0 24380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_249
timestamp 1621523292
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1621523292
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1621523292
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1621523292
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_270
timestamp 1621523292
transform 1 0 25944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_282
timestamp 1621523292
transform 1 0 27048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1621523292
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1621523292
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_298
timestamp 1621523292
transform 1 0 28520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_294
timestamp 1621523292
transform 1 0 28152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1621523292
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_310
timestamp 1621523292
transform 1 0 29624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_322
timestamp 1621523292
transform 1 0 30728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_306
timestamp 1621523292
transform 1 0 29256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_315
timestamp 1621523292
transform 1 0 30084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_327
timestamp 1621523292
transform 1 0 31188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1621523292
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_334
timestamp 1621523292
transform 1 0 31832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1621523292
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_339
timestamp 1621523292
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1621523292
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_355
timestamp 1621523292
transform 1 0 33764 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1621523292
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1621523292
transform 1 0 33396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_363
timestamp 1621523292
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1621523292
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_391
timestamp 1621523292
transform 1 0 37076 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1621523292
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1621523292
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1621523292
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_400
timestamp 1621523292
transform 1 0 37904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_412
timestamp 1621523292
transform 1 0 39008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_396
timestamp 1621523292
transform 1 0 37536 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_408
timestamp 1621523292
transform 1 0 38640 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1621523292
transform 1 0 40480 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_424
timestamp 1621523292
transform 1 0 40112 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_436
timestamp 1621523292
transform 1 0 41216 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_420
timestamp 1621523292
transform 1 0 39744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_429
timestamp 1621523292
transform 1 0 40572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1621523292
transform 1 0 43056 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_448
timestamp 1621523292
transform 1 0 42320 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_457
timestamp 1621523292
transform 1 0 43148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_441
timestamp 1621523292
transform 1 0 41676 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_453
timestamp 1621523292
transform 1 0 42780 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_469
timestamp 1621523292
transform 1 0 44252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_465
timestamp 1621523292
transform 1 0 43884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1621523292
transform 1 0 44988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1621523292
transform 1 0 45724 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_481
timestamp 1621523292
transform 1 0 45356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_493
timestamp 1621523292
transform 1 0 46460 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_486
timestamp 1621523292
transform 1 0 45816 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_498
timestamp 1621523292
transform 1 0 46920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1621523292
transform 1 0 48300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1621523292
transform 1 0 47564 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_514
timestamp 1621523292
transform 1 0 48392 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1621523292
transform 1 0 48024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_522
timestamp 1621523292
transform 1 0 49128 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1621523292
transform 1 0 50968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_526
timestamp 1621523292
transform 1 0 49496 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_538
timestamp 1621523292
transform 1 0 50600 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_534
timestamp 1621523292
transform 1 0 50232 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_543
timestamp 1621523292
transform 1 0 51060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_550
timestamp 1621523292
transform 1 0 51704 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_562
timestamp 1621523292
transform 1 0 52808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_555
timestamp 1621523292
transform 1 0 52164 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_567
timestamp 1621523292
transform 1 0 53268 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1621523292
transform 1 0 53544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_571
timestamp 1621523292
transform 1 0 53636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_583
timestamp 1621523292
transform 1 0 54740 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_579
timestamp 1621523292
transform 1 0 54372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_595
timestamp 1621523292
transform 1 0 55844 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_591
timestamp 1621523292
transform 1 0 55476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_596
timestamp 1621523292
transform 1 0 55936 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_591
timestamp 1621523292
transform 1 0 55476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1621523292
transform 1 0 55568 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1621523292
transform 1 0 55660 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_600
timestamp 1621523292
transform 1 0 56304 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_603
timestamp 1621523292
transform 1 0 56580 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1621523292
transform 1 0 56212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2262_
timestamp 1621523292
transform 1 0 56948 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2141_
timestamp 1621523292
transform 1 0 56304 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_608
timestamp 1621523292
transform 1 0 57040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1621523292
transform 1 0 57224 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1621523292
transform -1 0 58880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1621523292
transform -1 0 58880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output249
timestamp 1621523292
transform 1 0 57868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_615
timestamp 1621523292
transform 1 0 57684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1621523292
transform 1 0 58420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1621523292
transform 1 0 57500 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1621523292
transform 1 0 58236 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1621523292
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output291
timestamp 1621523292
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1621523292
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_11
timestamp 1621523292
transform 1 0 2116 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_23
timestamp 1621523292
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_35
timestamp 1621523292
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1621523292
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1621523292
transform 1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1621523292
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1621523292
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1621523292
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1621523292
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1621523292
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1621523292
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1621523292
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1621523292
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1621523292
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1621523292
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1621523292
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1621523292
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1621523292
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1621523292
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1621523292
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1621523292
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1621523292
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1621523292
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1621523292
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1621523292
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_241
timestamp 1621523292
transform 1 0 23276 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_253
timestamp 1621523292
transform 1 0 24380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_265
timestamp 1621523292
transform 1 0 25484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_277
timestamp 1621523292
transform 1 0 26588 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1621523292
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1621523292
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_298
timestamp 1621523292
transform 1 0 28520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_310
timestamp 1621523292
transform 1 0 29624 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_322
timestamp 1621523292
transform 1 0 30728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1621523292
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_334
timestamp 1621523292
transform 1 0 31832 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1621523292
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1621523292
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1621523292
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1621523292
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1621523292
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1621523292
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_400
timestamp 1621523292
transform 1 0 37904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_412
timestamp 1621523292
transform 1 0 39008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_424
timestamp 1621523292
transform 1 0 40112 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_436
timestamp 1621523292
transform 1 0 41216 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1621523292
transform 1 0 43056 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_448
timestamp 1621523292
transform 1 0 42320 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_457
timestamp 1621523292
transform 1 0 43148 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_469
timestamp 1621523292
transform 1 0 44252 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_481
timestamp 1621523292
transform 1 0 45356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_493
timestamp 1621523292
transform 1 0 46460 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1621523292
transform 1 0 48300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1621523292
transform 1 0 47564 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_514
timestamp 1621523292
transform 1 0 48392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_526
timestamp 1621523292
transform 1 0 49496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_538
timestamp 1621523292
transform 1 0 50600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1621523292
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_562
timestamp 1621523292
transform 1 0 52808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1621523292
transform 1 0 53544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_571
timestamp 1621523292
transform 1 0 53636 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_583
timestamp 1621523292
transform 1 0 54740 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1582_
timestamp 1621523292
transform 1 0 56856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2151_
timestamp 1621523292
transform 1 0 56212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_595
timestamp 1621523292
transform 1 0 55844 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_602
timestamp 1621523292
transform 1 0 56488 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_609
timestamp 1621523292
transform 1 0 57132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2300_
timestamp 1621523292
transform 1 0 57500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1621523292
transform -1 0 58880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1621523292
transform 1 0 58236 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1621523292
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1621523292
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1621523292
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1621523292
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1621523292
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1621523292
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1621523292
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1621523292
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1621523292
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1621523292
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1621523292
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1621523292
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1621523292
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1621523292
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1621523292
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1621523292
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1621523292
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1621523292
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1621523292
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1621523292
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1621523292
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1621523292
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1621523292
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1621523292
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1621523292
transform 1 0 20700 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1621523292
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1621523292
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1621523292
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1621523292
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1621523292
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_270
timestamp 1621523292
transform 1 0 25944 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_282
timestamp 1621523292
transform 1 0 27048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_294
timestamp 1621523292
transform 1 0 28152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1621523292
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_306
timestamp 1621523292
transform 1 0 29256 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1621523292
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1621523292
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1621523292
transform 1 0 32292 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1621523292
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1621523292
transform 1 0 33396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_363
timestamp 1621523292
transform 1 0 34500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1621523292
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1621523292
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_396
timestamp 1621523292
transform 1 0 37536 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_408
timestamp 1621523292
transform 1 0 38640 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1621523292
transform 1 0 40480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_420
timestamp 1621523292
transform 1 0 39744 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_429
timestamp 1621523292
transform 1 0 40572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_441
timestamp 1621523292
transform 1 0 41676 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_453
timestamp 1621523292
transform 1 0 42780 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_465
timestamp 1621523292
transform 1 0 43884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_477
timestamp 1621523292
transform 1 0 44988 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1621523292
transform 1 0 45724 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_486
timestamp 1621523292
transform 1 0 45816 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_498
timestamp 1621523292
transform 1 0 46920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_510
timestamp 1621523292
transform 1 0 48024 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_522
timestamp 1621523292
transform 1 0 49128 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1621523292
transform 1 0 50968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_534
timestamp 1621523292
transform 1 0 50232 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_543
timestamp 1621523292
transform 1 0 51060 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_555
timestamp 1621523292
transform 1 0 52164 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_567
timestamp 1621523292
transform 1 0 53268 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_579
timestamp 1621523292
transform 1 0 54372 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1580_
timestamp 1621523292
transform 1 0 57224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1621523292
transform 1 0 56212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1621523292
transform 1 0 55568 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_591
timestamp 1621523292
transform 1 0 55476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_595
timestamp 1621523292
transform 1 0 55844 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_600
timestamp 1621523292
transform 1 0 56304 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_608
timestamp 1621523292
transform 1 0 57040 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1621523292
transform -1 0 58880 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output211
timestamp 1621523292
transform 1 0 57868 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_613
timestamp 1621523292
transform 1 0 57500 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1621523292
transform 1 0 58236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1621523292
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output292
timestamp 1621523292
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1621523292
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_11
timestamp 1621523292
transform 1 0 2116 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_23
timestamp 1621523292
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1621523292
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1621523292
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1621523292
transform 1 0 5428 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1621523292
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1621523292
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1621523292
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1621523292
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1621523292
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1621523292
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1621523292
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1621523292
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1621523292
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1621523292
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1621523292
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1621523292
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1621523292
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1621523292
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1621523292
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1621523292
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1621523292
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1621523292
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1621523292
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1621523292
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1621523292
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1621523292
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1621523292
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1621523292
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1621523292
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1621523292
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_298
timestamp 1621523292
transform 1 0 28520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_310
timestamp 1621523292
transform 1 0 29624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1621523292
transform 1 0 30728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1621523292
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1621523292
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1621523292
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1621523292
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1621523292
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1621523292
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_391
timestamp 1621523292
transform 1 0 37076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1621523292
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_400
timestamp 1621523292
transform 1 0 37904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_412
timestamp 1621523292
transform 1 0 39008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_424
timestamp 1621523292
transform 1 0 40112 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_436
timestamp 1621523292
transform 1 0 41216 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1621523292
transform 1 0 43056 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_448
timestamp 1621523292
transform 1 0 42320 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_457
timestamp 1621523292
transform 1 0 43148 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_469
timestamp 1621523292
transform 1 0 44252 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_481
timestamp 1621523292
transform 1 0 45356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_493
timestamp 1621523292
transform 1 0 46460 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1621523292
transform 1 0 48300 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1621523292
transform 1 0 47564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_514
timestamp 1621523292
transform 1 0 48392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_526
timestamp 1621523292
transform 1 0 49496 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_538
timestamp 1621523292
transform 1 0 50600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1621523292
transform 1 0 51704 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_562
timestamp 1621523292
transform 1 0 52808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1621523292
transform 1 0 53544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_571
timestamp 1621523292
transform 1 0 53636 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_583
timestamp 1621523292
transform 1 0 54740 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_589
timestamp 1621523292
transform 1 0 55292 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1625_
timestamp 1621523292
transform 1 0 56672 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2143_
timestamp 1621523292
transform 1 0 56028 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2152_
timestamp 1621523292
transform 1 0 55384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2263_
timestamp 1621523292
transform 1 0 57316 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_593
timestamp 1621523292
transform 1 0 55660 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_600
timestamp 1621523292
transform 1 0 56304 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_607
timestamp 1621523292
transform 1 0 56948 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1621523292
transform -1 0 58880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_619
timestamp 1621523292
transform 1 0 58052 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1621523292
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output293
timestamp 1621523292
transform 1 0 1748 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1621523292
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_11
timestamp 1621523292
transform 1 0 2116 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1621523292
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_23
timestamp 1621523292
transform 1 0 3220 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1621523292
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1621523292
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1621523292
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1621523292
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1621523292
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1621523292
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1621523292
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1621523292
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1621523292
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1621523292
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1621523292
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1621523292
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1621523292
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1621523292
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1621523292
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1621523292
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1621523292
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1621523292
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1621523292
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1621523292
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1621523292
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1621523292
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1621523292
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1621523292
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1621523292
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1621523292
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1621523292
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_294
timestamp 1621523292
transform 1 0 28152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1621523292
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_306
timestamp 1621523292
transform 1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1621523292
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_327
timestamp 1621523292
transform 1 0 31188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_339
timestamp 1621523292
transform 1 0 32292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1621523292
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1621523292
transform 1 0 33396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_363
timestamp 1621523292
transform 1 0 34500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1621523292
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1621523292
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_396
timestamp 1621523292
transform 1 0 37536 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_408
timestamp 1621523292
transform 1 0 38640 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1621523292
transform 1 0 40480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_420
timestamp 1621523292
transform 1 0 39744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_429
timestamp 1621523292
transform 1 0 40572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_441
timestamp 1621523292
transform 1 0 41676 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_453
timestamp 1621523292
transform 1 0 42780 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_465
timestamp 1621523292
transform 1 0 43884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1621523292
transform 1 0 44988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1621523292
transform 1 0 45724 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_486
timestamp 1621523292
transform 1 0 45816 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_498
timestamp 1621523292
transform 1 0 46920 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_510
timestamp 1621523292
transform 1 0 48024 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_522
timestamp 1621523292
transform 1 0 49128 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1621523292
transform 1 0 50968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_534
timestamp 1621523292
transform 1 0 50232 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_543
timestamp 1621523292
transform 1 0 51060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_555
timestamp 1621523292
transform 1 0 52164 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_567
timestamp 1621523292
transform 1 0 53268 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_579
timestamp 1621523292
transform 1 0 54372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1621523292
transform 1 0 56212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output250
timestamp 1621523292
transform 1 0 56764 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_591
timestamp 1621523292
transform 1 0 55476 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_600
timestamp 1621523292
transform 1 0 56304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_604
timestamp 1621523292
transform 1 0 56672 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_609
timestamp 1621523292
transform 1 0 57132 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2301_
timestamp 1621523292
transform 1 0 57500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1621523292
transform -1 0 58880 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1621523292
transform 1 0 58236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1621523292
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1621523292
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output294
timestamp 1621523292
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1621523292
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1621523292
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1621523292
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_11
timestamp 1621523292
transform 1 0 2116 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1621523292
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1621523292
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1621523292
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_23
timestamp 1621523292
transform 1 0 3220 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1621523292
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1621523292
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1621523292
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1621523292
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1621523292
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1621523292
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1621523292
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1621523292
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1621523292
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1621523292
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1621523292
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_87
timestamp 1621523292
transform 1 0 9108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_94
timestamp 1621523292
transform 1 0 9752 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_106
timestamp 1621523292
transform 1 0 10856 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1621523292
transform 1 0 10212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1621523292
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1621523292
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1621523292
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_111
timestamp 1621523292
transform 1 0 11316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1621523292
transform 1 0 12420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1621523292
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1621523292
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1621523292
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_135
timestamp 1621523292
transform 1 0 13524 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1621523292
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1621523292
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1621523292
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1621523292
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1621523292
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1621523292
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1621523292
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1621523292
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1621523292
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1621523292
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1621523292
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1621523292
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1621523292
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1621523292
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1621523292
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1621523292
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1621523292
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1621523292
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1621523292
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1621523292
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1621523292
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1621523292
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1621523292
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1621523292
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1621523292
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1621523292
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1621523292
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1621523292
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1621523292
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1621523292
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1621523292
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1621523292
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1621523292
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_310
timestamp 1621523292
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1621523292
transform 1 0 30728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_306
timestamp 1621523292
transform 1 0 29256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1621523292
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_327
timestamp 1621523292
transform 1 0 31188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1621523292
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_334
timestamp 1621523292
transform 1 0 31832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_343
timestamp 1621523292
transform 1 0 32660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1621523292
transform 1 0 32292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1621523292
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_355
timestamp 1621523292
transform 1 0 33764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1621523292
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1621523292
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1621523292
transform 1 0 34500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1621523292
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_391
timestamp 1621523292
transform 1 0 37076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1621523292
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1621523292
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1621523292
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_400
timestamp 1621523292
transform 1 0 37904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1621523292
transform 1 0 39008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_396
timestamp 1621523292
transform 1 0 37536 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1621523292
transform 1 0 38640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1621523292
transform 1 0 40480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_424
timestamp 1621523292
transform 1 0 40112 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_436
timestamp 1621523292
transform 1 0 41216 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_420
timestamp 1621523292
transform 1 0 39744 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_429
timestamp 1621523292
transform 1 0 40572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1621523292
transform 1 0 43056 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_448
timestamp 1621523292
transform 1 0 42320 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_457
timestamp 1621523292
transform 1 0 43148 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_441
timestamp 1621523292
transform 1 0 41676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_453
timestamp 1621523292
transform 1 0 42780 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_469
timestamp 1621523292
transform 1 0 44252 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_465
timestamp 1621523292
transform 1 0 43884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1621523292
transform 1 0 44988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1621523292
transform 1 0 45724 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_481
timestamp 1621523292
transform 1 0 45356 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_493
timestamp 1621523292
transform 1 0 46460 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_486
timestamp 1621523292
transform 1 0 45816 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_498
timestamp 1621523292
transform 1 0 46920 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1621523292
transform 1 0 48300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1621523292
transform 1 0 47564 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_514
timestamp 1621523292
transform 1 0 48392 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_510
timestamp 1621523292
transform 1 0 48024 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_522
timestamp 1621523292
transform 1 0 49128 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1621523292
transform 1 0 50968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_526
timestamp 1621523292
transform 1 0 49496 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_538
timestamp 1621523292
transform 1 0 50600 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_534
timestamp 1621523292
transform 1 0 50232 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_543
timestamp 1621523292
transform 1 0 51060 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_550
timestamp 1621523292
transform 1 0 51704 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_562
timestamp 1621523292
transform 1 0 52808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_555
timestamp 1621523292
transform 1 0 52164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_567
timestamp 1621523292
transform 1 0 53268 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1621523292
transform 1 0 53544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_571
timestamp 1621523292
transform 1 0 53636 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_583
timestamp 1621523292
transform 1 0 54740 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_589
timestamp 1621523292
transform 1 0 55292 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_579
timestamp 1621523292
transform 1 0 54372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_595
timestamp 1621523292
transform 1 0 55844 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_591
timestamp 1621523292
transform 1 0 55476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_593
timestamp 1621523292
transform 1 0 55660 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1621523292
transform 1 0 55384 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2153_
timestamp 1621523292
transform 1 0 55568 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1620_
timestamp 1621523292
transform 1 0 56028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_600
timestamp 1621523292
transform 1 0 56304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_600
timestamp 1621523292
transform 1 0 56304 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 56488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1621523292
transform 1 0 56212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2264_
timestamp 1621523292
transform 1 0 56672 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_608
timestamp 1621523292
transform 1 0 57040 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output251
timestamp 1621523292
transform 1 0 57132 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1621523292
transform -1 0 58880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1621523292
transform -1 0 58880 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output212
timestamp 1621523292
transform 1 0 57868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output213
timestamp 1621523292
transform 1 0 57868 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_613
timestamp 1621523292
transform 1 0 57500 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1621523292
transform 1 0 58236 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_612
timestamp 1621523292
transform 1 0 57408 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_616
timestamp 1621523292
transform 1 0 57776 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1621523292
transform 1 0 58236 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1621523292
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1621523292
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1621523292
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1621523292
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1621523292
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1621523292
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1621523292
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1621523292
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1621523292
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1621523292
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_94
timestamp 1621523292
transform 1 0 9752 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1621523292
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1621523292
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_115
timestamp 1621523292
transform 1 0 11684 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_127
timestamp 1621523292
transform 1 0 12788 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1621523292
transform 1 0 13892 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_151
timestamp 1621523292
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1621523292
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_163
timestamp 1621523292
transform 1 0 16100 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1621523292
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1621523292
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1621523292
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1621523292
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1621523292
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1621523292
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_229
timestamp 1621523292
transform 1 0 22172 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_241
timestamp 1621523292
transform 1 0 23276 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_253
timestamp 1621523292
transform 1 0 24380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_265
timestamp 1621523292
transform 1 0 25484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_277
timestamp 1621523292
transform 1 0 26588 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1621523292
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1621523292
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1621523292
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1621523292
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1621523292
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1621523292
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1621523292
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1621523292
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_355
timestamp 1621523292
transform 1 0 33764 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1621523292
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1621523292
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1621523292
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1621523292
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_400
timestamp 1621523292
transform 1 0 37904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1621523292
transform 1 0 39008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_424
timestamp 1621523292
transform 1 0 40112 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_436
timestamp 1621523292
transform 1 0 41216 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1621523292
transform 1 0 43056 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_448
timestamp 1621523292
transform 1 0 42320 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_457
timestamp 1621523292
transform 1 0 43148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_469
timestamp 1621523292
transform 1 0 44252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1621523292
transform 1 0 45356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_493
timestamp 1621523292
transform 1 0 46460 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1621523292
transform 1 0 48300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1621523292
transform 1 0 47564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_514
timestamp 1621523292
transform 1 0 48392 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_526
timestamp 1621523292
transform 1 0 49496 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_538
timestamp 1621523292
transform 1 0 50600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_550
timestamp 1621523292
transform 1 0 51704 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_562
timestamp 1621523292
transform 1 0 52808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1621523292
transform 1 0 53544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_571
timestamp 1621523292
transform 1 0 53636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_583
timestamp 1621523292
transform 1 0 54740 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1621523292
transform 1 0 56856 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1624_
timestamp 1621523292
transform 1 0 56212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2184_
timestamp 1621523292
transform 1 0 55568 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_591
timestamp 1621523292
transform 1 0 55476 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_595
timestamp 1621523292
transform 1 0 55844 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_602
timestamp 1621523292
transform 1 0 56488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_609
timestamp 1621523292
transform 1 0 57132 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2302_
timestamp 1621523292
transform 1 0 57500 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1621523292
transform -1 0 58880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_621
timestamp 1621523292
transform 1 0 58236 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1621523292
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output295
timestamp 1621523292
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1621523292
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1621523292
transform 1 0 2116 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1621523292
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1621523292
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1621523292
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1621523292
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1621523292
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1621523292
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1621523292
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1621523292
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1621523292
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1621523292
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1621523292
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1621523292
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1621523292
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1621523292
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_144
timestamp 1621523292
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1621523292
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1621523292
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1621523292
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_192
timestamp 1621523292
transform 1 0 18768 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1621523292
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1621523292
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1621523292
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_225
timestamp 1621523292
transform 1 0 21804 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_237
timestamp 1621523292
transform 1 0 22908 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1621523292
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_249
timestamp 1621523292
transform 1 0 24012 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1621523292
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1621523292
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1621523292
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1621523292
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1621523292
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1621523292
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_315
timestamp 1621523292
transform 1 0 30084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_327
timestamp 1621523292
transform 1 0 31188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1621523292
transform 1 0 32292 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1621523292
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1621523292
transform 1 0 33396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1621523292
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1621523292
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_384
timestamp 1621523292
transform 1 0 36432 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_396
timestamp 1621523292
transform 1 0 37536 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_408
timestamp 1621523292
transform 1 0 38640 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1621523292
transform 1 0 40480 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_420
timestamp 1621523292
transform 1 0 39744 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_429
timestamp 1621523292
transform 1 0 40572 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_441
timestamp 1621523292
transform 1 0 41676 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_453
timestamp 1621523292
transform 1 0 42780 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_465
timestamp 1621523292
transform 1 0 43884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_477
timestamp 1621523292
transform 1 0 44988 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1621523292
transform 1 0 45724 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_486
timestamp 1621523292
transform 1 0 45816 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1621523292
transform 1 0 46920 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_510
timestamp 1621523292
transform 1 0 48024 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_522
timestamp 1621523292
transform 1 0 49128 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1621523292
transform 1 0 50968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_534
timestamp 1621523292
transform 1 0 50232 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_543
timestamp 1621523292
transform 1 0 51060 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_555
timestamp 1621523292
transform 1 0 52164 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_567
timestamp 1621523292
transform 1 0 53268 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_579
timestamp 1621523292
transform 1 0 54372 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1541_
timestamp 1621523292
transform 1 0 56764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1621523292
transform 1 0 56212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1621523292
transform 1 0 55568 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_591
timestamp 1621523292
transform 1 0 55476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_595
timestamp 1621523292
transform 1 0 55844 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_600
timestamp 1621523292
transform 1 0 56304 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_604
timestamp 1621523292
transform 1 0 56672 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_608
timestamp 1621523292
transform 1 0 57040 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2333_
timestamp 1621523292
transform 1 0 57408 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1621523292
transform -1 0 58880 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1621523292
transform 1 0 58236 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1621523292
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output296
timestamp 1621523292
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1621523292
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_11
timestamp 1621523292
transform 1 0 2116 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_23
timestamp 1621523292
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_35
timestamp 1621523292
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1621523292
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1621523292
transform 1 0 5428 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1621523292
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1621523292
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1621523292
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1621523292
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1621523292
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1621523292
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1621523292
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1621523292
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1621523292
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1621523292
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1621523292
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1621523292
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1621523292
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1621523292
transform 1 0 16928 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1621523292
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1621523292
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1621523292
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1621523292
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_220
timestamp 1621523292
transform 1 0 21344 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1621523292
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1621523292
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1621523292
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1621523292
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1621523292
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1621523292
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1621523292
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1621523292
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1621523292
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1621523292
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1621523292
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1621523292
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1621523292
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1621523292
transform 1 0 33764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1621523292
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1621523292
transform 1 0 35972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_391
timestamp 1621523292
transform 1 0 37076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1621523292
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1621523292
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1621523292
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_424
timestamp 1621523292
transform 1 0 40112 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_436
timestamp 1621523292
transform 1 0 41216 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1621523292
transform 1 0 43056 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_448
timestamp 1621523292
transform 1 0 42320 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_457
timestamp 1621523292
transform 1 0 43148 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_469
timestamp 1621523292
transform 1 0 44252 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_481
timestamp 1621523292
transform 1 0 45356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_493
timestamp 1621523292
transform 1 0 46460 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1621523292
transform 1 0 48300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1621523292
transform 1 0 47564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_514
timestamp 1621523292
transform 1 0 48392 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_526
timestamp 1621523292
transform 1 0 49496 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_538
timestamp 1621523292
transform 1 0 50600 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_550
timestamp 1621523292
transform 1 0 51704 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_562
timestamp 1621523292
transform 1 0 52808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1621523292
transform 1 0 53544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_571
timestamp 1621523292
transform 1 0 53636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_583
timestamp 1621523292
transform 1 0 54740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1623_
timestamp 1621523292
transform 1 0 55936 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2265_
timestamp 1621523292
transform 1 0 56580 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1621523292
transform 1 0 56396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_595
timestamp 1621523292
transform 1 0 55844 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_599
timestamp 1621523292
transform 1 0 56212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_611
timestamp 1621523292
transform 1 0 57316 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1621523292
transform -1 0 58880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output216
timestamp 1621523292
transform 1 0 57868 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1621523292
transform 1 0 58236 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1621523292
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1621523292
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1621523292
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1621523292
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1621523292
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1621523292
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1621523292
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1621523292
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1621523292
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1621523292
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1621523292
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1621523292
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1621523292
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1621523292
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1621523292
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1621523292
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1621523292
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1621523292
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1621523292
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_168
timestamp 1621523292
transform 1 0 16560 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_180
timestamp 1621523292
transform 1 0 17664 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_192
timestamp 1621523292
transform 1 0 18768 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1621523292
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1621523292
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_213
timestamp 1621523292
transform 1 0 20700 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_225
timestamp 1621523292
transform 1 0 21804 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_237
timestamp 1621523292
transform 1 0 22908 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1621523292
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_249
timestamp 1621523292
transform 1 0 24012 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1621523292
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_270
timestamp 1621523292
transform 1 0 25944 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_282
timestamp 1621523292
transform 1 0 27048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_294
timestamp 1621523292
transform 1 0 28152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1621523292
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1621523292
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1621523292
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1621523292
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_339
timestamp 1621523292
transform 1 0 32292 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1621523292
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_351
timestamp 1621523292
transform 1 0 33396 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_363
timestamp 1621523292
transform 1 0 34500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_372
timestamp 1621523292
transform 1 0 35328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_384
timestamp 1621523292
transform 1 0 36432 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_396
timestamp 1621523292
transform 1 0 37536 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_408
timestamp 1621523292
transform 1 0 38640 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1621523292
transform 1 0 40480 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_420
timestamp 1621523292
transform 1 0 39744 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_429
timestamp 1621523292
transform 1 0 40572 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_441
timestamp 1621523292
transform 1 0 41676 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_453
timestamp 1621523292
transform 1 0 42780 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_465
timestamp 1621523292
transform 1 0 43884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_477
timestamp 1621523292
transform 1 0 44988 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1621523292
transform 1 0 45724 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_486
timestamp 1621523292
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_498
timestamp 1621523292
transform 1 0 46920 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_510
timestamp 1621523292
transform 1 0 48024 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_522
timestamp 1621523292
transform 1 0 49128 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1621523292
transform 1 0 50968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_534
timestamp 1621523292
transform 1 0 50232 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_543
timestamp 1621523292
transform 1 0 51060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_555
timestamp 1621523292
transform 1 0 52164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_567
timestamp 1621523292
transform 1 0 53268 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2154_
timestamp 1621523292
transform 1 0 54924 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_579
timestamp 1621523292
transform 1 0 54372 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_588
timestamp 1621523292
transform 1 0 55200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1578_
timestamp 1621523292
transform 1 0 55568 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1621523292
transform 1 0 56212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output252
timestamp 1621523292
transform 1 0 56764 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_595
timestamp 1621523292
transform 1 0 55844 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_600
timestamp 1621523292
transform 1 0 56304 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_604
timestamp 1621523292
transform 1 0 56672 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_609
timestamp 1621523292
transform 1 0 57132 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2303_
timestamp 1621523292
transform 1 0 57500 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1621523292
transform -1 0 58880 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_621
timestamp 1621523292
transform 1 0 58236 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1621523292
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output297
timestamp 1621523292
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1621523292
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_11
timestamp 1621523292
transform 1 0 2116 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_23
timestamp 1621523292
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_35
timestamp 1621523292
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1621523292
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1621523292
transform 1 0 5428 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1621523292
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1621523292
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_70
timestamp 1621523292
transform 1 0 7544 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_82
timestamp 1621523292
transform 1 0 8648 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_94
timestamp 1621523292
transform 1 0 9752 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_106
timestamp 1621523292
transform 1 0 10856 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1621523292
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1621523292
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1621523292
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _1539_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 14720 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_139
timestamp 1621523292
transform 1 0 13892 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_147
timestamp 1621523292
transform 1 0 14628 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1621523292
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_154
timestamp 1621523292
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_166
timestamp 1621523292
transform 1 0 16376 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_170
timestamp 1621523292
transform 1 0 16744 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1621523292
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1621523292
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1621523292
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1621523292
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1621523292
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_220
timestamp 1621523292
transform 1 0 21344 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_229
timestamp 1621523292
transform 1 0 22172 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_241
timestamp 1621523292
transform 1 0 23276 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1621523292
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1621523292
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_277
timestamp 1621523292
transform 1 0 26588 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1621523292
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1621523292
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_298
timestamp 1621523292
transform 1 0 28520 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_310
timestamp 1621523292
transform 1 0 29624 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1621523292
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1621523292
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_334
timestamp 1621523292
transform 1 0 31832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1621523292
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1621523292
transform 1 0 33764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1621523292
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1621523292
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_391
timestamp 1621523292
transform 1 0 37076 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1621523292
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_400
timestamp 1621523292
transform 1 0 37904 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_412
timestamp 1621523292
transform 1 0 39008 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_424
timestamp 1621523292
transform 1 0 40112 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_436
timestamp 1621523292
transform 1 0 41216 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1621523292
transform 1 0 43056 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_448
timestamp 1621523292
transform 1 0 42320 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_457
timestamp 1621523292
transform 1 0 43148 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_469
timestamp 1621523292
transform 1 0 44252 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_481
timestamp 1621523292
transform 1 0 45356 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_493
timestamp 1621523292
transform 1 0 46460 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1621523292
transform 1 0 48300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_505
timestamp 1621523292
transform 1 0 47564 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_514
timestamp 1621523292
transform 1 0 48392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_526
timestamp 1621523292
transform 1 0 49496 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_538
timestamp 1621523292
transform 1 0 50600 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1621523292
transform 1 0 51704 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_562
timestamp 1621523292
transform 1 0 52808 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1621523292
transform 1 0 53544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1621523292
transform 1 0 54832 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_571
timestamp 1621523292
transform 1 0 53636 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_583
timestamp 1621523292
transform 1 0 54740 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_587
timestamp 1621523292
transform 1 0 55108 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1540_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 56764 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1577_
timestamp 1621523292
transform 1 0 56120 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2155_
timestamp 1621523292
transform 1 0 55476 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_594
timestamp 1621523292
transform 1 0 55752 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_601
timestamp 1621523292
transform 1 0 56396 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_611
timestamp 1621523292
transform 1 0 57316 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1621523292
transform -1 0 58880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output214
timestamp 1621523292
transform 1 0 57868 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1621523292
transform 1 0 58236 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1621523292
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1621523292
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output298
timestamp 1621523292
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1621523292
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1621523292
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1621523292
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1621523292
transform 1 0 2116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1621523292
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1621523292
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1621523292
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1621523292
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1621523292
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1621523292
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1621523292
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1621523292
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1621523292
transform 1 0 5428 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_55
timestamp 1621523292
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1621523292
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1621523292
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1621523292
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1621523292
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1621523292
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_70
timestamp 1621523292
transform 1 0 7544 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_82
timestamp 1621523292
transform 1 0 8648 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1703_
timestamp 1621523292
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1621523292
transform 1 0 9568 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2197_
timestamp 1621523292
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1621523292
transform 1 0 10212 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_106
timestamp 1621523292
transform 1 0 10856 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1621523292
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1621523292
transform 1 0 9844 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_108
timestamp 1621523292
transform 1 0 11040 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_4  _2196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 12052 0 1 16864
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1621523292
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_118
timestamp 1621523292
transform 1 0 11960 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_130
timestamp 1621523292
transform 1 0 13064 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_115
timestamp 1621523292
transform 1 0 11684 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1700_
timestamp 1621523292
transform 1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1702_
timestamp 1621523292
transform 1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2200_
timestamp 1621523292
transform 1 0 13616 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1621523292
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_139
timestamp 1621523292
transform 1 0 13892 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1621523292
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_132
timestamp 1621523292
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_145
timestamp 1621523292
transform 1 0 14444 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_152
timestamp 1621523292
transform 1 0 15088 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1621523292
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1621523292
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1621523292
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_164
timestamp 1621523292
transform 1 0 16192 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_170
timestamp 1621523292
transform 1 0 16744 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1621523292
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1621523292
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1621523292
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1621523292
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1621523292
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1621523292
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_201
timestamp 1621523292
transform 1 0 19596 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_213
timestamp 1621523292
transform 1 0 20700 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_208
timestamp 1621523292
transform 1 0 20240 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_216
timestamp 1621523292
transform 1 0 20976 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 21252 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1720_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 22724 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _1722_
timestamp 1621523292
transform 1 0 22816 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1621523292
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_225
timestamp 1621523292
transform 1 0 21804 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_233
timestamp 1621523292
transform 1 0 22540 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_222
timestamp 1621523292
transform 1 0 21528 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_229
timestamp 1621523292
transform 1 0 22172 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1525_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 24012 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1621523292
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1621523292
transform 1 0 24104 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_245
timestamp 1621523292
transform 1 0 23644 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_252
timestamp 1621523292
transform 1 0 24288 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_256
timestamp 1621523292
transform 1 0 24656 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_258
timestamp 1621523292
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_244
timestamp 1621523292
transform 1 0 23552 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_258
timestamp 1621523292
transform 1 0 24840 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_270
timestamp 1621523292
transform 1 0 25944 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_282
timestamp 1621523292
transform 1 0 27048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_270
timestamp 1621523292
transform 1 0 25944 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_282
timestamp 1621523292
transform 1 0 27048 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1621523292
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_294
timestamp 1621523292
transform 1 0 28152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1621523292
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1621523292
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1621523292
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_306
timestamp 1621523292
transform 1 0 29256 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1621523292
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1621523292
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1621523292
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1621523292
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1621523292
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1621523292
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1621523292
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1621523292
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1621523292
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1621523292
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1621523292
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1621523292
transform 1 0 33764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1621523292
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1621523292
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_384
timestamp 1621523292
transform 1 0 36432 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1621523292
transform 1 0 35972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_391
timestamp 1621523292
transform 1 0 37076 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1621523292
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_396
timestamp 1621523292
transform 1 0 37536 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_408
timestamp 1621523292
transform 1 0 38640 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1621523292
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1621523292
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1621523292
transform 1 0 40480 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_420
timestamp 1621523292
transform 1 0 39744 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_429
timestamp 1621523292
transform 1 0 40572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1621523292
transform 1 0 40112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1621523292
transform 1 0 41216 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1621523292
transform 1 0 43056 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_441
timestamp 1621523292
transform 1 0 41676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_453
timestamp 1621523292
transform 1 0 42780 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_448
timestamp 1621523292
transform 1 0 42320 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_457
timestamp 1621523292
transform 1 0 43148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_465
timestamp 1621523292
transform 1 0 43884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_477
timestamp 1621523292
transform 1 0 44988 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_469
timestamp 1621523292
transform 1 0 44252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1621523292
transform 1 0 45724 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_486
timestamp 1621523292
transform 1 0 45816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_498
timestamp 1621523292
transform 1 0 46920 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_481
timestamp 1621523292
transform 1 0 45356 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_493
timestamp 1621523292
transform 1 0 46460 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1621523292
transform 1 0 48300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_510
timestamp 1621523292
transform 1 0 48024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_522
timestamp 1621523292
transform 1 0 49128 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1621523292
transform 1 0 47564 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_514
timestamp 1621523292
transform 1 0 48392 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1621523292
transform 1 0 50968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_534
timestamp 1621523292
transform 1 0 50232 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_543
timestamp 1621523292
transform 1 0 51060 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_526
timestamp 1621523292
transform 1 0 49496 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_538
timestamp 1621523292
transform 1 0 50600 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_555
timestamp 1621523292
transform 1 0 52164 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_567
timestamp 1621523292
transform 1 0 53268 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_550
timestamp 1621523292
transform 1 0 51704 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_562
timestamp 1621523292
transform 1 0 52808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1621523292
transform 1 0 53544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_579
timestamp 1621523292
transform 1 0 54372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_571
timestamp 1621523292
transform 1 0 53636 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_583
timestamp 1621523292
transform 1 0 54740 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_589
timestamp 1621523292
transform 1 0 55292 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_593
timestamp 1621523292
transform 1 0 55660 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_595
timestamp 1621523292
transform 1 0 55844 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_591
timestamp 1621523292
transform 1 0 55476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1622_
timestamp 1621523292
transform 1 0 55568 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1621_
timestamp 1621523292
transform 1 0 55384 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1576_
timestamp 1621523292
transform 1 0 56028 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_605
timestamp 1621523292
transform 1 0 56764 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_601
timestamp 1621523292
transform 1 0 56396 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_604
timestamp 1621523292
transform 1 0 56672 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_600
timestamp 1621523292
transform 1 0 56304 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1621523292
transform 1 0 56212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2266_
timestamp 1621523292
transform 1 0 56764 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1575_
timestamp 1621523292
transform 1 0 56856 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_609
timestamp 1621523292
transform 1 0 57132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2304_
timestamp 1621523292
transform 1 0 57500 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1621523292
transform -1 0 58880 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1621523292
transform -1 0 58880 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output178
timestamp 1621523292
transform 1 0 57868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_613
timestamp 1621523292
transform 1 0 57500 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1621523292
transform 1 0 58236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1621523292
transform 1 0 58236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1621523292
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output299
timestamp 1621523292
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1621523292
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_11
timestamp 1621523292
transform 1 0 2116 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1621523292
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1621523292
transform 1 0 3220 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1621523292
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1621523292
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1621523292
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1621523292
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1621523292
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1621523292
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1621523292
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_2  _2198_
timestamp 1621523292
transform 1 0 10396 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_99
timestamp 1621523292
transform 1 0 10212 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1705_
timestamp 1621523292
transform 1 0 12052 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_110
timestamp 1621523292
transform 1 0 11224 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_118
timestamp 1621523292
transform 1 0 11960 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_122
timestamp 1621523292
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1621523292
transform 1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1770_
timestamp 1621523292
transform 1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1621523292
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1621523292
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_139
timestamp 1621523292
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1621523292
transform 1 0 14352 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_151
timestamp 1621523292
transform 1 0 14996 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 15364 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 16008 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_158
timestamp 1621523292
transform 1 0 15640 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1621523292
transform 1 0 16284 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1621523292
transform 1 0 17388 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_189
timestamp 1621523292
transform 1 0 18492 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2455_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 19964 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1621523292
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_197
timestamp 1621523292
transform 1 0 19228 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_201
timestamp 1621523292
transform 1 0 19596 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1621523292
transform 1 0 21804 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1721_
timestamp 1621523292
transform 1 0 22816 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1621523292
transform 1 0 21436 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_228
timestamp 1621523292
transform 1 0 22080 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1621523292
transform 1 0 24012 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1325_
timestamp 1621523292
transform 1 0 25208 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1621523292
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_245
timestamp 1621523292
transform 1 0 23644 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_252
timestamp 1621523292
transform 1 0 24288 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_256
timestamp 1621523292
transform 1 0 24656 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_258
timestamp 1621523292
transform 1 0 24840 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2523_
timestamp 1621523292
transform 1 0 25852 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_28_265
timestamp 1621523292
transform 1 0 25484 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_285
timestamp 1621523292
transform 1 0 27324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_297
timestamp 1621523292
transform 1 0 28428 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1621523292
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1621523292
transform 1 0 29532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_313
timestamp 1621523292
transform 1 0 29900 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1621523292
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1621523292
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1621523292
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1621523292
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1621523292
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1621523292
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1621523292
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1621523292
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_396
timestamp 1621523292
transform 1 0 37536 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_408
timestamp 1621523292
transform 1 0 38640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1621523292
transform 1 0 40480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_420
timestamp 1621523292
transform 1 0 39744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_429
timestamp 1621523292
transform 1 0 40572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_441
timestamp 1621523292
transform 1 0 41676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_453
timestamp 1621523292
transform 1 0 42780 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_465
timestamp 1621523292
transform 1 0 43884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 1621523292
transform 1 0 44988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1621523292
transform 1 0 45724 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_486
timestamp 1621523292
transform 1 0 45816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_498
timestamp 1621523292
transform 1 0 46920 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_510
timestamp 1621523292
transform 1 0 48024 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_522
timestamp 1621523292
transform 1 0 49128 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1621523292
transform 1 0 50968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_534
timestamp 1621523292
transform 1 0 50232 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_543
timestamp 1621523292
transform 1 0 51060 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_555
timestamp 1621523292
transform 1 0 52164 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_567
timestamp 1621523292
transform 1 0 53268 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_579
timestamp 1621523292
transform 1 0 54372 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_1  _2267_
timestamp 1621523292
transform 1 0 56672 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1621523292
transform 1 0 56212 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1621523292
transform 1 0 56488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_591
timestamp 1621523292
transform 1 0 55476 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_600
timestamp 1621523292
transform 1 0 56304 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1621523292
transform -1 0 58880 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output217
timestamp 1621523292
transform 1 0 57868 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_612
timestamp 1621523292
transform 1 0 57408 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_616
timestamp 1621523292
transform 1 0 57776 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_621
timestamp 1621523292
transform 1 0 58236 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1621523292
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1621523292
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1621523292
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1621523292
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_39
timestamp 1621523292
transform 1 0 4692 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1777_
timestamp 1621523292
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1621523292
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_47
timestamp 1621523292
transform 1 0 5428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_53
timestamp 1621523292
transform 1 0 5980 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1621523292
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_4  _2194_
timestamp 1621523292
transform 1 0 8280 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_29_70
timestamp 1621523292
transform 1 0 7544 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 10764 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1763_
timestamp 1621523292
transform 1 0 9936 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1621523292
transform 1 0 9476 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_95
timestamp 1621523292
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_101
timestamp 1621523292
transform 1 0 10396 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1765_
timestamp 1621523292
transform 1 0 12972 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2099_
timestamp 1621523292
transform 1 0 12328 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1621523292
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_110
timestamp 1621523292
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_115
timestamp 1621523292
transform 1 0 11684 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1621523292
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1621523292
transform 1 0 12604 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_4  _2199_
timestamp 1621523292
transform 1 0 13616 0 1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1621523292
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1621523292
transform 1 0 14812 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1766_
timestamp 1621523292
transform 1 0 15180 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1769_
timestamp 1621523292
transform 1 0 16100 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1621523292
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_156
timestamp 1621523292
transform 1 0 15456 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1621523292
transform 1 0 16008 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_166
timestamp 1621523292
transform 1 0 16376 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_170
timestamp 1621523292
transform 1 0 16744 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1621523292
transform 1 0 16928 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1452_
timestamp 1621523292
transform 1 0 18308 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1527_
timestamp 1621523292
transform 1 0 18952 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2101_
timestamp 1621523292
transform 1 0 17296 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_179
timestamp 1621523292
transform 1 0 17572 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_190
timestamp 1621523292
transform 1 0 18584 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1165_
timestamp 1621523292
transform 1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _1166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 20976 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1526_
timestamp 1621523292
transform 1 0 19688 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_197
timestamp 1621523292
transform 1 0 19228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_201
timestamp 1621523292
transform 1 0 19596 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_205
timestamp 1621523292
transform 1 0 19964 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_212
timestamp 1621523292
transform 1 0 20608 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1723_
timestamp 1621523292
transform 1 0 22724 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1621523292
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_223
timestamp 1621523292
transform 1 0 21620 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_227
timestamp 1621523292
transform 1 0 21988 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_229
timestamp 1621523292
transform 1 0 22172 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2456_
timestamp 1621523292
transform 1 0 23920 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1621523292
transform 1 0 23552 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1523_
timestamp 1621523292
transform 1 0 26036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_264
timestamp 1621523292
transform 1 0 25392 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_270
timestamp 1621523292
transform 1 0 25944 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_274
timestamp 1621523292
transform 1 0 26312 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_282
timestamp 1621523292
transform 1 0 27048 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1328_
timestamp 1621523292
transform 1 0 27784 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 1621523292
transform 1 0 28428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1621523292
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_286
timestamp 1621523292
transform 1 0 27416 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1621523292
transform 1 0 28060 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_300
timestamp 1621523292
transform 1 0 28704 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1522_
timestamp 1621523292
transform 1 0 29256 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_309
timestamp 1621523292
transform 1 0 29532 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_321
timestamp 1621523292
transform 1 0 30636 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1621523292
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_333
timestamp 1621523292
transform 1 0 31740 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_341
timestamp 1621523292
transform 1 0 32476 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1621523292
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_355
timestamp 1621523292
transform 1 0 33764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1621523292
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1621523292
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_391
timestamp 1621523292
transform 1 0 37076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1621523292
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1621523292
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_412
timestamp 1621523292
transform 1 0 39008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1621523292
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1621523292
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1621523292
transform 1 0 43056 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_448
timestamp 1621523292
transform 1 0 42320 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_457
timestamp 1621523292
transform 1 0 43148 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_469
timestamp 1621523292
transform 1 0 44252 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_481
timestamp 1621523292
transform 1 0 45356 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_493
timestamp 1621523292
transform 1 0 46460 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1621523292
transform 1 0 48300 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1621523292
transform 1 0 47564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_514
timestamp 1621523292
transform 1 0 48392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_526
timestamp 1621523292
transform 1 0 49496 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_538
timestamp 1621523292
transform 1 0 50600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_550
timestamp 1621523292
transform 1 0 51704 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_562
timestamp 1621523292
transform 1 0 52808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1621523292
transform 1 0 53544 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_571
timestamp 1621523292
transform 1 0 53636 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_583
timestamp 1621523292
transform 1 0 54740 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1621523292
transform 1 0 56856 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1621523292
transform 1 0 56212 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_595
timestamp 1621523292
transform 1 0 55844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_602
timestamp 1621523292
transform 1 0 56488 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_609
timestamp 1621523292
transform 1 0 57132 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2305_
timestamp 1621523292
transform 1 0 57500 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1621523292
transform -1 0 58880 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_621
timestamp 1621523292
transform 1 0 58236 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1697_
timestamp 1621523292
transform 1 0 2852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1621523292
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output301
timestamp 1621523292
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1621523292
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_11
timestamp 1621523292
transform 1 0 2116 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1621523292
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1621523292
transform 1 0 3128 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1621523292
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1621523292
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_42
timestamp 1621523292
transform 1 0 4968 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1771_
timestamp 1621523292
transform 1 0 5612 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1772_
timestamp 1621523292
transform 1 0 6256 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1780_
timestamp 1621523292
transform 1 0 6900 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_48
timestamp 1621523292
transform 1 0 5520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1621523292
transform 1 0 5888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1621523292
transform 1 0 6532 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1708_
timestamp 1621523292
transform 1 0 8188 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1709_
timestamp 1621523292
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1621523292
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_66
timestamp 1621523292
transform 1 0 7176 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1621523292
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_80
timestamp 1621523292
transform 1 0 8464 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_87
timestamp 1621523292
transform 1 0 9108 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1758_
timestamp 1621523292
transform 1 0 9844 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2489_
timestamp 1621523292
transform 1 0 11132 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_100
timestamp 1621523292
transform 1 0 10304 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_108
timestamp 1621523292
transform 1 0 11040 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1762_
timestamp 1621523292
transform 1 0 12972 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1621523292
transform 1 0 12604 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1761_
timestamp 1621523292
transform 1 0 13616 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2492_
timestamp 1621523292
transform 1 0 14720 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1621523292
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1621523292
transform 1 0 13248 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_139
timestamp 1621523292
transform 1 0 13892 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_144
timestamp 1621523292
transform 1 0 14352 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1465_
timestamp 1621523292
transform 1 0 16560 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1621523292
transform 1 0 16192 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_171
timestamp 1621523292
transform 1 0 16836 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2454_
timestamp 1621523292
transform 1 0 17664 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 1621523292
transform 1 0 17572 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_196
timestamp 1621523292
transform 1 0 19136 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1621523292
transform 1 0 19964 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1182_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 20608 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1621523292
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1621523292
transform 1 0 19596 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1621523292
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2521_
timestamp 1621523292
transform 1 0 21988 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_30_220
timestamp 1621523292
transform 1 0 21344 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1621523292
transform 1 0 21896 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1621523292
transform 1 0 24012 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1621523292
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_243
timestamp 1621523292
transform 1 0 23460 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_252
timestamp 1621523292
transform 1 0 24288 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_256
timestamp 1621523292
transform 1 0 24656 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_258
timestamp 1621523292
transform 1 0 24840 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 26588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 25484 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_264
timestamp 1621523292
transform 1 0 25392 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1621523292
transform 1 0 26220 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_281
timestamp 1621523292
transform 1 0 26956 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2457_
timestamp 1621523292
transform 1 0 27508 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_30_303
timestamp 1621523292
transform 1 0 28980 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1518_
timestamp 1621523292
transform 1 0 29348 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1521_
timestamp 1621523292
transform 1 0 30912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1621523292
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_310
timestamp 1621523292
transform 1 0 29624 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_315
timestamp 1621523292
transform 1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_323
timestamp 1621523292
transform 1 0 30820 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1621523292
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1621523292
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1621523292
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1621523292
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1621523292
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1621523292
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1621523292
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1621523292
transform 1 0 37536 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1621523292
transform 1 0 38640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1621523292
transform 1 0 40480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_420
timestamp 1621523292
transform 1 0 39744 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_429
timestamp 1621523292
transform 1 0 40572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_441
timestamp 1621523292
transform 1 0 41676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_453
timestamp 1621523292
transform 1 0 42780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_465
timestamp 1621523292
transform 1 0 43884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1621523292
transform 1 0 44988 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1621523292
transform 1 0 45724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_486
timestamp 1621523292
transform 1 0 45816 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_498
timestamp 1621523292
transform 1 0 46920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_510
timestamp 1621523292
transform 1 0 48024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_522
timestamp 1621523292
transform 1 0 49128 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1621523292
transform 1 0 50968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_534
timestamp 1621523292
transform 1 0 50232 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_543
timestamp 1621523292
transform 1 0 51060 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_555
timestamp 1621523292
transform 1 0 52164 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_567
timestamp 1621523292
transform 1 0 53268 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_579
timestamp 1621523292
transform 1 0 54372 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2156_
timestamp 1621523292
transform 1 0 57224 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1621523292
transform 1 0 56212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1621523292
transform 1 0 55568 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_591
timestamp 1621523292
transform 1 0 55476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_595
timestamp 1621523292
transform 1 0 55844 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_600
timestamp 1621523292
transform 1 0 56304 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_608
timestamp 1621523292
transform 1 0 57040 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1621523292
transform -1 0 58880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output179
timestamp 1621523292
transform 1 0 57868 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1621523292
transform 1 0 57500 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1621523292
transform 1 0 58236 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1694_
timestamp 1621523292
transform 1 0 2576 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1699_
timestamp 1621523292
transform 1 0 1932 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1621523292
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1621523292
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_12
timestamp 1621523292
transform 1 0 2208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_19
timestamp 1621523292
transform 1 0 2852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1696_
timestamp 1621523292
transform 1 0 3588 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1778_
timestamp 1621523292
transform 1 0 4508 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_30
timestamp 1621523292
transform 1 0 3864 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_36
timestamp 1621523292
transform 1 0 4416 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_40
timestamp 1621523292
transform 1 0 4784 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1690_
timestamp 1621523292
transform 1 0 5152 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1621523292
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1621523292
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1621523292
transform 1 0 5428 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1621523292
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_58
timestamp 1621523292
transform 1 0 6440 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_65
timestamp 1621523292
transform 1 0 7084 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_4  _2193_
timestamp 1621523292
transform 1 0 7820 0 1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_31_86
timestamp 1621523292
transform 1 0 9016 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1759_
timestamp 1621523292
transform 1 0 9752 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1764_
timestamp 1621523292
transform 1 0 10580 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1621523292
transform 1 0 10212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_108
timestamp 1621523292
transform 1 0 11040 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2490_
timestamp 1621523292
transform 1 0 12144 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1621523292
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_115
timestamp 1621523292
transform 1 0 11684 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_119
timestamp 1621523292
transform 1 0 12052 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 15088 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1475_
timestamp 1621523292
transform 1 0 13984 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_136
timestamp 1621523292
transform 1 0 13616 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_144
timestamp 1621523292
transform 1 0 14352 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1621523292
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1621523292
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1621523292
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_166
timestamp 1621523292
transform 1 0 16376 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_170
timestamp 1621523292
transform 1 0 16744 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_172
timestamp 1621523292
transform 1 0 16928 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1170_
timestamp 1621523292
transform 1 0 19044 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 1621523292
transform 1 0 18400 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1453_
timestamp 1621523292
transform 1 0 17296 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_183
timestamp 1621523292
transform 1 0 17940 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_187
timestamp 1621523292
transform 1 0 18308 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1621523292
transform 1 0 18676 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1621523292
transform 1 0 21160 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1621523292
transform 1 0 20056 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1621523292
transform 1 0 19688 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_209
timestamp 1621523292
transform 1 0 20332 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_217
timestamp 1621523292
transform 1 0 21068 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1724_
timestamp 1621523292
transform 1 0 23000 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1621523292
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_221
timestamp 1621523292
transform 1 0 21436 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_227
timestamp 1621523292
transform 1 0 21988 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_229
timestamp 1621523292
transform 1 0 22172 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1621523292
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1163_
timestamp 1621523292
transform 1 0 24196 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_247
timestamp 1621523292
transform 1 0 23828 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_258
timestamp 1621523292
transform 1 0 24840 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 25576 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1621523292
transform 1 0 26588 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_273
timestamp 1621523292
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_280
timestamp 1621523292
transform 1 0 26864 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1621523292
transform 1 0 27784 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1621523292
transform 1 0 28612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1621523292
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_284
timestamp 1621523292
transform 1 0 27232 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_286
timestamp 1621523292
transform 1 0 27416 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1621523292
transform 1 0 28060 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_302
timestamp 1621523292
transform 1 0 28888 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1311_
timestamp 1621523292
transform 1 0 30636 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1621523292
transform 1 0 29256 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1511_
timestamp 1621523292
transform 1 0 29900 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_309
timestamp 1621523292
transform 1 0 29532 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1621523292
transform 1 0 30176 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_320
timestamp 1621523292
transform 1 0 30544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_324
timestamp 1621523292
transform 1 0 30912 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1621523292
transform 1 0 31464 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1621523292
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_333
timestamp 1621523292
transform 1 0 31740 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_341
timestamp 1621523292
transform 1 0 32476 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_343
timestamp 1621523292
transform 1 0 32660 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_355
timestamp 1621523292
transform 1 0 33764 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1621523292
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1621523292
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_391
timestamp 1621523292
transform 1 0 37076 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1621523292
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1621523292
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1621523292
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1621523292
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1621523292
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1621523292
transform 1 0 43056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_448
timestamp 1621523292
transform 1 0 42320 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_457
timestamp 1621523292
transform 1 0 43148 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_469
timestamp 1621523292
transform 1 0 44252 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_481
timestamp 1621523292
transform 1 0 45356 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_493
timestamp 1621523292
transform 1 0 46460 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1621523292
transform 1 0 48300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1621523292
transform 1 0 47564 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_514
timestamp 1621523292
transform 1 0 48392 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_526
timestamp 1621523292
transform 1 0 49496 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_538
timestamp 1621523292
transform 1 0 50600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_550
timestamp 1621523292
transform 1 0 51704 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_562
timestamp 1621523292
transform 1 0 52808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1621523292
transform 1 0 53544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_571
timestamp 1621523292
transform 1 0 53636 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_583
timestamp 1621523292
transform 1 0 54740 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1573_
timestamp 1621523292
transform 1 0 57224 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1619_
timestamp 1621523292
transform 1 0 55936 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2157_
timestamp 1621523292
transform 1 0 56580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_595
timestamp 1621523292
transform 1 0 55844 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_599
timestamp 1621523292
transform 1 0 56212 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_606
timestamp 1621523292
transform 1 0 56856 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1621523292
transform -1 0 58880 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output218
timestamp 1621523292
transform 1 0 57868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_613
timestamp 1621523292
transform 1 0 57500 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_621
timestamp 1621523292
transform 1 0 58236 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2201_
timestamp 1621523292
transform 1 0 2300 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1621523292
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output302
timestamp 1621523292
transform 1 0 1564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1621523292
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1621523292
transform 1 0 1932 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2204_
timestamp 1621523292
transform 1 0 4232 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1621523292
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_22
timestamp 1621523292
transform 1 0 3128 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_28
timestamp 1621523292
transform 1 0 3680 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_30
timestamp 1621523292
transform 1 0 3864 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_43
timestamp 1621523292
transform 1 0 5060 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2206_
timestamp 1621523292
transform 1 0 7084 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_1  _2209_
timestamp 1621523292
transform 1 0 5428 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_55
timestamp 1621523292
transform 1 0 6164 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1621523292
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1693_
timestamp 1621523292
transform 1 0 8280 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1621523292
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_74
timestamp 1621523292
transform 1 0 7912 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_81
timestamp 1621523292
transform 1 0 8556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1621523292
transform 1 0 8924 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_87
timestamp 1621523292
transform 1 0 9108 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2493_
timestamp 1621523292
transform 1 0 9476 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_32_107
timestamp 1621523292
transform 1 0 10948 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1474_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 11592 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1476_
timestamp 1621523292
transform 1 0 12788 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_113
timestamp 1621523292
transform 1 0 11500 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1621523292
transform 1 0 12420 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1467_
timestamp 1621523292
transform 1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1621523292
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_136
timestamp 1621523292
transform 1 0 13616 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_142
timestamp 1621523292
transform 1 0 14168 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1621523292
transform 1 0 14352 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_148
timestamp 1621523292
transform 1 0 14720 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_152
timestamp 1621523292
transform 1 0 15088 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1454_
timestamp 1621523292
transform 1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2496_
timestamp 1621523292
transform 1 0 16376 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_158
timestamp 1621523292
transform 1 0 15640 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_162
timestamp 1621523292
transform 1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1621523292
transform 1 0 18860 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1621523292
transform 1 0 18216 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_182
timestamp 1621523292
transform 1 0 17848 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_189
timestamp 1621523292
transform 1 0 18492 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_196
timestamp 1621523292
transform 1 0 19136 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _1183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 20424 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1621523292
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_201
timestamp 1621523292
transform 1 0 19596 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1621523292
transform 1 0 20332 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_218
timestamp 1621523292
transform 1 0 21160 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1333_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 21528 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1334_
timestamp 1621523292
transform 1 0 22632 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_230
timestamp 1621523292
transform 1 0 22264 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1324_
timestamp 1621523292
transform 1 0 23736 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1326_
timestamp 1621523292
transform 1 0 25208 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1621523292
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_242
timestamp 1621523292
transform 1 0 23368 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1621523292
transform 1 0 24380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_258
timestamp 1621523292
transform 1 0 24840 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1159_
timestamp 1621523292
transform 1 0 26588 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_32_270
timestamp 1621523292
transform 1 0 25944 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1621523292
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1621523292
transform 1 0 27600 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1306_
timestamp 1621523292
transform 1 0 28244 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1621523292
transform 1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1621523292
transform 1 0 27232 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_291
timestamp 1621523292
transform 1 0 27876 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_298
timestamp 1621523292
transform 1 0 28520 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_305
timestamp 1621523292
transform 1 0 29164 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2460_
timestamp 1621523292
transform 1 0 30912 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1621523292
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_313
timestamp 1621523292
transform 1 0 29900 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_315
timestamp 1621523292
transform 1 0 30084 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_323
timestamp 1621523292
transform 1 0 30820 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1621523292
transform 1 0 32752 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_340
timestamp 1621523292
transform 1 0 32384 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_347
timestamp 1621523292
transform 1 0 33028 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1621523292
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_359
timestamp 1621523292
transform 1 0 34132 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_372
timestamp 1621523292
transform 1 0 35328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_384
timestamp 1621523292
transform 1 0 36432 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_396
timestamp 1621523292
transform 1 0 37536 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_408
timestamp 1621523292
transform 1 0 38640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1621523292
transform 1 0 40480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_420
timestamp 1621523292
transform 1 0 39744 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_429
timestamp 1621523292
transform 1 0 40572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_441
timestamp 1621523292
transform 1 0 41676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_453
timestamp 1621523292
transform 1 0 42780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1621523292
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_477
timestamp 1621523292
transform 1 0 44988 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1621523292
transform 1 0 45724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_486
timestamp 1621523292
transform 1 0 45816 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_498
timestamp 1621523292
transform 1 0 46920 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_510
timestamp 1621523292
transform 1 0 48024 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_522
timestamp 1621523292
transform 1 0 49128 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1621523292
transform 1 0 50968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_534
timestamp 1621523292
transform 1 0 50232 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_543
timestamp 1621523292
transform 1 0 51060 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_555
timestamp 1621523292
transform 1 0 52164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_567
timestamp 1621523292
transform 1 0 53268 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1538_
timestamp 1621523292
transform 1 0 54832 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1706_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 53636 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_32_580
timestamp 1621523292
transform 1 0 54464 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2268_
timestamp 1621523292
transform 1 0 56672 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1621523292
transform 1 0 56212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_590
timestamp 1621523292
transform 1 0 55384 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_598
timestamp 1621523292
transform 1 0 56120 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_600
timestamp 1621523292
transform 1 0 56304 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1621523292
transform -1 0 58880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output180
timestamp 1621523292
transform 1 0 57868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_612
timestamp 1621523292
transform 1 0 57408 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_616
timestamp 1621523292
transform 1 0 57776 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1621523292
transform 1 0 58236 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1621523292
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_3
timestamp 1621523292
transform 1 0 1380 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output303
timestamp 1621523292
transform 1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1621523292
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1621523292
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1686_
timestamp 1621523292
transform 1 0 1932 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1621523292
transform 1 0 2760 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1621523292
transform 1 0 2116 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_18
timestamp 1621523292
transform 1 0 2760 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_12
timestamp 1621523292
transform 1 0 2208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_2  _2203_
timestamp 1621523292
transform 1 0 2852 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1682_
timestamp 1621523292
transform 1 0 2484 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_30
timestamp 1621523292
transform 1 0 3864 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_25
timestamp 1621523292
transform 1 0 3404 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_28
timestamp 1621523292
transform 1 0 3680 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1621523292
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1683_
timestamp 1621523292
transform 1 0 3128 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_37
timestamp 1621523292
transform 1 0 4508 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_39
timestamp 1621523292
transform 1 0 4692 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1621523292
transform 1 0 4416 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1684_
timestamp 1621523292
transform 1 0 4232 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2210_
timestamp 1621523292
transform 1 0 5060 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1621523292
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_51
timestamp 1621523292
transform 1 0 5796 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_44
timestamp 1621523292
transform 1 0 5152 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_51
timestamp 1621523292
transform 1 0 5796 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1688_
timestamp 1621523292
transform 1 0 5520 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_58
timestamp 1621523292
transform 1 0 6440 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_58
timestamp 1621523292
transform 1 0 6440 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1621523292
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_2  _2207_
timestamp 1621523292
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1698_
timestamp 1621523292
transform 1 0 6164 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2208_
timestamp 1621523292
transform 1 0 6992 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_71
timestamp 1621523292
transform 1 0 7636 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_73
timestamp 1621523292
transform 1 0 7820 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_78
timestamp 1621523292
transform 1 0 8280 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1776_
timestamp 1621523292
transform 1 0 8188 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1691_
timestamp 1621523292
transform 1 0 8004 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_82
timestamp 1621523292
transform 1 0 8648 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_85
timestamp 1621523292
transform 1 0 8924 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1621523292
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1775_
timestamp 1621523292
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_87
timestamp 1621523292
transform 1 0 9108 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1464_
timestamp 1621523292
transform 1 0 10120 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1756_
timestamp 1621523292
transform 1 0 9476 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2494_
timestamp 1621523292
transform 1 0 9476 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1621523292
transform 1 0 9752 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_107
timestamp 1621523292
transform 1 0 10948 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_107
timestamp 1621523292
transform 1 0 10948 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_113
timestamp 1621523292
transform 1 0 11500 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1621523292
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1621523292
transform 1 0 11500 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1621523292
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1459_
timestamp 1621523292
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_130
timestamp 1621523292
transform 1 0 13064 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_130
timestamp 1621523292
transform 1 0 13064 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_122
timestamp 1621523292
transform 1 0 12328 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1463_
timestamp 1621523292
transform 1 0 13156 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2488_
timestamp 1621523292
transform 1 0 11592 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_34_139
timestamp 1621523292
transform 1 0 13892 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1621523292
transform 1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1528_
timestamp 1621523292
transform 1 0 13616 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1472_
timestamp 1621523292
transform 1 0 13892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_144
timestamp 1621523292
transform 1 0 14352 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_152
timestamp 1621523292
transform 1 0 15088 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_143
timestamp 1621523292
transform 1 0 14260 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1621523292
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1457_
timestamp 1621523292
transform 1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2495_
timestamp 1621523292
transform 1 0 14720 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  _1442_
timestamp 1621523292
transform 1 0 16928 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1621523292
transform 1 0 16192 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1455_
timestamp 1621523292
transform 1 0 15548 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1621523292
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_156
timestamp 1621523292
transform 1 0 15456 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_160
timestamp 1621523292
transform 1 0 15824 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_167
timestamp 1621523292
transform 1 0 16468 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_172
timestamp 1621523292
transform 1 0 16928 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_164
timestamp 1621523292
transform 1 0 16192 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1621523292
transform 1 0 18860 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1340_
timestamp 1621523292
transform 1 0 17756 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2520_
timestamp 1621523292
transform 1 0 17664 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1621523292
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_176
timestamp 1621523292
transform 1 0 17296 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_180
timestamp 1621523292
transform 1 0 17664 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_184
timestamp 1621523292
transform 1 0 18032 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_192
timestamp 1621523292
transform 1 0 18768 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_196
timestamp 1621523292
transform 1 0 19136 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1178_
timestamp 1621523292
transform 1 0 19964 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1331_
timestamp 1621523292
transform 1 0 20700 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1336_
timestamp 1621523292
transform 1 0 19504 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2452_
timestamp 1621523292
transform 1 0 20700 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1621523292
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_209
timestamp 1621523292
transform 1 0 20332 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1621523292
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1621523292
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1329_
timestamp 1621523292
transform 1 0 23000 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2522_
timestamp 1621523292
transform 1 0 22540 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1621523292
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1621523292
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_229
timestamp 1621523292
transform 1 0 22172 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1621523292
transform 1 0 22908 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_229
timestamp 1621523292
transform 1 0 22172 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _1184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 25208 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _1314_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 24196 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1621523292
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_245
timestamp 1621523292
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_258
timestamp 1621523292
transform 1 0 24840 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_249
timestamp 1621523292
transform 1 0 24012 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1621523292
transform 1 0 24840 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_262
timestamp 1621523292
transform 1 0 25208 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1621523292
transform 1 0 25300 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 26404 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 26128 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_271
timestamp 1621523292
transform 1 0 26036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_280
timestamp 1621523292
transform 1 0 26864 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_266
timestamp 1621523292
transform 1 0 25576 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_281
timestamp 1621523292
transform 1 0 26956 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1621523292
transform 1 0 27324 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1621523292
transform 1 0 28152 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1313_
timestamp 1621523292
transform 1 0 28796 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2459_
timestamp 1621523292
transform 1 0 27784 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1621523292
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_284
timestamp 1621523292
transform 1 0 27232 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_286
timestamp 1621523292
transform 1 0 27416 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_288
timestamp 1621523292
transform 1 0 27600 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_297
timestamp 1621523292
transform 1 0 28428 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1307_
timestamp 1621523292
transform 1 0 31004 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2526_
timestamp 1621523292
transform 1 0 29624 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1621523292
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1621523292
transform 1 0 29256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_326
timestamp 1621523292
transform 1 0 31096 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_310
timestamp 1621523292
transform 1 0 29624 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_315
timestamp 1621523292
transform 1 0 30084 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_323
timestamp 1621523292
transform 1 0 30820 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_332
timestamp 1621523292
transform 1 0 31648 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1621523292
transform 1 0 32108 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1134_
timestamp 1621523292
transform 1 0 31464 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_34_349
timestamp 1621523292
transform 1 0 33212 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_340
timestamp 1621523292
transform 1 0 32384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_343
timestamp 1621523292
transform 1 0 32660 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_341
timestamp 1621523292
transform 1 0 32476 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1621523292
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _1188_
timestamp 1621523292
transform 1 0 32568 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2527_
timestamp 1621523292
transform 1 0 33028 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__o21ai_1  _1189_
timestamp 1621523292
transform 1 0 33580 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1621523292
transform 1 0 34316 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1519_
timestamp 1621523292
transform 1 0 34868 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1621523292
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_363
timestamp 1621523292
transform 1 0 34500 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_370
timestamp 1621523292
transform 1 0 35144 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_357
timestamp 1621523292
transform 1 0 33948 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_364
timestamp 1621523292
transform 1 0 34592 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_370
timestamp 1621523292
transform 1 0 35144 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1725_
timestamp 1621523292
transform 1 0 36892 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1726_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 36064 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1729_
timestamp 1621523292
transform 1 0 36064 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_33_378
timestamp 1621523292
transform 1 0 35880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_385
timestamp 1621523292
transform 1 0 36524 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_372
timestamp 1621523292
transform 1 0 35328 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_385
timestamp 1621523292
transform 1 0 36524 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_393
timestamp 1621523292
transform 1 0 37260 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1621523292
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_397
timestamp 1621523292
transform 1 0 37628 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_400
timestamp 1621523292
transform 1 0 37904 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_412
timestamp 1621523292
transform 1 0 39008 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_405
timestamp 1621523292
transform 1 0 38364 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1621523292
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_424
timestamp 1621523292
transform 1 0 40112 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_436
timestamp 1621523292
transform 1 0 41216 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_417
timestamp 1621523292
transform 1 0 39468 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_425
timestamp 1621523292
transform 1 0 40204 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1621523292
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1621523292
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_448
timestamp 1621523292
transform 1 0 42320 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1621523292
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1621523292
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1621523292
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1621523292
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_465
timestamp 1621523292
transform 1 0 43884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1621523292
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1621523292
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1621523292
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_493
timestamp 1621523292
transform 1 0 46460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1621523292
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_498
timestamp 1621523292
transform 1 0 46920 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1621523292
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1621523292
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_514
timestamp 1621523292
transform 1 0 48392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_510
timestamp 1621523292
transform 1 0 48024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_522
timestamp 1621523292
transform 1 0 49128 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1621523292
transform 1 0 50968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_526
timestamp 1621523292
transform 1 0 49496 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_538
timestamp 1621523292
transform 1 0 50600 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_534
timestamp 1621523292
transform 1 0 50232 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_543
timestamp 1621523292
transform 1 0 51060 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_550
timestamp 1621523292
transform 1 0 51704 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_562
timestamp 1621523292
transform 1 0 52808 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_555
timestamp 1621523292
transform 1 0 52164 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_567
timestamp 1621523292
transform 1 0 53268 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1618_
timestamp 1621523292
transform 1 0 55016 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2158_
timestamp 1621523292
transform 1 0 54924 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1621523292
transform 1 0 53544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1621523292
transform 1 0 54372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_571
timestamp 1621523292
transform 1 0 53636 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_582
timestamp 1621523292
transform 1 0 54648 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_589
timestamp 1621523292
transform 1 0 55292 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_579
timestamp 1621523292
transform 1 0 54372 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_588
timestamp 1621523292
transform 1 0 55200 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_595
timestamp 1621523292
transform 1 0 55844 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_596
timestamp 1621523292
transform 1 0 55936 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1614_
timestamp 1621523292
transform 1 0 55660 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1621523292
transform 1 0 55568 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_600
timestamp 1621523292
transform 1 0 56304 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1621523292
transform 1 0 56488 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1621523292
transform 1 0 56212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__ebufn_1  _2269_
timestamp 1621523292
transform 1 0 56672 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1545_
timestamp 1621523292
transform 1 0 56672 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_608
timestamp 1621523292
transform 1 0 57040 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2306_
timestamp 1621523292
transform 1 0 57500 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1621523292
transform -1 0 58880 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1621523292
transform -1 0 58880 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output219
timestamp 1621523292
transform 1 0 57868 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_612
timestamp 1621523292
transform 1 0 57408 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_621
timestamp 1621523292
transform 1 0 58236 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_612
timestamp 1621523292
transform 1 0 57408 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_616
timestamp 1621523292
transform 1 0 57776 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_621
timestamp 1621523292
transform 1 0 58236 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1680_
timestamp 1621523292
transform 1 0 2484 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1621523292
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output304
timestamp 1621523292
transform 1 0 1748 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1621523292
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_11
timestamp 1621523292
transform 1 0 2116 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_18
timestamp 1621523292
transform 1 0 2760 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1669_
timestamp 1621523292
transform 1 0 4784 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2202_
timestamp 1621523292
transform 1 0 3312 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_35_33
timestamp 1621523292
transform 1 0 4140 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_39
timestamp 1621523292
transform 1 0 4692 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_43
timestamp 1621523292
transform 1 0 5060 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1687_
timestamp 1621523292
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1621523292
transform 1 0 6808 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1621523292
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1621523292
transform 1 0 5704 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_56
timestamp 1621523292
transform 1 0 6256 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1621523292
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_65
timestamp 1621523292
transform 1 0 7084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1768_
timestamp 1621523292
transform 1 0 7544 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2497_
timestamp 1621523292
transform 1 0 8556 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_69
timestamp 1621523292
transform 1 0 7452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_75
timestamp 1621523292
transform 1 0 8004 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1461_
timestamp 1621523292
transform 1 0 10396 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1621523292
transform 1 0 10028 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1479_
timestamp 1621523292
transform 1 0 12052 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1621523292
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_110
timestamp 1621523292
transform 1 0 11224 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1621523292
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_128
timestamp 1621523292
transform 1 0 12880 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1449_
timestamp 1621523292
transform 1 0 14628 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1478_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 13248 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_138
timestamp 1621523292
transform 1 0 13800 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_146
timestamp 1621523292
transform 1 0 14536 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1621523292
transform 1 0 14904 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1456_
timestamp 1621523292
transform 1 0 15272 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1621523292
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_161
timestamp 1621523292
transform 1 0 15916 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1621523292
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_172
timestamp 1621523292
transform 1 0 16928 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2453_
timestamp 1621523292
transform 1 0 17756 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_180
timestamp 1621523292
transform 1 0 17664 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1621523292
transform 1 0 20792 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1335_
timestamp 1621523292
transform 1 0 19596 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_197
timestamp 1621523292
transform 1 0 19228 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_208
timestamp 1621523292
transform 1 0 20240 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_217
timestamp 1621523292
transform 1 0 21068 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1621523292
transform 1 0 21436 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1330_
timestamp 1621523292
transform 1 0 22908 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1621523292
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_224
timestamp 1621523292
transform 1 0 21712 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_229
timestamp 1621523292
transform 1 0 22172 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1153_
timestamp 1621523292
transform 1 0 25116 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1316_
timestamp 1621523292
transform 1 0 24104 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_246
timestamp 1621523292
transform 1 0 23736 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_254
timestamp 1621523292
transform 1 0 24472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_260
timestamp 1621523292
transform 1 0 25024 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_1  _1149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 26312 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_35_266
timestamp 1621523292
transform 1 0 25576 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1621523292
transform 1 0 26956 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1621523292
transform 1 0 29072 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1150_
timestamp 1621523292
transform 1 0 27784 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1621523292
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1621523292
transform 1 0 27416 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_297
timestamp 1621523292
transform 1 0 28428 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_303
timestamp 1621523292
transform 1 0 28980 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1621523292
transform 1 0 29716 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1312_
timestamp 1621523292
transform 1 0 30360 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_35_307
timestamp 1621523292
transform 1 0 29348 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_314
timestamp 1621523292
transform 1 0 29992 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_325
timestamp 1621523292
transform 1 0 31004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1130_
timestamp 1621523292
transform 1 0 33120 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1276_
timestamp 1621523292
transform 1 0 31372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1621523292
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_333
timestamp 1621523292
transform 1 0 31740 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_341
timestamp 1621523292
transform 1 0 32476 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_343
timestamp 1621523292
transform 1 0 32660 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_347
timestamp 1621523292
transform 1 0 33028 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2461_
timestamp 1621523292
transform 1 0 34132 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_35_355
timestamp 1621523292
transform 1 0 33764 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1728_
timestamp 1621523292
transform 1 0 36064 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_35_375
timestamp 1621523292
transform 1 0 35604 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_379
timestamp 1621523292
transform 1 0 35972 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_385
timestamp 1621523292
transform 1 0 36524 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1621523292
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_397
timestamp 1621523292
transform 1 0 37628 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_400
timestamp 1621523292
transform 1 0 37904 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_412
timestamp 1621523292
transform 1 0 39008 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_424
timestamp 1621523292
transform 1 0 40112 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_436
timestamp 1621523292
transform 1 0 41216 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1621523292
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_448
timestamp 1621523292
transform 1 0 42320 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_457
timestamp 1621523292
transform 1 0 43148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_469
timestamp 1621523292
transform 1 0 44252 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1621523292
transform 1 0 45356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_493
timestamp 1621523292
transform 1 0 46460 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1621523292
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1621523292
transform 1 0 47564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_514
timestamp 1621523292
transform 1 0 48392 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_526
timestamp 1621523292
transform 1 0 49496 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_538
timestamp 1621523292
transform 1 0 50600 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_550
timestamp 1621523292
transform 1 0 51704 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_562
timestamp 1621523292
transform 1 0 52808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1571_
timestamp 1621523292
transform 1 0 55016 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1621523292
transform 1 0 53544 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_571
timestamp 1621523292
transform 1 0 53636 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_583
timestamp 1621523292
transform 1 0 54740 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_589
timestamp 1621523292
transform 1 0 55292 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1570_
timestamp 1621523292
transform 1 0 56856 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2272_
timestamp 1621523292
transform 1 0 55660 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_601
timestamp 1621523292
transform 1 0 56396 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_605
timestamp 1621523292
transform 1 0 56764 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_609
timestamp 1621523292
transform 1 0 57132 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2307_
timestamp 1621523292
transform 1 0 57500 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1621523292
transform -1 0 58880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1621523292
transform 1 0 58236 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1681_
timestamp 1621523292
transform 1 0 3036 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2211_
timestamp 1621523292
transform 1 0 1932 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1621523292
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1621523292
transform 1 0 1380 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_17
timestamp 1621523292
transform 1 0 2668 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2205_
timestamp 1621523292
transform 1 0 4232 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1621523292
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1621523292
transform 1 0 3312 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_28
timestamp 1621523292
transform 1 0 3680 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_30
timestamp 1621523292
transform 1 0 3864 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_43
timestamp 1621523292
transform 1 0 5060 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _1537_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 5428 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1779_
timestamp 1621523292
transform 1 0 6624 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_36_54
timestamp 1621523292
transform 1 0 6072 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_65
timestamp 1621523292
transform 1 0 7084 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1767_
timestamp 1621523292
transform 1 0 8280 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1773_
timestamp 1621523292
transform 1 0 7452 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1621523292
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_74
timestamp 1621523292
transform 1 0 7912 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_81
timestamp 1621523292
transform 1 0 8556 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1621523292
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_87
timestamp 1621523292
transform 1 0 9108 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1415_
timestamp 1621523292
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1451_
timestamp 1621523292
transform 1 0 9936 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_36_95
timestamp 1621523292
transform 1 0 9844 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_105
timestamp 1621523292
transform 1 0 10764 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1621523292
transform 1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1458_
timestamp 1621523292
transform 1 0 11868 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1621523292
transform 1 0 11500 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_121
timestamp 1621523292
transform 1 0 12236 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1621523292
transform 1 0 12880 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1370_
timestamp 1621523292
transform 1 0 13248 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1621523292
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1621523292
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_136
timestamp 1621523292
transform 1 0 13616 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_142
timestamp 1621523292
transform 1 0 14168 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_144
timestamp 1621523292
transform 1 0 14352 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1621523292
transform 1 0 15088 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1446_
timestamp 1621523292
transform 1 0 15456 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2498_
timestamp 1621523292
transform 1 0 16100 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1621523292
transform 1 0 15732 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1448_
timestamp 1621523292
transform 1 0 17940 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1621523292
transform 1 0 17572 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_190
timestamp 1621523292
transform 1 0 18584 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1177_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 20056 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1273_
timestamp 1621523292
transform 1 0 20884 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1621523292
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_198
timestamp 1621523292
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_201
timestamp 1621523292
transform 1 0 19596 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_205
timestamp 1621523292
transform 1 0 19964 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1621523292
transform 1 0 20516 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1621523292
transform 1 0 21620 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1719_
timestamp 1621523292
transform 1 0 22540 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_219
timestamp 1621523292
transform 1 0 21252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_226
timestamp 1621523292
transform 1 0 21896 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_232
timestamp 1621523292
transform 1 0 22448 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_239
timestamp 1621523292
transform 1 0 23092 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1315_
timestamp 1621523292
transform 1 0 23920 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1520_
timestamp 1621523292
transform 1 0 25208 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1621523292
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_247
timestamp 1621523292
transform 1 0 23828 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1621523292
transform 1 0 24380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_258
timestamp 1621523292
transform 1 0 24840 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2525_
timestamp 1621523292
transform 1 0 26220 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_36_266
timestamp 1621523292
transform 1 0 25576 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_272
timestamp 1621523292
transform 1 0 26128 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2462_
timestamp 1621523292
transform 1 0 28152 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_36_289
timestamp 1621523292
transform 1 0 27692 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_293
timestamp 1621523292
transform 1 0 28060 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o31a_1  _1297_
timestamp 1621523292
transform 1 0 30728 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1621523292
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_310
timestamp 1621523292
transform 1 0 29624 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_315
timestamp 1621523292
transform 1 0 30084 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_321
timestamp 1621523292
transform 1 0 30636 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1309_
timestamp 1621523292
transform 1 0 32016 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1310_
timestamp 1621523292
transform 1 0 33120 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_329
timestamp 1621523292
transform 1 0 31372 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_335
timestamp 1621523292
transform 1 0 31924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_344
timestamp 1621523292
transform 1 0 32752 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1621523292
transform 1 0 34224 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1621523292
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_356
timestamp 1621523292
transform 1 0 33856 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1621523292
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1727_
timestamp 1621523292
transform 1 0 36064 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1730_
timestamp 1621523292
transform 1 0 36892 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_36_372
timestamp 1621523292
transform 1 0 35328 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_385
timestamp 1621523292
transform 1 0 36524 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_394
timestamp 1621523292
transform 1 0 37352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_406
timestamp 1621523292
transform 1 0 38456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1621523292
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_418
timestamp 1621523292
transform 1 0 39560 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_426
timestamp 1621523292
transform 1 0 40296 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1621523292
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1621523292
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_453
timestamp 1621523292
transform 1 0 42780 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_465
timestamp 1621523292
transform 1 0 43884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1621523292
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1621523292
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1621523292
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1621523292
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_510
timestamp 1621523292
transform 1 0 48024 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_522
timestamp 1621523292
transform 1 0 49128 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1621523292
transform 1 0 50968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_534
timestamp 1621523292
transform 1 0 50232 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_543
timestamp 1621523292
transform 1 0 51060 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_555
timestamp 1621523292
transform 1 0 52164 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_567
timestamp 1621523292
transform 1 0 53268 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1616_
timestamp 1621523292
transform 1 0 54924 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_579
timestamp 1621523292
transform 1 0 54372 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_588
timestamp 1621523292
transform 1 0 55200 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1615_
timestamp 1621523292
transform 1 0 55568 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2271_
timestamp 1621523292
transform 1 0 56672 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1621523292
transform 1 0 56212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_595
timestamp 1621523292
transform 1 0 55844 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_600
timestamp 1621523292
transform 1 0 56304 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1621523292
transform -1 0 58880 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output181
timestamp 1621523292
transform 1 0 57868 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_612
timestamp 1621523292
transform 1 0 57408 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_616
timestamp 1621523292
transform 1 0 57776 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_621
timestamp 1621523292
transform 1 0 58236 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2212_
timestamp 1621523292
transform 1 0 1748 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1621523292
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1621523292
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_15
timestamp 1621523292
transform 1 0 2484 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1670_
timestamp 1621523292
transform 1 0 4508 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _2215_
timestamp 1621523292
transform 1 0 3312 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_23
timestamp 1621523292
transform 1 0 3220 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_32
timestamp 1621523292
transform 1 0 4048 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_36
timestamp 1621523292
transform 1 0 4416 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_43
timestamp 1621523292
transform 1 0 5060 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1438_
timestamp 1621523292
transform 1 0 5704 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1621523292
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_49
timestamp 1621523292
transform 1 0 5612 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_53
timestamp 1621523292
transform 1 0 5980 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_58
timestamp 1621523292
transform 1 0 6440 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1774_
timestamp 1621523292
transform 1 0 7360 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2502_
timestamp 1621523292
transform 1 0 8464 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_37_66
timestamp 1621523292
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_73
timestamp 1621523292
transform 1 0 7820 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_79
timestamp 1621523292
transform 1 0 8372 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1435_
timestamp 1621523292
transform 1 0 10304 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_37_96
timestamp 1621523292
transform 1 0 9936 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_109
timestamp 1621523292
transform 1 0 11132 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2501_
timestamp 1621523292
transform 1 0 12052 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1621523292
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1621523292
transform 1 0 11500 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_115
timestamp 1621523292
transform 1 0 11684 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1450_
timestamp 1621523292
transform 1 0 13892 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1460_
timestamp 1621523292
transform 1 0 14628 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_135
timestamp 1621523292
transform 1 0 13524 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_143
timestamp 1621523292
transform 1 0 14260 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_151
timestamp 1621523292
transform 1 0 14996 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1621523292
transform 1 0 16192 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1443_
timestamp 1621523292
transform 1 0 15548 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1621523292
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_160
timestamp 1621523292
transform 1 0 15824 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_167
timestamp 1621523292
transform 1 0 16468 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_172
timestamp 1621523292
transform 1 0 16928 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1621523292
transform 1 0 17572 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1176_
timestamp 1621523292
transform 1 0 18952 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1621523292
transform 1 0 18216 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_178
timestamp 1621523292
transform 1 0 17480 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_182
timestamp 1621523292
transform 1 0 17848 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_190
timestamp 1621523292
transform 1 0 18584 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 19964 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1344_
timestamp 1621523292
transform 1 0 20976 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_201
timestamp 1621523292
transform 1 0 19596 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_211
timestamp 1621523292
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_215
timestamp 1621523292
transform 1 0 20884 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1264_
timestamp 1621523292
transform 1 0 22540 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1621523292
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_224
timestamp 1621523292
transform 1 0 21712 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_229
timestamp 1621523292
transform 1 0 22172 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1621523292
transform 1 0 22908 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1318_
timestamp 1621523292
transform 1 0 24564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1321_
timestamp 1621523292
transform 1 0 23736 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1621523292
transform 1 0 23644 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1621523292
transform 1 0 24196 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1319_
timestamp 1621523292
transform 1 0 25668 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_263
timestamp 1621523292
transform 1 0 25300 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_275
timestamp 1621523292
transform 1 0 26404 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_283
timestamp 1621523292
transform 1 0 27140 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a22o_1  _1142_
timestamp 1621523292
transform 1 0 29072 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1621523292
transform 1 0 27784 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1289_
timestamp 1621523292
transform 1 0 28428 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1621523292
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_286
timestamp 1621523292
transform 1 0 27416 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1621523292
transform 1 0 28060 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_300
timestamp 1621523292
transform 1 0 28704 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1621523292
transform 1 0 30820 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1299_
timestamp 1621523292
transform 1 0 30084 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_311
timestamp 1621523292
transform 1 0 29716 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_319
timestamp 1621523292
transform 1 0 30452 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1621523292
transform 1 0 33028 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1144_
timestamp 1621523292
transform 1 0 31648 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1621523292
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_328
timestamp 1621523292
transform 1 0 31280 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_337
timestamp 1621523292
transform 1 0 32108 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_341
timestamp 1621523292
transform 1 0 32476 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1621523292
transform 1 0 32660 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1621523292
transform 1 0 34132 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_350
timestamp 1621523292
transform 1 0 33304 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_358
timestamp 1621523292
transform 1 0 34040 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_362
timestamp 1621523292
transform 1 0 34408 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_370
timestamp 1621523292
transform 1 0 35144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1621523292
transform 1 0 35328 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1517_
timestamp 1621523292
transform 1 0 35972 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_375
timestamp 1621523292
transform 1 0 35604 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_382
timestamp 1621523292
transform 1 0 36248 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1621523292
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_394
timestamp 1621523292
transform 1 0 37352 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_398
timestamp 1621523292
transform 1 0 37720 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1621523292
transform 1 0 37904 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1621523292
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_424
timestamp 1621523292
transform 1 0 40112 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_436
timestamp 1621523292
transform 1 0 41216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1621523292
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_448
timestamp 1621523292
transform 1 0 42320 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1621523292
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1621523292
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_481
timestamp 1621523292
transform 1 0 45356 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_493
timestamp 1621523292
transform 1 0 46460 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1621523292
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1621523292
transform 1 0 47564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_514
timestamp 1621523292
transform 1 0 48392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_526
timestamp 1621523292
transform 1 0 49496 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_538
timestamp 1621523292
transform 1 0 50600 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1621523292
transform 1 0 51704 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_562
timestamp 1621523292
transform 1 0 52808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1617_
timestamp 1621523292
transform 1 0 54832 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1621523292
transform 1 0 53544 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_571
timestamp 1621523292
transform 1 0 53636 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_583
timestamp 1621523292
transform 1 0 54740 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_587
timestamp 1621523292
transform 1 0 55108 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2270_
timestamp 1621523292
transform 1 0 55476 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output220
timestamp 1621523292
transform 1 0 56764 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_599
timestamp 1621523292
transform 1 0 56212 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_609
timestamp 1621523292
transform 1 0 57132 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2308_
timestamp 1621523292
transform 1 0 57500 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1621523292
transform -1 0 58880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1621523292
transform 1 0 58236 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1676_
timestamp 1621523292
transform 1 0 2484 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1621523292
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output305
timestamp 1621523292
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1621523292
transform 1 0 1380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_11
timestamp 1621523292
transform 1 0 2116 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_18
timestamp 1621523292
transform 1 0 2760 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1621523292
transform 1 0 3128 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2500_
timestamp 1621523292
transform 1 0 4600 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1621523292
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_25
timestamp 1621523292
transform 1 0 3404 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_30
timestamp 1621523292
transform 1 0 3864 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1432_
timestamp 1621523292
transform 1 0 6900 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_54
timestamp 1621523292
transform 1 0 6072 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_62
timestamp 1621523292
transform 1 0 6808 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1430_
timestamp 1621523292
transform 1 0 7820 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1621523292
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_66
timestamp 1621523292
transform 1 0 7176 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_72
timestamp 1621523292
transform 1 0 7728 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_76
timestamp 1621523292
transform 1 0 8096 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1621523292
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_87
timestamp 1621523292
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1398_
timestamp 1621523292
transform 1 0 10120 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1434_
timestamp 1621523292
transform 1 0 9476 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1437_
timestamp 1621523292
transform 1 0 10948 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_38_94
timestamp 1621523292
transform 1 0 9752 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_101
timestamp 1621523292
transform 1 0 10396 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1416_
timestamp 1621523292
transform 1 0 12144 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_116
timestamp 1621523292
transform 1 0 11776 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_123
timestamp 1621523292
transform 1 0 12420 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_131
timestamp 1621523292
transform 1 0 13156 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1436_
timestamp 1621523292
transform 1 0 13248 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2499_
timestamp 1621523292
transform 1 0 14720 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1621523292
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_136
timestamp 1621523292
transform 1 0 13616 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_142
timestamp 1621523292
transform 1 0 14168 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_144
timestamp 1621523292
transform 1 0 14352 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1441_
timestamp 1621523292
transform 1 0 16928 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_164
timestamp 1621523292
transform 1 0 16192 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2519_
timestamp 1621523292
transform 1 0 17664 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_176
timestamp 1621523292
transform 1 0 17296 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_196
timestamp 1621523292
transform 1 0 19136 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1339_
timestamp 1621523292
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1621523292
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_201
timestamp 1621523292
transform 1 0 19596 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_213
timestamp 1621523292
transform 1 0 20700 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2518_
timestamp 1621523292
transform 1 0 21620 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_38_221
timestamp 1621523292
transform 1 0 21436 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_239
timestamp 1621523292
transform 1 0 23092 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1258_
timestamp 1621523292
transform 1 0 25208 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1322_
timestamp 1621523292
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1621523292
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1621523292
transform 1 0 24380 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_258
timestamp 1621523292
transform 1 0 24840 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2458_
timestamp 1621523292
transform 1 0 25944 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_38_266
timestamp 1621523292
transform 1 0 25576 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1621523292
transform 1 0 27784 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _1305_
timestamp 1621523292
transform 1 0 28704 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_286
timestamp 1621523292
transform 1 0 27416 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_293
timestamp 1621523292
transform 1 0 28060 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_299
timestamp 1621523292
transform 1 0 28612 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1191_
timestamp 1621523292
transform 1 0 31004 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1621523292
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_308
timestamp 1621523292
transform 1 0 29440 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_315
timestamp 1621523292
transform 1 0 30084 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_323
timestamp 1621523292
transform 1 0 30820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a221o_1  _1301_
timestamp 1621523292
transform 1 0 32200 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_334
timestamp 1621523292
transform 1 0 31832 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_346
timestamp 1621523292
transform 1 0 32936 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1138_
timestamp 1621523292
transform 1 0 33948 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1621523292
transform 1 0 33304 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1621523292
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_353
timestamp 1621523292
transform 1 0 33580 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_364
timestamp 1621523292
transform 1 0 34592 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_370
timestamp 1621523292
transform 1 0 35144 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1621523292
transform 1 0 35972 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_372
timestamp 1621523292
transform 1 0 35328 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_378
timestamp 1621523292
transform 1 0 35880 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_382
timestamp 1621523292
transform 1 0 36248 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_394
timestamp 1621523292
transform 1 0 37352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_406
timestamp 1621523292
transform 1 0 38456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1621523292
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_418
timestamp 1621523292
transform 1 0 39560 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_426
timestamp 1621523292
transform 1 0 40296 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1621523292
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1621523292
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1621523292
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1621523292
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1621523292
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1621523292
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1621523292
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_498
timestamp 1621523292
transform 1 0 46920 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_510
timestamp 1621523292
transform 1 0 48024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_522
timestamp 1621523292
transform 1 0 49128 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1621523292
transform 1 0 50968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_534
timestamp 1621523292
transform 1 0 50232 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_543
timestamp 1621523292
transform 1 0 51060 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_555
timestamp 1621523292
transform 1 0 52164 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_567
timestamp 1621523292
transform 1 0 53268 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1608_
timestamp 1621523292
transform 1 0 55292 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1613_
timestamp 1621523292
transform 1 0 54648 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_579
timestamp 1621523292
transform 1 0 54372 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_585
timestamp 1621523292
transform 1 0 54924 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2159_
timestamp 1621523292
transform 1 0 57224 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1621523292
transform 1 0 56212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_592
timestamp 1621523292
transform 1 0 55568 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_598
timestamp 1621523292
transform 1 0 56120 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_600
timestamp 1621523292
transform 1 0 56304 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_608
timestamp 1621523292
transform 1 0 57040 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1621523292
transform -1 0 58880 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output182
timestamp 1621523292
transform 1 0 57868 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_613
timestamp 1621523292
transform 1 0 57500 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_621
timestamp 1621523292
transform 1 0 58236 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2214_
timestamp 1621523292
transform 1 0 2116 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2216_
timestamp 1621523292
transform 1 0 1380 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2217_
timestamp 1621523292
transform 1 0 2484 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1621523292
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1621523292
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output306
timestamp 1621523292
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1621523292
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_19
timestamp 1621523292
transform 1 0 2852 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1621523292
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1440_
timestamp 1621523292
transform 1 0 4692 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2213_
timestamp 1621523292
transform 1 0 3220 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2506_
timestamp 1621523292
transform 1 0 4232 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1621523292
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_31
timestamp 1621523292
transform 1 0 3956 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_42
timestamp 1621523292
transform 1 0 4968 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_23
timestamp 1621523292
transform 1 0 3220 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_30
timestamp 1621523292
transform 1 0 3864 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1421_
timestamp 1621523292
transform 1 0 6072 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1439_
timestamp 1621523292
transform 1 0 5336 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2503_
timestamp 1621523292
transform 1 0 6808 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1621523292
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_53
timestamp 1621523292
transform 1 0 5980 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_58
timestamp 1621523292
transform 1 0 6440 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_50
timestamp 1621523292
transform 1 0 5704 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_61
timestamp 1621523292
transform 1 0 6716 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1393_
timestamp 1621523292
transform 1 0 8372 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1431_
timestamp 1621523292
transform 1 0 7268 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1489_
timestamp 1621523292
transform 1 0 8648 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1621523292
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_78
timestamp 1621523292
transform 1 0 8280 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_74
timestamp 1621523292
transform 1 0 7912 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_78
timestamp 1621523292
transform 1 0 8280 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_82
timestamp 1621523292
transform 1 0 8648 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_87
timestamp 1621523292
transform 1 0 9108 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1395_
timestamp 1621523292
transform 1 0 9568 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1473_
timestamp 1621523292
transform 1 0 10488 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2504_
timestamp 1621523292
transform 1 0 9476 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_39_88
timestamp 1621523292
transform 1 0 9200 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_95
timestamp 1621523292
transform 1 0 9844 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_101
timestamp 1621523292
transform 1 0 10396 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_108
timestamp 1621523292
transform 1 0 11040 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_107
timestamp 1621523292
transform 1 0 10948 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1418_
timestamp 1621523292
transform 1 0 11316 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1427_
timestamp 1621523292
transform 1 0 12696 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2507_
timestamp 1621523292
transform 1 0 12052 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1621523292
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_115
timestamp 1621523292
transform 1 0 11684 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_120
timestamp 1621523292
transform 1 0 12144 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_129
timestamp 1621523292
transform 1 0 12972 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_137
timestamp 1621523292
transform 1 0 13708 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_135
timestamp 1621523292
transform 1 0 13524 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1428_
timestamp 1621523292
transform 1 0 13340 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_144
timestamp 1621523292
transform 1 0 14352 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_143
timestamp 1621523292
transform 1 0 14260 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1621523292
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1433_
timestamp 1621523292
transform 1 0 13892 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_148
timestamp 1621523292
transform 1 0 14720 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_147
timestamp 1621523292
transform 1 0 14628 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1743_
timestamp 1621523292
transform 1 0 14812 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1445_
timestamp 1621523292
transform 1 0 14720 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1323_
timestamp 1621523292
transform 1 0 16192 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2546_
timestamp 1621523292
transform 1 0 15824 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1621523292
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_155
timestamp 1621523292
transform 1 0 15364 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_163
timestamp 1621523292
transform 1 0 16100 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_167
timestamp 1621523292
transform 1 0 16468 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_172
timestamp 1621523292
transform 1 0 16928 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_153
timestamp 1621523292
transform 1 0 15180 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_159
timestamp 1621523292
transform 1 0 15732 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1246_
timestamp 1621523292
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2100_
timestamp 1621523292
transform 1 0 17664 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1621523292
transform 1 0 17848 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1621523292
transform 1 0 18952 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_180
timestamp 1621523292
transform 1 0 17664 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_190
timestamp 1621523292
transform 1 0 18584 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_176
timestamp 1621523292
transform 1 0 17296 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_188
timestamp 1621523292
transform 1 0 18400 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_196
timestamp 1621523292
transform 1 0 19136 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 20056 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1621523292
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1621523292
transform 1 0 20240 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_202
timestamp 1621523292
transform 1 0 19688 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_211
timestamp 1621523292
transform 1 0 20516 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_201
timestamp 1621523292
transform 1 0 19596 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_207
timestamp 1621523292
transform 1 0 20148 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_216
timestamp 1621523292
transform 1 0 20976 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1621523292
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_224
timestamp 1621523292
transform 1 0 21712 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1621523292
transform 1 0 21252 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1069_
timestamp 1621523292
transform 1 0 21896 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_230
timestamp 1621523292
transform 1 0 22264 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 1621523292
transform 1 0 22172 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1621523292
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1222_
timestamp 1621523292
transform 1 0 22632 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1217_
timestamp 1621523292
transform 1 0 22540 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_238
timestamp 1621523292
transform 1 0 23000 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_237
timestamp 1621523292
transform 1 0 22908 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1065_
timestamp 1621523292
transform 1 0 24104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1226_
timestamp 1621523292
transform 1 0 23368 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2524_
timestamp 1621523292
transform 1 0 23644 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1621523292
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1621523292
transform 1 0 25116 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_246
timestamp 1621523292
transform 1 0 23736 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_253
timestamp 1621523292
transform 1 0 24380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_258
timestamp 1621523292
transform 1 0 24840 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_264
timestamp 1621523292
transform 1 0 25392 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1621523292
transform 1 0 25484 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1152_
timestamp 1621523292
transform 1 0 25484 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_40_272
timestamp 1621523292
transform 1 0 26128 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_277
timestamp 1621523292
transform 1 0 26588 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_273
timestamp 1621523292
transform 1 0 26220 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1259_
timestamp 1621523292
transform 1 0 26496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1621523292
transform 1 0 26680 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_280
timestamp 1621523292
transform 1 0 26864 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_281
timestamp 1621523292
transform 1 0 26956 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2528_
timestamp 1621523292
transform 1 0 27784 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1621523292
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1621523292
transform 1 0 27784 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1621523292
transform 1 0 28888 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1621523292
transform 1 0 27416 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_288
timestamp 1621523292
transform 1 0 27600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_298
timestamp 1621523292
transform 1 0 28520 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_310
timestamp 1621523292
transform 1 0 29624 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_314
timestamp 1621523292
transform 1 0 29992 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_306
timestamp 1621523292
transform 1 0 29256 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1621523292
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_315
timestamp 1621523292
transform 1 0 30084 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_320
timestamp 1621523292
transform 1 0 30544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1304_
timestamp 1621523292
transform 1 0 30452 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1298_
timestamp 1621523292
transform 1 0 30084 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_40_324
timestamp 1621523292
transform 1 0 30912 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1190_
timestamp 1621523292
transform 1 0 30912 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_40_332
timestamp 1621523292
transform 1 0 31648 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_338
timestamp 1621523292
transform 1 0 32200 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1621523292
transform 1 0 31556 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1621523292
transform 1 0 31924 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1277_
timestamp 1621523292
transform 1 0 31280 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_343
timestamp 1621523292
transform 1 0 32660 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_343
timestamp 1621523292
transform 1 0 32660 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1621523292
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o211a_1  _1302_
timestamp 1621523292
transform 1 0 33028 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1621523292
transform 1 0 32384 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2529_
timestamp 1621523292
transform 1 0 33028 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1621523292
transform 1 0 34132 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2463_
timestamp 1621523292
transform 1 0 34776 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1621523292
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_355
timestamp 1621523292
transform 1 0 33764 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_362
timestamp 1621523292
transform 1 0 34408 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1621523292
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1621523292
transform 1 0 35788 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1621523292
transform 1 0 36616 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_382
timestamp 1621523292
transform 1 0 36248 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_389
timestamp 1621523292
transform 1 0 36892 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_372
timestamp 1621523292
transform 1 0 35328 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_376
timestamp 1621523292
transform 1 0 35696 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_380
timestamp 1621523292
transform 1 0 36064 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_392
timestamp 1621523292
transform 1 0 37168 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1621523292
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_397
timestamp 1621523292
transform 1 0 37628 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1621523292
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_412
timestamp 1621523292
transform 1 0 39008 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_404
timestamp 1621523292
transform 1 0 38272 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1621523292
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_424
timestamp 1621523292
transform 1 0 40112 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_436
timestamp 1621523292
transform 1 0 41216 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_416
timestamp 1621523292
transform 1 0 39376 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_429
timestamp 1621523292
transform 1 0 40572 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1621523292
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_448
timestamp 1621523292
transform 1 0 42320 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1621523292
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_441
timestamp 1621523292
transform 1 0 41676 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_453
timestamp 1621523292
transform 1 0 42780 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1621523292
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_465
timestamp 1621523292
transform 1 0 43884 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_477
timestamp 1621523292
transform 1 0 44988 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1621523292
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1621523292
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1621523292
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_486
timestamp 1621523292
transform 1 0 45816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_498
timestamp 1621523292
transform 1 0 46920 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1621523292
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1621523292
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_514
timestamp 1621523292
transform 1 0 48392 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_510
timestamp 1621523292
transform 1 0 48024 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_522
timestamp 1621523292
transform 1 0 49128 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1621523292
transform 1 0 50968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_526
timestamp 1621523292
transform 1 0 49496 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_538
timestamp 1621523292
transform 1 0 50600 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_534
timestamp 1621523292
transform 1 0 50232 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_543
timestamp 1621523292
transform 1 0 51060 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_550
timestamp 1621523292
transform 1 0 51704 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_562
timestamp 1621523292
transform 1 0 52808 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_555
timestamp 1621523292
transform 1 0 52164 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_567
timestamp 1621523292
transform 1 0 53268 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1621523292
transform 1 0 53544 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1621523292
transform 1 0 55200 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_571
timestamp 1621523292
transform 1 0 53636 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_583
timestamp 1621523292
transform 1 0 54740 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_587
timestamp 1621523292
transform 1 0 55108 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_579
timestamp 1621523292
transform 1 0 54372 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_598
timestamp 1621523292
transform 1 0 56120 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_594
timestamp 1621523292
transform 1 0 55752 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_598
timestamp 1621523292
transform 1 0 56120 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2273_
timestamp 1621523292
transform 1 0 55384 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1612_
timestamp 1621523292
transform 1 0 55476 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_600
timestamp 1621523292
transform 1 0 56304 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_606
timestamp 1621523292
transform 1 0 56856 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_602
timestamp 1621523292
transform 1 0 56488 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1621523292
transform 1 0 56580 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1621523292
transform 1 0 56212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_608
timestamp 1621523292
transform 1 0 57040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1621523292
transform 1 0 57224 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2160_
timestamp 1621523292
transform 1 0 57224 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1621523292
transform -1 0 58880 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1621523292
transform -1 0 58880 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output183
timestamp 1621523292
transform 1 0 57868 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output221
timestamp 1621523292
transform 1 0 57868 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_613
timestamp 1621523292
transform 1 0 57500 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1621523292
transform 1 0 58236 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1621523292
transform 1 0 57500 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1621523292
transform 1 0 58236 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2218_
timestamp 1621523292
transform 1 0 1932 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1621523292
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_3
timestamp 1621523292
transform 1 0 1380 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_17
timestamp 1621523292
transform 1 0 2668 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1422_
timestamp 1621523292
transform 1 0 4692 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1786_
timestamp 1621523292
transform 1 0 3496 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_41_25
timestamp 1621523292
transform 1 0 3404 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_31
timestamp 1621523292
transform 1 0 3956 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_42
timestamp 1621523292
transform 1 0 4968 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1419_
timestamp 1621523292
transform 1 0 5336 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1621523292
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_49
timestamp 1621523292
transform 1 0 5612 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_58
timestamp 1621523292
transform 1 0 6440 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1411_
timestamp 1621523292
transform 1 0 7360 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1412_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 8004 0 1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__fill_2  FILLER_41_66
timestamp 1621523292
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1621523292
transform 1 0 7636 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_85
timestamp 1621523292
transform 1 0 8924 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1394_
timestamp 1621523292
transform 1 0 9292 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1429_
timestamp 1621523292
transform 1 0 10120 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_41_92
timestamp 1621523292
transform 1 0 9568 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_107
timestamp 1621523292
transform 1 0 10948 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1426_
timestamp 1621523292
transform 1 0 12604 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1621523292
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_113
timestamp 1621523292
transform 1 0 11500 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_115
timestamp 1621523292
transform 1 0 11684 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_123
timestamp 1621523292
transform 1 0 12420 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_128
timestamp 1621523292
transform 1 0 12880 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1379_
timestamp 1621523292
transform 1 0 13248 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2480_
timestamp 1621523292
transform 1 0 14536 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_41_137
timestamp 1621523292
transform 1 0 13708 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_145
timestamp 1621523292
transform 1 0 14444 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1621523292
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_162
timestamp 1621523292
transform 1 0 16008 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_170
timestamp 1621523292
transform 1 0 16744 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_172
timestamp 1621523292
transform 1 0 16928 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1535_
timestamp 1621523292
transform 1 0 17296 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2451_
timestamp 1621523292
transform 1 0 18308 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_41_181
timestamp 1621523292
transform 1 0 17756 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1231_
timestamp 1621523292
transform 1 0 20240 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1621523292
transform 1 0 20976 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_203
timestamp 1621523292
transform 1 0 19780 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_207
timestamp 1621523292
transform 1 0 20148 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_212
timestamp 1621523292
transform 1 0 20608 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1621523292
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1621523292
transform 1 0 22724 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_224
timestamp 1621523292
transform 1 0 21712 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_229
timestamp 1621523292
transform 1 0 22172 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1221_
timestamp 1621523292
transform 1 0 23828 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1223_
timestamp 1621523292
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_243
timestamp 1621523292
transform 1 0 23460 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_251
timestamp 1621523292
transform 1 0 24196 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_259
timestamp 1621523292
transform 1 0 24932 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2534_
timestamp 1621523292
transform 1 0 25484 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1621523292
transform 1 0 26956 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1621523292
transform 1 0 27784 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2530_
timestamp 1621523292
transform 1 0 29072 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1621523292
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_286
timestamp 1621523292
transform 1 0 27416 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_294
timestamp 1621523292
transform 1 0 28152 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_302
timestamp 1621523292
transform 1 0 28888 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1621523292
transform 1 0 30912 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_320
timestamp 1621523292
transform 1 0 30544 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_327
timestamp 1621523292
transform 1 0 31188 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1118_
timestamp 1621523292
transform 1 0 33212 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1295_
timestamp 1621523292
transform 1 0 31556 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1621523292
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_338
timestamp 1621523292
transform 1 0 32200 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_343
timestamp 1621523292
transform 1 0 32660 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2464_
timestamp 1621523292
transform 1 0 34592 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_41_356
timestamp 1621523292
transform 1 0 33856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1732_
timestamp 1621523292
transform 1 0 36432 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_41_380
timestamp 1621523292
transform 1 0 36064 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_389
timestamp 1621523292
transform 1 0 36892 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1621523292
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_397
timestamp 1621523292
transform 1 0 37628 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_400
timestamp 1621523292
transform 1 0 37904 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_412
timestamp 1621523292
transform 1 0 39008 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_424
timestamp 1621523292
transform 1 0 40112 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_436
timestamp 1621523292
transform 1 0 41216 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1621523292
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_448
timestamp 1621523292
transform 1 0 42320 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_457
timestamp 1621523292
transform 1 0 43148 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_469
timestamp 1621523292
transform 1 0 44252 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_481
timestamp 1621523292
transform 1 0 45356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_493
timestamp 1621523292
transform 1 0 46460 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1621523292
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1621523292
transform 1 0 47564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_514
timestamp 1621523292
transform 1 0 48392 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_526
timestamp 1621523292
transform 1 0 49496 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_538
timestamp 1621523292
transform 1 0 50600 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_550
timestamp 1621523292
transform 1 0 51704 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_562
timestamp 1621523292
transform 1 0 52808 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2275_
timestamp 1621523292
transform 1 0 54464 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1621523292
transform 1 0 53544 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_571
timestamp 1621523292
transform 1 0 53636 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_579
timestamp 1621523292
transform 1 0 54372 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_588
timestamp 1621523292
transform 1 0 55200 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1569_
timestamp 1621523292
transform 1 0 56856 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2274_
timestamp 1621523292
transform 1 0 55568 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_600
timestamp 1621523292
transform 1 0 56304 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_609
timestamp 1621523292
transform 1 0 57132 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2309_
timestamp 1621523292
transform 1 0 57500 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1621523292
transform -1 0 58880 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_621
timestamp 1621523292
transform 1 0 58236 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1787_
timestamp 1621523292
transform 1 0 2944 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1621523292
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output307
timestamp 1621523292
transform 1 0 1748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1621523292
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_11
timestamp 1621523292
transform 1 0 2116 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_19
timestamp 1621523292
transform 1 0 2852 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1425_
timestamp 1621523292
transform 1 0 5060 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1781_
timestamp 1621523292
transform 1 0 4232 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1621523292
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_25
timestamp 1621523292
transform 1 0 3404 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_30
timestamp 1621523292
transform 1 0 3864 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_39
timestamp 1621523292
transform 1 0 4692 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1410_
timestamp 1621523292
transform 1 0 6716 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1424_
timestamp 1621523292
transform 1 0 5704 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_42_46
timestamp 1621523292
transform 1 0 5336 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_57
timestamp 1621523292
transform 1 0 6348 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_65
timestamp 1621523292
transform 1 0 7084 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1413_
timestamp 1621523292
transform 1 0 7452 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1621523292
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1621523292
transform 1 0 8096 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_84
timestamp 1621523292
transform 1 0 8832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_87
timestamp 1621523292
transform 1 0 9108 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1381_
timestamp 1621523292
transform 1 0 9476 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2513_
timestamp 1621523292
transform 1 0 10764 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_95
timestamp 1621523292
transform 1 0 9844 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_103
timestamp 1621523292
transform 1 0 10580 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1377_
timestamp 1621523292
transform 1 0 12880 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_121
timestamp 1621523292
transform 1 0 12236 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_127
timestamp 1621523292
transform 1 0 12788 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_131
timestamp 1621523292
transform 1 0 13156 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1345_
timestamp 1621523292
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1380_
timestamp 1621523292
transform 1 0 13524 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1621523292
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_139
timestamp 1621523292
transform 1 0 13892 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_144
timestamp 1621523292
transform 1 0 14352 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_148
timestamp 1621523292
transform 1 0 14720 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1621523292
transform 1 0 15824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1531_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 16468 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1621523292
transform 1 0 15364 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_159
timestamp 1621523292
transform 1 0 15732 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_163
timestamp 1621523292
transform 1 0 16100 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_171
timestamp 1621523292
transform 1 0 16836 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1343_
timestamp 1621523292
transform 1 0 17204 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1536_
timestamp 1621523292
transform 1 0 17940 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_179
timestamp 1621523292
transform 1 0 17572 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_191
timestamp 1621523292
transform 1 0 18676 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2487_
timestamp 1621523292
transform 1 0 19964 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1621523292
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_199
timestamp 1621523292
transform 1 0 19412 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_201
timestamp 1621523292
transform 1 0 19596 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2540_
timestamp 1621523292
transform 1 0 21804 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_42_221
timestamp 1621523292
transform 1 0 21436 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1227_
timestamp 1621523292
transform 1 0 23828 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1275_
timestamp 1621523292
transform 1 0 25208 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1621523292
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_241
timestamp 1621523292
transform 1 0 23276 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_251
timestamp 1621523292
transform 1 0 24196 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_258
timestamp 1621523292
transform 1 0 24840 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2468_
timestamp 1621523292
transform 1 0 26864 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 1621523292
transform 1 0 26036 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_279
timestamp 1621523292
transform 1 0 26772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1296_
timestamp 1621523292
transform 1 0 28796 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_42_296
timestamp 1621523292
transform 1 0 28336 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_300
timestamp 1621523292
transform 1 0 28704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1195_
timestamp 1621523292
transform 1 0 31096 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1621523292
transform 1 0 30452 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1621523292
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_310
timestamp 1621523292
transform 1 0 29624 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_315
timestamp 1621523292
transform 1 0 30084 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_322
timestamp 1621523292
transform 1 0 30728 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1279_
timestamp 1621523292
transform 1 0 32292 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_42_335
timestamp 1621523292
transform 1 0 31924 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_346
timestamp 1621523292
transform 1 0 32936 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1186_
timestamp 1621523292
transform 1 0 33764 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1621523292
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_354
timestamp 1621523292
transform 1 0 33672 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_362
timestamp 1621523292
transform 1 0 34408 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_370
timestamp 1621523292
transform 1 0 35144 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1621523292
transform 1 0 35696 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1516_
timestamp 1621523292
transform 1 0 37168 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1733_
timestamp 1621523292
transform 1 0 36340 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_42_372
timestamp 1621523292
transform 1 0 35328 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_379
timestamp 1621523292
transform 1 0 35972 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_388
timestamp 1621523292
transform 1 0 36800 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_395
timestamp 1621523292
transform 1 0 37444 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_407
timestamp 1621523292
transform 1 0 38548 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1621523292
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_419
timestamp 1621523292
transform 1 0 39652 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_427
timestamp 1621523292
transform 1 0 40388 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_429
timestamp 1621523292
transform 1 0 40572 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_441
timestamp 1621523292
transform 1 0 41676 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_453
timestamp 1621523292
transform 1 0 42780 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_465
timestamp 1621523292
transform 1 0 43884 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1621523292
transform 1 0 44988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1621523292
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_486
timestamp 1621523292
transform 1 0 45816 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_498
timestamp 1621523292
transform 1 0 46920 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1621523292
transform 1 0 48024 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_522
timestamp 1621523292
transform 1 0 49128 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1621523292
transform 1 0 50968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_534
timestamp 1621523292
transform 1 0 50232 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_543
timestamp 1621523292
transform 1 0 51060 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_555
timestamp 1621523292
transform 1 0 52164 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_567
timestamp 1621523292
transform 1 0 53268 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_579
timestamp 1621523292
transform 1 0 54372 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_587
timestamp 1621523292
transform 1 0 55108 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1583_
timestamp 1621523292
transform 1 0 57040 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1611_
timestamp 1621523292
transform 1 0 55384 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1621523292
transform 1 0 56212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_593
timestamp 1621523292
transform 1 0 55660 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_600
timestamp 1621523292
transform 1 0 56304 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1568_
timestamp 1621523292
transform 1 0 57960 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1621523292
transform -1 0 58880 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_614
timestamp 1621523292
transform 1 0 57592 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1621523292
transform 1 0 58236 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2219_
timestamp 1621523292
transform 1 0 1932 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1621523292
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_3
timestamp 1621523292
transform 1 0 1380 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_17
timestamp 1621523292
transform 1 0 2668 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1782_
timestamp 1621523292
transform 1 0 3496 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2505_
timestamp 1621523292
transform 1 0 4508 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_43_25
timestamp 1621523292
transform 1 0 3404 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_31
timestamp 1621523292
transform 1 0 3956 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2508_
timestamp 1621523292
transform 1 0 6900 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1621523292
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_53
timestamp 1621523292
transform 1 0 5980 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_58
timestamp 1621523292
transform 1 0 6440 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_62
timestamp 1621523292
transform 1 0 6808 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2514_
timestamp 1621523292
transform 1 0 8740 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_43_79
timestamp 1621523292
transform 1 0 8372 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1621523292
transform 1 0 10580 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1621523292
transform 1 0 10212 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_106
timestamp 1621523292
transform 1 0 10856 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2509_
timestamp 1621523292
transform 1 0 12052 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1621523292
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_115
timestamp 1621523292
transform 1 0 11684 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1251_
timestamp 1621523292
transform 1 0 14904 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1420_
timestamp 1621523292
transform 1 0 13892 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_135
timestamp 1621523292
transform 1 0 13524 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_143
timestamp 1621523292
transform 1 0 14260 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_149
timestamp 1621523292
transform 1 0 14812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1621523292
transform 1 0 16192 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1621523292
transform 1 0 15548 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1621523292
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_153
timestamp 1621523292
transform 1 0 15180 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_160
timestamp 1621523292
transform 1 0 15824 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_167
timestamp 1621523292
transform 1 0 16468 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_172
timestamp 1621523292
transform 1 0 16928 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1228_
timestamp 1621523292
transform 1 0 18860 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1621523292
transform 1 0 17756 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_180
timestamp 1621523292
transform 1 0 17664 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1621523292
transform 1 0 18492 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1066_
timestamp 1621523292
transform 1 0 20240 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1621523292
transform 1 0 20976 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_202
timestamp 1621523292
transform 1 0 19688 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_212
timestamp 1621523292
transform 1 0 20608 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1621523292
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1621523292
transform 1 0 22540 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_224
timestamp 1621523292
transform 1 0 21712 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_229
timestamp 1621523292
transform 1 0 22172 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2535_
timestamp 1621523292
transform 1 0 24104 0 1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_43_241
timestamp 1621523292
transform 1 0 23276 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_249
timestamp 1621523292
transform 1 0 24012 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1272_
timestamp 1621523292
transform 1 0 25944 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_43_266
timestamp 1621523292
transform 1 0 25576 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_279
timestamp 1621523292
transform 1 0 26772 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1508_
timestamp 1621523292
transform 1 0 27784 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1514_
timestamp 1621523292
transform 1 0 28520 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1621523292
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1621523292
transform 1 0 27416 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_294
timestamp 1621523292
transform 1 0 28152 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_302
timestamp 1621523292
transform 1 0 28888 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1621523292
transform 1 0 29256 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1621523292
transform 1 0 29992 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1196_
timestamp 1621523292
transform 1 0 30636 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_309
timestamp 1621523292
transform 1 0 29532 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_313
timestamp 1621523292
transform 1 0 29900 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_317
timestamp 1621523292
transform 1 0 30268 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1127_
timestamp 1621523292
transform 1 0 31740 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1290_
timestamp 1621523292
transform 1 0 33028 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1621523292
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_329
timestamp 1621523292
transform 1 0 31372 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_338
timestamp 1621523292
transform 1 0 32200 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_343
timestamp 1621523292
transform 1 0 32660 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1621523292
transform 1 0 34776 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1187_
timestamp 1621523292
transform 1 0 34040 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_354
timestamp 1621523292
transform 1 0 33672 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_362
timestamp 1621523292
transform 1 0 34408 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_369
timestamp 1621523292
transform 1 0 35052 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1621523292
transform 1 0 35604 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1734_
timestamp 1621523292
transform 1 0 36248 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_43_378
timestamp 1621523292
transform 1 0 35880 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_387
timestamp 1621523292
transform 1 0 36708 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1621523292
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_400
timestamp 1621523292
transform 1 0 37904 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_412
timestamp 1621523292
transform 1 0 39008 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_424
timestamp 1621523292
transform 1 0 40112 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_436
timestamp 1621523292
transform 1 0 41216 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1621523292
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_448
timestamp 1621523292
transform 1 0 42320 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1621523292
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1621523292
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_481
timestamp 1621523292
transform 1 0 45356 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_493
timestamp 1621523292
transform 1 0 46460 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1621523292
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1621523292
transform 1 0 47564 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_514
timestamp 1621523292
transform 1 0 48392 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_526
timestamp 1621523292
transform 1 0 49496 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_538
timestamp 1621523292
transform 1 0 50600 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_550
timestamp 1621523292
transform 1 0 51704 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_562
timestamp 1621523292
transform 1 0 52808 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1609_
timestamp 1621523292
transform 1 0 55292 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1621523292
transform 1 0 53544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_571
timestamp 1621523292
transform 1 0 53636 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_583
timestamp 1621523292
transform 1 0 54740 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _1564_
timestamp 1621523292
transform 1 0 57224 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1610_
timestamp 1621523292
transform 1 0 55936 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1621523292
transform 1 0 56580 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_592
timestamp 1621523292
transform 1 0 55568 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_599
timestamp 1621523292
transform 1 0 56212 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_606
timestamp 1621523292
transform 1 0 56856 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1621523292
transform -1 0 58880 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output222
timestamp 1621523292
transform 1 0 57868 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_613
timestamp 1621523292
transform 1 0 57500 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_621
timestamp 1621523292
transform 1 0 58236 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2220_
timestamp 1621523292
transform 1 0 1840 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1621523292
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output308
timestamp 1621523292
transform 1 0 2944 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_3
timestamp 1621523292
transform 1 0 1380 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_7
timestamp 1621523292
transform 1 0 1748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1621523292
transform 1 0 2576 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1789_
timestamp 1621523292
transform 1 0 4508 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1621523292
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1621523292
transform 1 0 3312 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_28
timestamp 1621523292
transform 1 0 3680 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_30
timestamp 1621523292
transform 1 0 3864 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_36
timestamp 1621523292
transform 1 0 4416 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_40
timestamp 1621523292
transform 1 0 4784 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1414_
timestamp 1621523292
transform 1 0 6808 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1423_
timestamp 1621523292
transform 1 0 6164 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2102_
timestamp 1621523292
transform 1 0 5152 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_47
timestamp 1621523292
transform 1 0 5428 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1621523292
transform 1 0 6440 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_65
timestamp 1621523292
transform 1 0 7084 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1383_
timestamp 1621523292
transform 1 0 8372 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1384_
timestamp 1621523292
transform 1 0 7452 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1621523292
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_72
timestamp 1621523292
transform 1 0 7728 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_78
timestamp 1621523292
transform 1 0 8280 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_82
timestamp 1621523292
transform 1 0 8648 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_87
timestamp 1621523292
transform 1 0 9108 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1396_
timestamp 1621523292
transform 1 0 9752 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1399_
timestamp 1621523292
transform 1 0 10948 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_44_93
timestamp 1621523292
transform 1 0 9660 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_103
timestamp 1621523292
transform 1 0 10580 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1409_
timestamp 1621523292
transform 1 0 12144 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_116
timestamp 1621523292
transform 1 0 11776 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_129
timestamp 1621523292
transform 1 0 12972 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1392_
timestamp 1621523292
transform 1 0 13524 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2478_
timestamp 1621523292
transform 1 0 14720 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1621523292
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_139
timestamp 1621523292
transform 1 0 13892 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_144
timestamp 1621523292
transform 1 0 14352 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1213_
timestamp 1621523292
transform 1 0 16560 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_44_164
timestamp 1621523292
transform 1 0 16192 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1495_
timestamp 1621523292
transform 1 0 17572 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1621523292
transform 1 0 18308 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1621523292
transform 1 0 17204 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_183
timestamp 1621523292
transform 1 0 17940 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_195
timestamp 1621523292
transform 1 0 19044 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1621523292
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1621523292
transform 1 0 20148 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_199
timestamp 1621523292
transform 1 0 19412 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_201
timestamp 1621523292
transform 1 0 19596 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1621523292
transform 1 0 20884 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1234_
timestamp 1621523292
transform 1 0 23184 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1249_
timestamp 1621523292
transform 1 0 22356 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1250_
timestamp 1621523292
transform 1 0 21252 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1621523292
transform 1 0 21988 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_235
timestamp 1621523292
transform 1 0 22724 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_239
timestamp 1621523292
transform 1 0 23092 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _1274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 25208 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1294_
timestamp 1621523292
transform 1 0 23920 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1621523292
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_244
timestamp 1621523292
transform 1 0 23552 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_252
timestamp 1621523292
transform 1 0 24288 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_256
timestamp 1621523292
transform 1 0 24656 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1621523292
transform 1 0 24840 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1106_
timestamp 1621523292
transform 1 0 26588 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_44_269
timestamp 1621523292
transform 1 0 25852 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2532_
timestamp 1621523292
transform 1 0 28152 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_44_284
timestamp 1621523292
transform 1 0 27232 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_292
timestamp 1621523292
transform 1 0 27968 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  _1280_
timestamp 1621523292
transform 1 0 30912 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1621523292
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_310
timestamp 1621523292
transform 1 0 29624 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_315
timestamp 1621523292
transform 1 0 30084 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_323
timestamp 1621523292
transform 1 0 30820 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _1287_
timestamp 1621523292
transform 1 0 31740 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1292_
timestamp 1621523292
transform 1 0 32568 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_329
timestamp 1621523292
transform 1 0 31372 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_338
timestamp 1621523292
transform 1 0 32200 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1114_
timestamp 1621523292
transform 1 0 33672 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1621523292
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_350
timestamp 1621523292
transform 1 0 33304 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_361
timestamp 1621523292
transform 1 0 34316 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_369
timestamp 1621523292
transform 1 0 35052 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _1515_
timestamp 1621523292
transform 1 0 37076 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1735_
timestamp 1621523292
transform 1 0 36248 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_44_372
timestamp 1621523292
transform 1 0 35328 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_380
timestamp 1621523292
transform 1 0 36064 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_387
timestamp 1621523292
transform 1 0 36708 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_394
timestamp 1621523292
transform 1 0 37352 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_406
timestamp 1621523292
transform 1 0 38456 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1621523292
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_418
timestamp 1621523292
transform 1 0 39560 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_426
timestamp 1621523292
transform 1 0 40296 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_429
timestamp 1621523292
transform 1 0 40572 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_441
timestamp 1621523292
transform 1 0 41676 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_453
timestamp 1621523292
transform 1 0 42780 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_465
timestamp 1621523292
transform 1 0 43884 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_477
timestamp 1621523292
transform 1 0 44988 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1621523292
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_486
timestamp 1621523292
transform 1 0 45816 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_498
timestamp 1621523292
transform 1 0 46920 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_510
timestamp 1621523292
transform 1 0 48024 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_522
timestamp 1621523292
transform 1 0 49128 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1621523292
transform 1 0 50968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_534
timestamp 1621523292
transform 1 0 50232 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_543
timestamp 1621523292
transform 1 0 51060 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_555
timestamp 1621523292
transform 1 0 52164 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_567
timestamp 1621523292
transform 1 0 53268 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_1  _2276_
timestamp 1621523292
transform 1 0 55108 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_579
timestamp 1621523292
transform 1 0 54372 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _2161_
timestamp 1621523292
transform 1 0 56856 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1621523292
transform 1 0 56212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_595
timestamp 1621523292
transform 1 0 55844 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_600
timestamp 1621523292
transform 1 0 56304 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_609
timestamp 1621523292
transform 1 0 57132 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2310_
timestamp 1621523292
transform 1 0 57500 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1621523292
transform -1 0 58880 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_621
timestamp 1621523292
transform 1 0 58236 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1675_
timestamp 1621523292
transform 1 0 2576 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2221_
timestamp 1621523292
transform 1 0 1472 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1621523292
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_3
timestamp 1621523292
transform 1 0 1380 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_12
timestamp 1621523292
transform 1 0 2208 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_19
timestamp 1621523292
transform 1 0 2852 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1677_
timestamp 1621523292
transform 1 0 3220 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1621523292
transform 1 0 3864 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1788_
timestamp 1621523292
transform 1 0 4508 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_26
timestamp 1621523292
transform 1 0 3496 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1621523292
transform 1 0 4140 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_40
timestamp 1621523292
transform 1 0 4784 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1707_
timestamp 1621523292
transform 1 0 5244 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2515_
timestamp 1621523292
transform 1 0 6808 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1621523292
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_44
timestamp 1621523292
transform 1 0 5152 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1621523292
transform 1 0 5520 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_56
timestamp 1621523292
transform 1 0 6256 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_58
timestamp 1621523292
transform 1 0 6440 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1371_
timestamp 1621523292
transform 1 0 8648 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_78
timestamp 1621523292
transform 1 0 8280 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_86
timestamp 1621523292
transform 1 0 9016 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1388_
timestamp 1621523292
transform 1 0 9660 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1407_
timestamp 1621523292
transform 1 0 10396 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_45_92
timestamp 1621523292
transform 1 0 9568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_97
timestamp 1621523292
transform 1 0 10028 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1391_
timestamp 1621523292
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1417_
timestamp 1621523292
transform 1 0 12696 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1621523292
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_110
timestamp 1621523292
transform 1 0 11224 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1621523292
transform 1 0 11684 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_122
timestamp 1621523292
transform 1 0 12328 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_130
timestamp 1621523292
transform 1 0 13064 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1390_
timestamp 1621523292
transform 1 0 14904 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1397_
timestamp 1621523292
transform 1 0 13432 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1406_
timestamp 1621523292
transform 1 0 14168 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_138
timestamp 1621523292
transform 1 0 13800 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1621523292
transform 1 0 14536 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1621523292
transform 1 0 16192 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1621523292
transform 1 0 15548 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1621523292
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1621523292
transform 1 0 15180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_160
timestamp 1621523292
transform 1 0 15824 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_167
timestamp 1621523292
transform 1 0 16468 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1621523292
transform 1 0 16928 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1621523292
transform 1 0 18308 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1215_
timestamp 1621523292
transform 1 0 17296 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2544_
timestamp 1621523292
transform 1 0 18952 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_183
timestamp 1621523292
transform 1 0 17940 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1621523292
transform 1 0 18584 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1241_
timestamp 1621523292
transform 1 0 20976 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_210
timestamp 1621523292
transform 1 0 20424 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2474_
timestamp 1621523292
transform 1 0 22632 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1621523292
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_220
timestamp 1621523292
transform 1 0 21344 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1621523292
transform 1 0 22172 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_233
timestamp 1621523292
transform 1 0 22540 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__or2_2  _1109_
timestamp 1621523292
transform 1 0 25208 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1502_
timestamp 1621523292
transform 1 0 24472 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_250
timestamp 1621523292
transform 1 0 24104 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_258
timestamp 1621523292
transform 1 0 24840 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1260_
timestamp 1621523292
transform 1 0 26036 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_267
timestamp 1621523292
transform 1 0 25668 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_278
timestamp 1621523292
transform 1 0 26680 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1197_
timestamp 1621523292
transform 1 0 27784 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1288_
timestamp 1621523292
transform 1 0 28888 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1621523292
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_284
timestamp 1621523292
transform 1 0 27232 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1621523292
transform 1 0 27416 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_296
timestamp 1621523292
transform 1 0 28336 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1125_
timestamp 1621523292
transform 1 0 29992 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_45_310
timestamp 1621523292
transform 1 0 29624 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_321
timestamp 1621523292
transform 1 0 30636 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1621523292
transform 1 0 31464 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1293_
timestamp 1621523292
transform 1 0 33028 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1621523292
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_329
timestamp 1621523292
transform 1 0 31372 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_335
timestamp 1621523292
transform 1 0 31924 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_341
timestamp 1621523292
transform 1 0 32476 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_343
timestamp 1621523292
transform 1 0 32660 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1621523292
transform 1 0 34132 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2465_
timestamp 1621523292
transform 1 0 34776 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_45_355
timestamp 1621523292
transform 1 0 33764 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_362
timestamp 1621523292
transform 1 0 34408 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_382
timestamp 1621523292
transform 1 0 36248 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1621523292
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_394
timestamp 1621523292
transform 1 0 37352 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_398
timestamp 1621523292
transform 1 0 37720 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_400
timestamp 1621523292
transform 1 0 37904 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_412
timestamp 1621523292
transform 1 0 39008 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_424
timestamp 1621523292
transform 1 0 40112 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_436
timestamp 1621523292
transform 1 0 41216 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1621523292
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_448
timestamp 1621523292
transform 1 0 42320 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_457
timestamp 1621523292
transform 1 0 43148 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_469
timestamp 1621523292
transform 1 0 44252 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1621523292
transform 1 0 45356 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_493
timestamp 1621523292
transform 1 0 46460 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1621523292
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1621523292
transform 1 0 47564 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_514
timestamp 1621523292
transform 1 0 48392 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_526
timestamp 1621523292
transform 1 0 49496 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_538
timestamp 1621523292
transform 1 0 50600 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_550
timestamp 1621523292
transform 1 0 51704 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_562
timestamp 1621523292
transform 1 0 52808 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2277_
timestamp 1621523292
transform 1 0 55292 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1621523292
transform 1 0 53544 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_571
timestamp 1621523292
transform 1 0 53636 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_583
timestamp 1621523292
transform 1 0 54740 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1567_
timestamp 1621523292
transform 1 0 57224 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2162_
timestamp 1621523292
transform 1 0 56580 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_598
timestamp 1621523292
transform 1 0 56120 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_602
timestamp 1621523292
transform 1 0 56488 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_606
timestamp 1621523292
transform 1 0 56856 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1621523292
transform -1 0 58880 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output184
timestamp 1621523292
transform 1 0 57868 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_613
timestamp 1621523292
transform 1 0 57500 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1621523292
transform 1 0 58236 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_3
timestamp 1621523292
transform 1 0 1380 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_3
timestamp 1621523292
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output310
timestamp 1621523292
transform 1 0 1748 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output309
timestamp 1621523292
transform 1 0 1748 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1621523292
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1621523292
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_15
timestamp 1621523292
transform 1 0 2484 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_11
timestamp 1621523292
transform 1 0 2116 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_11
timestamp 1621523292
transform 1 0 2116 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2222_
timestamp 1621523292
transform 1 0 2576 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1621523292
transform 1 0 2484 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_18
timestamp 1621523292
transform 1 0 2760 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_30
timestamp 1621523292
transform 1 0 3864 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_25
timestamp 1621523292
transform 1 0 3404 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1621523292
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1674_
timestamp 1621523292
transform 1 0 3128 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_39
timestamp 1621523292
transform 1 0 4692 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_41
timestamp 1621523292
transform 1 0 4876 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1785_
timestamp 1621523292
transform 1 0 5060 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1784_
timestamp 1621523292
transform 1 0 4416 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1783_
timestamp 1621523292
transform 1 0 4600 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_24
timestamp 1621523292
transform 1 0 3312 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1404_
timestamp 1621523292
transform 1 0 7084 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_4  _2195_
timestamp 1621523292
transform 1 0 5244 0 -1 27744
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1621523292
transform 1 0 6348 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_58
timestamp 1621523292
transform 1 0 6440 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_46
timestamp 1621523292
transform 1 0 5336 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_54
timestamp 1621523292
transform 1 0 6072 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_58
timestamp 1621523292
transform 1 0 6440 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_64
timestamp 1621523292
transform 1 0 6992 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_72
timestamp 1621523292
transform 1 0 7728 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1621523292
transform 1 0 7820 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1386_
timestamp 1621523292
transform 1 0 7176 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_47_80
timestamp 1621523292
transform 1 0 8464 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1621523292
transform 1 0 9108 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1621523292
transform 1 0 8924 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_81
timestamp 1621523292
transform 1 0 8556 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1621523292
transform 1 0 9016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _1346_
timestamp 1621523292
transform 1 0 8188 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2516_
timestamp 1621523292
transform 1 0 8556 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_1  _1382_
timestamp 1621523292
transform 1 0 9476 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1389_
timestamp 1621523292
transform 1 0 10856 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2510_
timestamp 1621523292
transform 1 0 11040 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_46_98
timestamp 1621523292
transform 1 0 10120 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_106
timestamp 1621523292
transform 1 0 10856 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_97
timestamp 1621523292
transform 1 0 10028 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_105
timestamp 1621523292
transform 1 0 10764 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1494_
timestamp 1621523292
transform 1 0 12052 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1750_
timestamp 1621523292
transform 1 0 12696 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1621523292
transform 1 0 11592 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_124
timestamp 1621523292
transform 1 0 12512 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_110
timestamp 1621523292
transform 1 0 11224 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_115
timestamp 1621523292
transform 1 0 11684 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_122
timestamp 1621523292
transform 1 0 12328 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_132
timestamp 1621523292
transform 1 0 13248 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_138
timestamp 1621523292
transform 1 0 13800 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_132
timestamp 1621523292
transform 1 0 13248 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_1  _1408_
timestamp 1621523292
transform 1 0 13432 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1373_
timestamp 1621523292
transform 1 0 13616 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1621523292
transform 1 0 14720 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_144
timestamp 1621523292
transform 1 0 14352 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1621523292
transform 1 0 13984 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_144
timestamp 1621523292
transform 1 0 14352 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_142
timestamp 1621523292
transform 1 0 14168 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1621523292
transform 1 0 14260 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1481_
timestamp 1621523292
transform 1 0 14444 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_152
timestamp 1621523292
transform 1 0 15088 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1621523292
transform 1 0 15088 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_155
timestamp 1621523292
transform 1 0 15364 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_161
timestamp 1621523292
transform 1 0 15916 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1532_
timestamp 1621523292
transform 1 0 15180 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1071_
timestamp 1621523292
transform 1 0 15732 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_47_170
timestamp 1621523292
transform 1 0 16744 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_166
timestamp 1621523292
transform 1 0 16376 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_169
timestamp 1621523292
transform 1 0 16652 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1218_
timestamp 1621523292
transform 1 0 16284 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_172
timestamp 1621523292
transform 1 0 16928 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1621523292
transform 1 0 16836 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _1225_
timestamp 1621523292
transform 1 0 17020 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1621523292
transform 1 0 17296 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1534_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 18032 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2545_
timestamp 1621523292
transform 1 0 17940 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1621523292
transform 1 0 17664 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_191
timestamp 1621523292
transform 1 0 18676 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_179
timestamp 1621523292
transform 1 0 17572 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_199
timestamp 1621523292
transform 1 0 19412 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1621523292
transform 1 0 19596 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_199
timestamp 1621523292
transform 1 0 19412 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1621523292
transform 1 0 19504 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a221o_1  _1482_
timestamp 1621523292
transform 1 0 19964 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1219_
timestamp 1621523292
transform 1 0 19780 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_211
timestamp 1621523292
transform 1 0 20516 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1621523292
transform 1 0 20148 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1621523292
transform 1 0 20700 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1244_
timestamp 1621523292
transform 1 0 20608 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_217
timestamp 1621523292
transform 1 0 21068 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 21160 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_220
timestamp 1621523292
transform 1 0 21344 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_221
timestamp 1621523292
transform 1 0 21436 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1621523292
transform 1 0 21804 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_235
timestamp 1621523292
transform 1 0 22724 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_229
timestamp 1621523292
transform 1 0 22172 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1621523292
transform 1 0 22080 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1621523292
transform 1 0 22080 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _1206_
timestamp 1621523292
transform 1 0 22816 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1094_
timestamp 1621523292
transform 1 0 22448 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_46_239
timestamp 1621523292
transform 1 0 23092 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1621523292
transform 1 0 23460 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_246
timestamp 1621523292
transform 1 0 23736 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1621523292
transform 1 0 23828 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1621523292
transform 1 0 23460 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_250
timestamp 1621523292
transform 1 0 24104 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1621523292
transform 1 0 24380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1621523292
transform 1 0 24748 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _1270_
timestamp 1621523292
transform 1 0 24472 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1621523292
transform 1 0 24104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_261
timestamp 1621523292
transform 1 0 25116 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_258
timestamp 1621523292
transform 1 0 24840 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1621523292
transform 1 0 26496 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 25484 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1198_
timestamp 1621523292
transform 1 0 25944 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2469_
timestamp 1621523292
transform 1 0 27140 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_46_264
timestamp 1621523292
transform 1 0 25392 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_272
timestamp 1621523292
transform 1 0 26128 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1621523292
transform 1 0 26772 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_269
timestamp 1621523292
transform 1 0 25852 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_277
timestamp 1621523292
transform 1 0 26588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1621523292
transform 1 0 28980 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1261_
timestamp 1621523292
transform 1 0 27784 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2466_
timestamp 1621523292
transform 1 0 29072 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1621523292
transform 1 0 27324 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_299
timestamp 1621523292
transform 1 0 28612 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_286
timestamp 1621523292
transform 1 0 27416 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_297
timestamp 1621523292
transform 1 0 28428 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_303
timestamp 1621523292
transform 1 0 28980 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o32a_1  _1194_
timestamp 1621523292
transform 1 0 30912 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1281_
timestamp 1621523292
transform 1 0 30820 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1621523292
transform 1 0 29992 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_306
timestamp 1621523292
transform 1 0 29256 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_315
timestamp 1621523292
transform 1 0 30084 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_327
timestamp 1621523292
transform 1 0 31188 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_320
timestamp 1621523292
transform 1 0 30544 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1621523292
transform 1 0 32568 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1621523292
transform 1 0 33028 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1621523292
transform 1 0 31556 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1621523292
transform 1 0 32568 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_334
timestamp 1621523292
transform 1 0 31832 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_46_345
timestamp 1621523292
transform 1 0 32844 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_332
timestamp 1621523292
transform 1 0 31648 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_340
timestamp 1621523292
transform 1 0 32384 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_343
timestamp 1621523292
transform 1 0 32660 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1621523292
transform 1 0 33672 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1513_
timestamp 1621523292
transform 1 0 34316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2531_
timestamp 1621523292
transform 1 0 33396 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1621523292
transform 1 0 35236 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_367
timestamp 1621523292
transform 1 0 34868 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_350
timestamp 1621523292
transform 1 0 33304 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_357
timestamp 1621523292
transform 1 0 33948 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_364
timestamp 1621523292
transform 1 0 34592 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1731_
timestamp 1621523292
transform 1 0 35696 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1736_
timestamp 1621523292
transform 1 0 36156 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1739_
timestamp 1621523292
transform 1 0 35328 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_46_372
timestamp 1621523292
transform 1 0 35328 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_380
timestamp 1621523292
transform 1 0 36064 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_392
timestamp 1621523292
transform 1 0 37168 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_377
timestamp 1621523292
transform 1 0 35788 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_386
timestamp 1621523292
transform 1 0 36616 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1621523292
transform 1 0 37812 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_404
timestamp 1621523292
transform 1 0 38272 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_398
timestamp 1621523292
transform 1 0 37720 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_400
timestamp 1621523292
transform 1 0 37904 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_412
timestamp 1621523292
transform 1 0 39008 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1621523292
transform 1 0 40480 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_416
timestamp 1621523292
transform 1 0 39376 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_429
timestamp 1621523292
transform 1 0 40572 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_424
timestamp 1621523292
transform 1 0 40112 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_436
timestamp 1621523292
transform 1 0 41216 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1621523292
transform 1 0 43056 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_441
timestamp 1621523292
transform 1 0 41676 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_453
timestamp 1621523292
transform 1 0 42780 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_448
timestamp 1621523292
transform 1 0 42320 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_457
timestamp 1621523292
transform 1 0 43148 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_465
timestamp 1621523292
transform 1 0 43884 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_477
timestamp 1621523292
transform 1 0 44988 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_469
timestamp 1621523292
transform 1 0 44252 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1621523292
transform 1 0 45724 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_486
timestamp 1621523292
transform 1 0 45816 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_498
timestamp 1621523292
transform 1 0 46920 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_481
timestamp 1621523292
transform 1 0 45356 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_493
timestamp 1621523292
transform 1 0 46460 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1621523292
transform 1 0 48300 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_510
timestamp 1621523292
transform 1 0 48024 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_522
timestamp 1621523292
transform 1 0 49128 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_505
timestamp 1621523292
transform 1 0 47564 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_514
timestamp 1621523292
transform 1 0 48392 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1621523292
transform 1 0 50968 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_534
timestamp 1621523292
transform 1 0 50232 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_543
timestamp 1621523292
transform 1 0 51060 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_526
timestamp 1621523292
transform 1 0 49496 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_538
timestamp 1621523292
transform 1 0 50600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_555
timestamp 1621523292
transform 1 0 52164 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_567
timestamp 1621523292
transform 1 0 53268 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_550
timestamp 1621523292
transform 1 0 51704 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_562
timestamp 1621523292
transform 1 0 52808 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1606_
timestamp 1621523292
transform 1 0 55292 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1621523292
transform 1 0 53544 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_579
timestamp 1621523292
transform 1 0 54372 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_571
timestamp 1621523292
transform 1 0 53636 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_583
timestamp 1621523292
transform 1 0 54740 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_598
timestamp 1621523292
transform 1 0 56120 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_592
timestamp 1621523292
transform 1 0 55568 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_595
timestamp 1621523292
transform 1 0 55844 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_591
timestamp 1621523292
transform 1 0 55476 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1621523292
transform 1 0 55568 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_602
timestamp 1621523292
transform 1 0 56488 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_604
timestamp 1621523292
transform 1 0 56672 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_600
timestamp 1621523292
transform 1 0 56304 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output223
timestamp 1621523292
transform 1 0 56764 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1621523292
transform 1 0 56212 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1604_
timestamp 1621523292
transform 1 0 56212 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_609
timestamp 1621523292
transform 1 0 57132 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1566_
timestamp 1621523292
transform 1 0 57224 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2311_
timestamp 1621523292
transform 1 0 57500 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1621523292
transform -1 0 58880 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1621523292
transform -1 0 58880 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output185
timestamp 1621523292
transform 1 0 57868 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1621523292
transform 1 0 58236 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_613
timestamp 1621523292
transform 1 0 57500 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1621523292
transform 1 0 58236 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2103_
timestamp 1621523292
transform 1 0 2576 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2223_
timestamp 1621523292
transform 1 0 1472 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1621523292
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_3
timestamp 1621523292
transform 1 0 1380 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_12
timestamp 1621523292
transform 1 0 2208 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1621523292
transform 1 0 2852 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1790_
timestamp 1621523292
transform 1 0 4508 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1621523292
transform 1 0 3772 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_27
timestamp 1621523292
transform 1 0 3588 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_30
timestamp 1621523292
transform 1 0 3864 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_36
timestamp 1621523292
transform 1 0 4416 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_40
timestamp 1621523292
transform 1 0 4784 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1387_
timestamp 1621523292
transform 1 0 6992 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2511_
timestamp 1621523292
transform 1 0 5152 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_60
timestamp 1621523292
transform 1 0 6624 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1401_
timestamp 1621523292
transform 1 0 7636 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1621523292
transform 1 0 9016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_67
timestamp 1621523292
transform 1 0 7268 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_78
timestamp 1621523292
transform 1 0 8280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_87
timestamp 1621523292
transform 1 0 9108 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1374_
timestamp 1621523292
transform 1 0 9476 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1471_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 10672 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_98
timestamp 1621523292
transform 1 0 10120 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__o32a_1  _1470_
timestamp 1621523292
transform 1 0 12328 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_116
timestamp 1621523292
transform 1 0 11776 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1621523292
transform 1 0 13064 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1462_
timestamp 1621523292
transform 1 0 13432 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2479_
timestamp 1621523292
transform 1 0 14720 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1621523292
transform 1 0 14260 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_138
timestamp 1621523292
transform 1 0 13800 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_142
timestamp 1621523292
transform 1 0 14168 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_144
timestamp 1621523292
transform 1 0 14352 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1240_
timestamp 1621523292
transform 1 0 16560 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_164
timestamp 1621523292
transform 1 0 16192 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_171
timestamp 1621523292
transform 1 0 16836 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1621523292
transform 1 0 18400 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1752_
timestamp 1621523292
transform 1 0 17204 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_48_184
timestamp 1621523292
transform 1 0 18032 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_196
timestamp 1621523292
transform 1 0 19136 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2541_
timestamp 1621523292
transform 1 0 19964 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1621523292
transform 1 0 19504 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_201
timestamp 1621523292
transform 1 0 19596 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1091_
timestamp 1621523292
transform 1 0 21804 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1205_
timestamp 1621523292
transform 1 0 22908 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1621523292
transform 1 0 21436 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1621523292
transform 1 0 22448 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_236
timestamp 1621523292
transform 1 0 22816 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1621523292
transform 1 0 23920 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1621523292
transform 1 0 24748 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_244
timestamp 1621523292
transform 1 0 23552 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_251
timestamp 1621523292
transform 1 0 24196 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_258
timestamp 1621523292
transform 1 0 24840 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _1111_
timestamp 1621523292
transform 1 0 25484 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1248_
timestamp 1621523292
transform 1 0 26680 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_264
timestamp 1621523292
transform 1 0 25392 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_274
timestamp 1621523292
transform 1 0 26312 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_281
timestamp 1621523292
transform 1 0 26956 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1265_
timestamp 1621523292
transform 1 0 27416 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1266_
timestamp 1621523292
transform 1 0 28520 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_285
timestamp 1621523292
transform 1 0 27324 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_294
timestamp 1621523292
transform 1 0 28152 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _1120_
timestamp 1621523292
transform 1 0 30820 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1621523292
transform 1 0 29992 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_306
timestamp 1621523292
transform 1 0 29256 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_315
timestamp 1621523292
transform 1 0 30084 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1283_
timestamp 1621523292
transform 1 0 31648 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2533_
timestamp 1621523292
transform 1 0 33028 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_48_328
timestamp 1621523292
transform 1 0 31280 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_340
timestamp 1621523292
transform 1 0 32384 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_346
timestamp 1621523292
transform 1 0 32936 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1621523292
transform 1 0 35236 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_363
timestamp 1621523292
transform 1 0 34500 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1737_
timestamp 1621523292
transform 1 0 35696 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_372
timestamp 1621523292
transform 1 0 35328 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_380
timestamp 1621523292
transform 1 0 36064 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_392
timestamp 1621523292
transform 1 0 37168 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_404
timestamp 1621523292
transform 1 0 38272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1621523292
transform 1 0 40480 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_416
timestamp 1621523292
transform 1 0 39376 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_429
timestamp 1621523292
transform 1 0 40572 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_441
timestamp 1621523292
transform 1 0 41676 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_453
timestamp 1621523292
transform 1 0 42780 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_465
timestamp 1621523292
transform 1 0 43884 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_477
timestamp 1621523292
transform 1 0 44988 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1621523292
transform 1 0 45724 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_486
timestamp 1621523292
transform 1 0 45816 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_498
timestamp 1621523292
transform 1 0 46920 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_510
timestamp 1621523292
transform 1 0 48024 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_522
timestamp 1621523292
transform 1 0 49128 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1621523292
transform 1 0 50968 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_534
timestamp 1621523292
transform 1 0 50232 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_543
timestamp 1621523292
transform 1 0 51060 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_555
timestamp 1621523292
transform 1 0 52164 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_567
timestamp 1621523292
transform 1 0 53268 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__ebufn_2  _2278_
timestamp 1621523292
transform 1 0 55016 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1621523292
transform 1 0 54372 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_582
timestamp 1621523292
transform 1 0 54648 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2280_
timestamp 1621523292
transform 1 0 56672 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1621523292
transform 1 0 56212 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_595
timestamp 1621523292
transform 1 0 55844 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_600
timestamp 1621523292
transform 1 0 56304 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1621523292
transform -1 0 58880 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output224
timestamp 1621523292
transform 1 0 57868 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_613
timestamp 1621523292
transform 1 0 57500 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_621
timestamp 1621523292
transform 1 0 58236 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1621523292
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output312
timestamp 1621523292
transform 1 0 1748 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_3
timestamp 1621523292
transform 1 0 1380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_11
timestamp 1621523292
transform 1 0 2116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1621523292
transform 1 0 3220 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1621523292
transform 1 0 4324 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 1621523292
transform 1 0 5704 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2512_
timestamp 1621523292
transform 1 0 6808 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1621523292
transform 1 0 6348 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_47
timestamp 1621523292
transform 1 0 5428 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_53
timestamp 1621523292
transform 1 0 5980 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_58
timestamp 1621523292
transform 1 0 6440 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2517_
timestamp 1621523292
transform 1 0 8740 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_49_78
timestamp 1621523292
transform 1 0 8280 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_82
timestamp 1621523292
transform 1 0 8648 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1347_
timestamp 1621523292
transform 1 0 10580 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1621523292
transform 1 0 10212 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_106
timestamp 1621523292
transform 1 0 10856 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_2  _1368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 13064 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1468_
timestamp 1621523292
transform 1 0 12052 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1621523292
transform 1 0 11592 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_115
timestamp 1621523292
transform 1 0 11684 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_122
timestamp 1621523292
transform 1 0 12328 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1621523292
transform 1 0 14996 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1480_
timestamp 1621523292
transform 1 0 14076 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_137
timestamp 1621523292
transform 1 0 13708 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1621523292
transform 1 0 14536 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_150
timestamp 1621523292
transform 1 0 14904 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _1753_
timestamp 1621523292
transform 1 0 15640 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1621523292
transform 1 0 16836 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1621523292
transform 1 0 15272 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_167
timestamp 1621523292
transform 1 0 16468 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_172
timestamp 1621523292
transform 1 0 16928 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1236_
timestamp 1621523292
transform 1 0 18860 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1751_
timestamp 1621523292
transform 1 0 17296 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_49_185
timestamp 1621523292
transform 1 0 18124 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1245_
timestamp 1621523292
transform 1 0 20424 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_200
timestamp 1621523292
transform 1 0 19504 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_208
timestamp 1621523292
transform 1 0 20240 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_218
timestamp 1621523292
transform 1 0 21160 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _1207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 22908 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1621523292
transform 1 0 22080 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_226
timestamp 1621523292
transform 1 0 21896 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_229
timestamp 1621523292
transform 1 0 22172 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 1621523292
transform 1 0 25024 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _1208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 23736 0 1 28832
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_49_242
timestamp 1621523292
transform 1 0 23368 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_256
timestamp 1621523292
transform 1 0 24656 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1200_
timestamp 1621523292
transform 1 0 25852 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_49_263
timestamp 1621523292
transform 1 0 25300 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_278
timestamp 1621523292
transform 1 0 26680 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1262_
timestamp 1621523292
transform 1 0 27784 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _2537_
timestamp 1621523292
transform 1 0 28796 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1621523292
transform 1 0 27324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_284
timestamp 1621523292
transform 1 0 27232 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_286
timestamp 1621523292
transform 1 0 27416 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_297
timestamp 1621523292
transform 1 0 28428 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1621523292
transform 1 0 30912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_317
timestamp 1621523292
transform 1 0 30268 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_323
timestamp 1621523292
transform 1 0 30820 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_327
timestamp 1621523292
transform 1 0 31188 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1121_
timestamp 1621523292
transform 1 0 31556 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1284_
timestamp 1621523292
transform 1 0 33028 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1621523292
transform 1 0 32568 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_338
timestamp 1621523292
transform 1 0 32200 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_343
timestamp 1621523292
transform 1 0 32660 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_355
timestamp 1621523292
transform 1 0 33764 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_367
timestamp 1621523292
transform 1 0 34868 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1738_
timestamp 1621523292
transform 1 0 35420 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1740_
timestamp 1621523292
transform 1 0 36248 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_378
timestamp 1621523292
transform 1 0 35880 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_387
timestamp 1621523292
transform 1 0 36708 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1621523292
transform 1 0 37812 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_400
timestamp 1621523292
transform 1 0 37904 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_412
timestamp 1621523292
transform 1 0 39008 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_424
timestamp 1621523292
transform 1 0 40112 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_436
timestamp 1621523292
transform 1 0 41216 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1621523292
transform 1 0 43056 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_448
timestamp 1621523292
transform 1 0 42320 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_457
timestamp 1621523292
transform 1 0 43148 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_469
timestamp 1621523292
transform 1 0 44252 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_481
timestamp 1621523292
transform 1 0 45356 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_493
timestamp 1621523292
transform 1 0 46460 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1621523292
transform 1 0 48300 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_505
timestamp 1621523292
transform 1 0 47564 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_514
timestamp 1621523292
transform 1 0 48392 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_526
timestamp 1621523292
transform 1 0 49496 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_538
timestamp 1621523292
transform 1 0 50600 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_550
timestamp 1621523292
transform 1 0 51704 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_562
timestamp 1621523292
transform 1 0 52808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1603_
timestamp 1621523292
transform 1 0 54832 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2163_
timestamp 1621523292
transform 1 0 54188 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1621523292
transform 1 0 53544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_571
timestamp 1621523292
transform 1 0 53636 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_580
timestamp 1621523292
transform 1 0 54464 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_587
timestamp 1621523292
transform 1 0 55108 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1565_
timestamp 1621523292
transform 1 0 56120 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1601_
timestamp 1621523292
transform 1 0 55476 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output225
timestamp 1621523292
transform 1 0 56764 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_594
timestamp 1621523292
transform 1 0 55752 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_601
timestamp 1621523292
transform 1 0 56396 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_609
timestamp 1621523292
transform 1 0 57132 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2312_
timestamp 1621523292
transform 1 0 57500 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1621523292
transform -1 0 58880 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_621
timestamp 1621523292
transform 1 0 58236 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1621523292
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output313
timestamp 1621523292
transform 1 0 1748 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1621523292
transform 1 0 1380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_11
timestamp 1621523292
transform 1 0 2116 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1621523292
transform 1 0 3772 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_23
timestamp 1621523292
transform 1 0 3220 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_30
timestamp 1621523292
transform 1 0 3864 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_42
timestamp 1621523292
transform 1 0 4968 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1402_
timestamp 1621523292
transform 1 0 7084 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1403_
timestamp 1621523292
transform 1 0 6440 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1621523292
transform 1 0 6072 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_61
timestamp 1621523292
transform 1 0 6716 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1400_
timestamp 1621523292
transform 1 0 8096 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1621523292
transform 1 0 9016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_68
timestamp 1621523292
transform 1 0 7360 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_79
timestamp 1621523292
transform 1 0 8372 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1621523292
transform 1 0 8924 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_87
timestamp 1621523292
transform 1 0 9108 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1375_
timestamp 1621523292
transform 1 0 9476 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2491_
timestamp 1621523292
transform 1 0 10488 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_50_94
timestamp 1621523292
transform 1 0 9752 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1477_
timestamp 1621523292
transform 1 0 12328 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_118
timestamp 1621523292
transform 1 0 11960 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_131
timestamp 1621523292
transform 1 0 13156 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1621523292
transform 1 0 13616 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2477_
timestamp 1621523292
transform 1 0 14720 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1621523292
transform 1 0 14260 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_135
timestamp 1621523292
transform 1 0 13524 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_139
timestamp 1621523292
transform 1 0 13892 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_144
timestamp 1621523292
transform 1 0 14352 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1074_
timestamp 1621523292
transform 1 0 16560 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_164
timestamp 1621523292
transform 1 0 16192 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_171
timestamp 1621523292
transform 1 0 16836 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1212_
timestamp 1621523292
transform 1 0 18400 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _1754_
timestamp 1621523292
transform 1 0 17204 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_50_184
timestamp 1621523292
transform 1 0 18032 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_195
timestamp 1621523292
transform 1 0 19044 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1621523292
transform 1 0 19964 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2475_
timestamp 1621523292
transform 1 0 20884 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1621523292
transform 1 0 19504 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_199
timestamp 1621523292
transform 1 0 19412 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_201
timestamp 1621523292
transform 1 0 19596 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_208
timestamp 1621523292
transform 1 0 20240 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_214
timestamp 1621523292
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _1239_
timestamp 1621523292
transform 1 0 22724 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_231
timestamp 1621523292
transform 1 0 22356 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_239
timestamp 1621523292
transform 1 0 23092 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1238_
timestamp 1621523292
transform 1 0 23828 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1621523292
transform 1 0 25208 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1621523292
transform 1 0 24748 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1621523292
transform 1 0 24380 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1621523292
transform 1 0 24840 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1199_
timestamp 1621523292
transform 1 0 26128 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_50_265
timestamp 1621523292
transform 1 0 25484 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_271
timestamp 1621523292
transform 1 0 26036 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_279
timestamp 1621523292
transform 1 0 26772 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1621523292
transform 1 0 28980 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1102_
timestamp 1621523292
transform 1 0 27968 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1621523292
transform 1 0 27324 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_288
timestamp 1621523292
transform 1 0 27600 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_299
timestamp 1621523292
transform 1 0 28612 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2467_
timestamp 1621523292
transform 1 0 30452 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1621523292
transform 1 0 29992 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_306
timestamp 1621523292
transform 1 0 29256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_315
timestamp 1621523292
transform 1 0 30084 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1621523292
transform 1 0 32292 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_335
timestamp 1621523292
transform 1 0 31924 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_342
timestamp 1621523292
transform 1 0 32568 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1621523292
transform 1 0 35236 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_354
timestamp 1621523292
transform 1 0 33672 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_366
timestamp 1621523292
transform 1 0 34776 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_370
timestamp 1621523292
transform 1 0 35144 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_372
timestamp 1621523292
transform 1 0 35328 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1621523292
transform 1 0 36432 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_396
timestamp 1621523292
transform 1 0 37536 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_408
timestamp 1621523292
transform 1 0 38640 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1621523292
transform 1 0 40480 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_420
timestamp 1621523292
transform 1 0 39744 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_429
timestamp 1621523292
transform 1 0 40572 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_441
timestamp 1621523292
transform 1 0 41676 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_453
timestamp 1621523292
transform 1 0 42780 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_465
timestamp 1621523292
transform 1 0 43884 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_477
timestamp 1621523292
transform 1 0 44988 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1621523292
transform 1 0 45724 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_486
timestamp 1621523292
transform 1 0 45816 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_498
timestamp 1621523292
transform 1 0 46920 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_510
timestamp 1621523292
transform 1 0 48024 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_522
timestamp 1621523292
transform 1 0 49128 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1621523292
transform 1 0 50968 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_534
timestamp 1621523292
transform 1 0 50232 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_543
timestamp 1621523292
transform 1 0 51060 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_555
timestamp 1621523292
transform 1 0 52164 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_567
timestamp 1621523292
transform 1 0 53268 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1602_
timestamp 1621523292
transform 1 0 54372 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2281_
timestamp 1621523292
transform 1 0 55016 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1621523292
transform 1 0 53728 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_571
timestamp 1621523292
transform 1 0 53636 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_575
timestamp 1621523292
transform 1 0 54004 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_582
timestamp 1621523292
transform 1 0 54648 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2279_
timestamp 1621523292
transform 1 0 56672 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1621523292
transform 1 0 56212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_595
timestamp 1621523292
transform 1 0 55844 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_600
timestamp 1621523292
transform 1 0 56304 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1621523292
transform -1 0 58880 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output186
timestamp 1621523292
transform 1 0 57868 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1621523292
transform 1 0 57500 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1621523292
transform 1 0 58236 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1621523292
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1621523292
transform 1 0 1380 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_6
timestamp 1621523292
transform 1 0 1656 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_18
timestamp 1621523292
transform 1 0 2760 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_30
timestamp 1621523292
transform 1 0 3864 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_42
timestamp 1621523292
transform 1 0 4968 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1621523292
transform 1 0 6348 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_54
timestamp 1621523292
transform 1 0 6072 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_58
timestamp 1621523292
transform 1 0 6440 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_70
timestamp 1621523292
transform 1 0 7544 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_82
timestamp 1621523292
transform 1 0 8648 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1533_
timestamp 1621523292
transform 1 0 10948 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 10304 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_wb_clk_i
timestamp 1621523292
transform 1 0 9476 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_90
timestamp 1621523292
transform 1 0 9384 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_94
timestamp 1621523292
transform 1 0 9752 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_103
timestamp 1621523292
transform 1 0 10580 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _1367_
timestamp 1621523292
transform 1 0 12420 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1621523292
transform 1 0 11592 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_110
timestamp 1621523292
transform 1 0 11224 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_115
timestamp 1621523292
transform 1 0 11684 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1621523292
transform 1 0 15088 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 13616 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_132
timestamp 1621523292
transform 1 0 13248 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_142
timestamp 1621523292
transform 1 0 14168 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_150
timestamp 1621523292
transform 1 0 14904 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o32a_1  _1211_
timestamp 1621523292
transform 1 0 15732 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1621523292
transform 1 0 16836 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_155
timestamp 1621523292
transform 1 0 15364 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_167
timestamp 1621523292
transform 1 0 16468 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_172
timestamp 1621523292
transform 1 0 16928 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _1075_
timestamp 1621523292
transform 1 0 17296 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1229_
timestamp 1621523292
transform 1 0 18308 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_51_183
timestamp 1621523292
transform 1 0 17940 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_194
timestamp 1621523292
transform 1 0 18952 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1621523292
transform 1 0 20608 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1237_
timestamp 1621523292
transform 1 0 19412 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_51_198
timestamp 1621523292
transform 1 0 19320 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_208
timestamp 1621523292
transform 1 0 20240 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_215
timestamp 1621523292
transform 1 0 20884 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1621523292
transform 1 0 21344 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1621523292
transform 1 0 22816 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1621523292
transform 1 0 22080 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_219
timestamp 1621523292
transform 1 0 21252 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_223
timestamp 1621523292
transform 1 0 21620 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_227
timestamp 1621523292
transform 1 0 21988 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_229
timestamp 1621523292
transform 1 0 22172 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_235
timestamp 1621523292
transform 1 0 22724 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_239
timestamp 1621523292
transform 1 0 23092 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2538_
timestamp 1621523292
transform 1 0 23460 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_51_259
timestamp 1621523292
transform 1 0 24932 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1621523292
transform 1 0 26588 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1268_
timestamp 1621523292
transform 1 0 25484 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_51_272
timestamp 1621523292
transform 1 0 26128 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_276
timestamp 1621523292
transform 1 0 26496 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_280
timestamp 1621523292
transform 1 0 26864 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1621523292
transform 1 0 27784 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1621523292
transform 1 0 28520 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1263_
timestamp 1621523292
transform 1 0 29164 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1621523292
transform 1 0 27324 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_284
timestamp 1621523292
transform 1 0 27232 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_286
timestamp 1621523292
transform 1 0 27416 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1621523292
transform 1 0 28060 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_297
timestamp 1621523292
transform 1 0 28428 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_301
timestamp 1621523292
transform 1 0 28796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1509_
timestamp 1621523292
transform 1 0 29808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1510_
timestamp 1621523292
transform 1 0 30452 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1621523292
transform 1 0 31096 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_308
timestamp 1621523292
transform 1 0 29440 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_315
timestamp 1621523292
transform 1 0 30084 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_322
timestamp 1621523292
transform 1 0 30728 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1621523292
transform 1 0 32568 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_329
timestamp 1621523292
transform 1 0 31372 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1621523292
transform 1 0 32476 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1621523292
transform 1 0 32660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1621523292
transform 1 0 33764 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1621523292
transform 1 0 34868 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_371
timestamp 1621523292
transform 1 0 35236 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _1741_
timestamp 1621523292
transform 1 0 35328 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1742_
timestamp 1621523292
transform 1 0 36156 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_51_377
timestamp 1621523292
transform 1 0 35788 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_386
timestamp 1621523292
transform 1 0 36616 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1621523292
transform 1 0 37812 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_398
timestamp 1621523292
transform 1 0 37720 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_400
timestamp 1621523292
transform 1 0 37904 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_412
timestamp 1621523292
transform 1 0 39008 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_424
timestamp 1621523292
transform 1 0 40112 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_436
timestamp 1621523292
transform 1 0 41216 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1621523292
transform 1 0 43056 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_448
timestamp 1621523292
transform 1 0 42320 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_457
timestamp 1621523292
transform 1 0 43148 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_469
timestamp 1621523292
transform 1 0 44252 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_481
timestamp 1621523292
transform 1 0 45356 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_493
timestamp 1621523292
transform 1 0 46460 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1621523292
transform 1 0 48300 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1621523292
transform 1 0 47564 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_514
timestamp 1621523292
transform 1 0 48392 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_526
timestamp 1621523292
transform 1 0 49496 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_538
timestamp 1621523292
transform 1 0 50600 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_550
timestamp 1621523292
transform 1 0 51704 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_562
timestamp 1621523292
transform 1 0 52808 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1605_
timestamp 1621523292
transform 1 0 54556 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2282_
timestamp 1621523292
transform 1 0 55200 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1621523292
transform 1 0 53544 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_571
timestamp 1621523292
transform 1 0 53636 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_579
timestamp 1621523292
transform 1 0 54372 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_584
timestamp 1621523292
transform 1 0 54832 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output187
timestamp 1621523292
transform 1 0 56764 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_597
timestamp 1621523292
transform 1 0 56028 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_609
timestamp 1621523292
transform 1 0 57132 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2313_
timestamp 1621523292
transform 1 0 57500 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1621523292
transform -1 0 58880 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_621
timestamp 1621523292
transform 1 0 58236 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1621523292
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1621523292
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1621523292
transform 1 0 1380 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_6
timestamp 1621523292
transform 1 0 1656 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_18
timestamp 1621523292
transform 1 0 2760 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1621523292
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1621523292
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1621523292
transform 1 0 3772 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_26
timestamp 1621523292
transform 1 0 3496 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_30
timestamp 1621523292
transform 1 0 3864 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_42
timestamp 1621523292
transform 1 0 4968 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1621523292
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1621523292
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1621523292
transform 1 0 6348 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_54
timestamp 1621523292
transform 1 0 6072 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_51
timestamp 1621523292
transform 1 0 5796 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_58
timestamp 1621523292
transform 1 0 6440 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1621523292
transform 1 0 9016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_66
timestamp 1621523292
transform 1 0 7176 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_78
timestamp 1621523292
transform 1 0 8280 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_87
timestamp 1621523292
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_70
timestamp 1621523292
transform 1 0 7544 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_82
timestamp 1621523292
transform 1 0 8648 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1760_
timestamp 1621523292
transform 1 0 10948 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_wb_clk_i
timestamp 1621523292
transform 1 0 10304 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_99
timestamp 1621523292
transform 1 0 10212 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_103
timestamp 1621523292
transform 1 0 10580 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_94
timestamp 1621523292
transform 1 0 9752 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_106
timestamp 1621523292
transform 1 0 10856 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1362_
timestamp 1621523292
transform 1 0 12420 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1365_
timestamp 1621523292
transform 1 0 11776 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1372_
timestamp 1621523292
transform 1 0 12420 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1621523292
transform 1 0 11592 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_110
timestamp 1621523292
transform 1 0 11224 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_119
timestamp 1621523292
transform 1 0 12052 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_115
timestamp 1621523292
transform 1 0 11684 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_139
timestamp 1621523292
transform 1 0 13892 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_132
timestamp 1621523292
transform 1 0 13248 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_139
timestamp 1621523292
transform 1 0 13892 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_132
timestamp 1621523292
transform 1 0 13248 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 13616 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1621523292
transform 1 0 13616 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_148
timestamp 1621523292
transform 1 0 14720 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_144
timestamp 1621523292
transform 1 0 14352 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1621523292
transform 1 0 14260 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1497_
timestamp 1621523292
transform 1 0 14444 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_152
timestamp 1621523292
transform 1 0 15088 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1621523292
transform 1 0 15272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1744_
timestamp 1621523292
transform 1 0 15456 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2543_
timestamp 1621523292
transform 1 0 15916 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1621523292
transform 1 0 16836 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1621523292
transform 1 0 15548 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_162
timestamp 1621523292
transform 1 0 16008 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_170
timestamp 1621523292
transform 1 0 16744 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_172
timestamp 1621523292
transform 1 0 16928 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1621523292
transform 1 0 18860 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1079_
timestamp 1621523292
transform 1 0 19044 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1232_
timestamp 1621523292
transform 1 0 17756 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1621523292
transform 1 0 17572 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_177
timestamp 1621523292
transform 1 0 17388 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_189
timestamp 1621523292
transform 1 0 18492 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_196
timestamp 1621523292
transform 1 0 19136 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_178
timestamp 1621523292
transform 1 0 17480 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_187
timestamp 1621523292
transform 1 0 18308 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1621523292
transform 1 0 20056 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1254_
timestamp 1621523292
transform 1 0 20976 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2542_
timestamp 1621523292
transform 1 0 19964 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1621523292
transform 1 0 19504 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_201
timestamp 1621523292
transform 1 0 19596 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_202
timestamp 1621523292
transform 1 0 19688 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_209
timestamp 1621523292
transform 1 0 20332 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_215
timestamp 1621523292
transform 1 0 20884 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_224
timestamp 1621523292
transform 1 0 21712 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_228
timestamp 1621523292
transform 1 0 22080 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_221
timestamp 1621523292
transform 1 0 21436 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1621523292
transform 1 0 22080 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1621523292
transform 1 0 21804 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_229
timestamp 1621523292
transform 1 0 22172 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_236
timestamp 1621523292
transform 1 0 22816 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1257_
timestamp 1621523292
transform 1 0 23000 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1252_
timestamp 1621523292
transform 1 0 22540 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_53_240
timestamp 1621523292
transform 1 0 23184 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _1256_
timestamp 1621523292
transform 1 0 23552 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1269_
timestamp 1621523292
transform 1 0 25208 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2536_
timestamp 1621523292
transform 1 0 25116 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1621523292
transform 1 0 24748 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_247
timestamp 1621523292
transform 1 0 23828 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_255
timestamp 1621523292
transform 1 0 24564 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1621523292
transform 1 0 24840 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_251
timestamp 1621523292
transform 1 0 24196 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_259
timestamp 1621523292
transform 1 0 24932 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_1  _1098_
timestamp 1621523292
transform 1 0 26404 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_52_271
timestamp 1621523292
transform 1 0 26036 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_282
timestamp 1621523292
transform 1 0 27048 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_277
timestamp 1621523292
transform 1 0 26588 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1507_
timestamp 1621523292
transform 1 0 27784 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2470_
timestamp 1621523292
transform 1 0 27416 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1621523292
transform 1 0 27324 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_302
timestamp 1621523292
transform 1 0 28888 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1621523292
transform 1 0 27416 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1621523292
transform 1 0 28060 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_305
timestamp 1621523292
transform 1 0 29164 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1621523292
transform 1 0 29256 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1621523292
transform 1 0 29992 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_309
timestamp 1621523292
transform 1 0 29532 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_313
timestamp 1621523292
transform 1 0 29900 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_315
timestamp 1621523292
transform 1 0 30084 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_327
timestamp 1621523292
transform 1 0 31188 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_317
timestamp 1621523292
transform 1 0 30268 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1917_
timestamp 1621523292
transform 1 0 33028 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1621523292
transform 1 0 32568 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_339
timestamp 1621523292
transform 1 0 32292 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_329
timestamp 1621523292
transform 1 0 31372 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 1621523292
transform 1 0 32476 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_343
timestamp 1621523292
transform 1 0 32660 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1915_
timestamp 1621523292
transform 1 0 33948 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1919_
timestamp 1621523292
transform 1 0 34592 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1621523292
transform 1 0 35236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_351
timestamp 1621523292
transform 1 0 33396 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_363
timestamp 1621523292
transform 1 0 34500 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_353
timestamp 1621523292
transform 1 0 33580 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_360
timestamp 1621523292
transform 1 0 34224 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1621523292
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_372
timestamp 1621523292
transform 1 0 35328 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_384
timestamp 1621523292
transform 1 0 36432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1621523292
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_391
timestamp 1621523292
transform 1 0 37076 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1621523292
transform 1 0 37812 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_396
timestamp 1621523292
transform 1 0 37536 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_408
timestamp 1621523292
transform 1 0 38640 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_400
timestamp 1621523292
transform 1 0 37904 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1621523292
transform 1 0 39008 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1621523292
transform 1 0 40480 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_420
timestamp 1621523292
transform 1 0 39744 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_429
timestamp 1621523292
transform 1 0 40572 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_424
timestamp 1621523292
transform 1 0 40112 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1621523292
transform 1 0 41216 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1621523292
transform 1 0 43056 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_441
timestamp 1621523292
transform 1 0 41676 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_453
timestamp 1621523292
transform 1 0 42780 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_448
timestamp 1621523292
transform 1 0 42320 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_457
timestamp 1621523292
transform 1 0 43148 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_465
timestamp 1621523292
transform 1 0 43884 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_477
timestamp 1621523292
transform 1 0 44988 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_469
timestamp 1621523292
transform 1 0 44252 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1621523292
transform 1 0 45724 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_486
timestamp 1621523292
transform 1 0 45816 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_498
timestamp 1621523292
transform 1 0 46920 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_481
timestamp 1621523292
transform 1 0 45356 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_493
timestamp 1621523292
transform 1 0 46460 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1621523292
transform 1 0 48300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_510
timestamp 1621523292
transform 1 0 48024 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_522
timestamp 1621523292
transform 1 0 49128 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1621523292
transform 1 0 47564 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_514
timestamp 1621523292
transform 1 0 48392 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1621523292
transform 1 0 50968 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_534
timestamp 1621523292
transform 1 0 50232 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_543
timestamp 1621523292
transform 1 0 51060 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_526
timestamp 1621523292
transform 1 0 49496 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_538
timestamp 1621523292
transform 1 0 50600 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1621523292
transform 1 0 52900 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_555
timestamp 1621523292
transform 1 0 52164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_567
timestamp 1621523292
transform 1 0 53268 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1621523292
transform 1 0 51704 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_562
timestamp 1621523292
transform 1 0 52808 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_566
timestamp 1621523292
transform 1 0 53176 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_571
timestamp 1621523292
transform 1 0 53636 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_574
timestamp 1621523292
transform 1 0 53912 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1621523292
transform 1 0 53544 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2164_
timestamp 1621523292
transform 1 0 53636 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_581
timestamp 1621523292
transform 1 0 54556 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2283_
timestamp 1621523292
transform 1 0 54372 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1600_
timestamp 1621523292
transform 1 0 54280 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1593_
timestamp 1621523292
transform 1 0 54924 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_588
timestamp 1621523292
transform 1 0 55200 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_588
timestamp 1621523292
transform 1 0 55200 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_595
timestamp 1621523292
transform 1 0 55844 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_600
timestamp 1621523292
transform 1 0 56304 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_595
timestamp 1621523292
transform 1 0 55844 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1621523292
transform 1 0 56212 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1592_
timestamp 1621523292
transform 1 0 55568 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1591_
timestamp 1621523292
transform 1 0 55568 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1589_
timestamp 1621523292
transform 1 0 56212 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_602
timestamp 1621523292
transform 1 0 56488 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1621523292
transform 1 0 56856 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1621523292
transform 1 0 56488 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_4  _2291_
timestamp 1621523292
transform 1 0 57040 0 1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__ebufn_4  _2290_
timestamp 1621523292
transform 1 0 56672 0 -1 31008
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1621523292
transform -1 0 58880 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1621523292
transform -1 0 58880 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_617
timestamp 1621523292
transform 1 0 57868 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_621
timestamp 1621523292
transform 1 0 58236 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1621523292
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1621523292
transform 1 0 1380 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_6
timestamp 1621523292
transform 1 0 1656 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_18
timestamp 1621523292
transform 1 0 2760 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1621523292
transform 1 0 3772 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_26
timestamp 1621523292
transform 1 0 3496 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_30
timestamp 1621523292
transform 1 0 3864 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_42
timestamp 1621523292
transform 1 0 4968 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_54
timestamp 1621523292
transform 1 0 6072 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1621523292
transform 1 0 9016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_66
timestamp 1621523292
transform 1 0 7176 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_78
timestamp 1621523292
transform 1 0 8280 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_87
timestamp 1621523292
transform 1 0 9108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_99
timestamp 1621523292
transform 1 0 10212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _1378_
timestamp 1621523292
transform 1 0 12420 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_111
timestamp 1621523292
transform 1 0 11316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1364_
timestamp 1621523292
transform 1 0 13616 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1498_
timestamp 1621523292
transform 1 0 14904 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1621523292
transform 1 0 14260 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_132
timestamp 1621523292
transform 1 0 13248 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_139
timestamp 1621523292
transform 1 0 13892 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_144
timestamp 1621523292
transform 1 0 14352 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1499_
timestamp 1621523292
transform 1 0 15548 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1530_
timestamp 1621523292
transform 1 0 16192 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 16836 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1621523292
transform 1 0 15180 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_160
timestamp 1621523292
transform 1 0 15824 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1621523292
transform 1 0 16468 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_174
timestamp 1621523292
transform 1 0 17112 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2476_
timestamp 1621523292
transform 1 0 17664 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_196
timestamp 1621523292
transform 1 0 19136 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1621523292
transform 1 0 21160 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _1749_
timestamp 1621523292
transform 1 0 19964 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1621523292
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_201
timestamp 1621523292
transform 1 0 19596 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_214
timestamp 1621523292
transform 1 0 20792 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1088_
timestamp 1621523292
transform 1 0 22264 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1504_
timestamp 1621523292
transform 1 0 23092 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1621523292
transform 1 0 21896 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_235
timestamp 1621523292
transform 1 0 22724 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1747_
timestamp 1621523292
transform 1 0 25208 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1621523292
transform 1 0 24748 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_242
timestamp 1621523292
transform 1 0 23368 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_254
timestamp 1621523292
transform 1 0 24472 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_258
timestamp 1621523292
transform 1 0 24840 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1621523292
transform 1 0 26404 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2471_
timestamp 1621523292
transform 1 0 27048 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_54_271
timestamp 1621523292
transform 1 0 26036 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_278
timestamp 1621523292
transform 1 0 26680 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_298
timestamp 1621523292
transform 1 0 28520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1621523292
transform 1 0 29992 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_310
timestamp 1621523292
transform 1 0 29624 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_315
timestamp 1621523292
transform 1 0 30084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_327
timestamp 1621523292
transform 1 0 31188 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2392_
timestamp 1621523292
transform 1 0 32108 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_54_335
timestamp 1621523292
transform 1 0 31924 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_1  _1920_
timestamp 1621523292
transform 1 0 34224 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1621523292
transform 1 0 35236 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_353
timestamp 1621523292
transform 1 0 33580 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_359
timestamp 1621523292
transform 1 0 34132 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_367
timestamp 1621523292
transform 1 0 34868 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1918_
timestamp 1621523292
transform 1 0 35696 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_372
timestamp 1621523292
transform 1 0 35328 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_379
timestamp 1621523292
transform 1 0 35972 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_391
timestamp 1621523292
transform 1 0 37076 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_403
timestamp 1621523292
transform 1 0 38180 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1621523292
transform 1 0 40480 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_415
timestamp 1621523292
transform 1 0 39284 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_427
timestamp 1621523292
transform 1 0 40388 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_429
timestamp 1621523292
transform 1 0 40572 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_441
timestamp 1621523292
transform 1 0 41676 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_453
timestamp 1621523292
transform 1 0 42780 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_465
timestamp 1621523292
transform 1 0 43884 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_477
timestamp 1621523292
transform 1 0 44988 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1621523292
transform 1 0 45724 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_486
timestamp 1621523292
transform 1 0 45816 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_498
timestamp 1621523292
transform 1 0 46920 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_510
timestamp 1621523292
transform 1 0 48024 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_522
timestamp 1621523292
transform 1 0 49128 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1621523292
transform 1 0 50968 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_534
timestamp 1621523292
transform 1 0 50232 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_543
timestamp 1621523292
transform 1 0 51060 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_555
timestamp 1621523292
transform 1 0 52164 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_567
timestamp 1621523292
transform 1 0 53268 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1594_
timestamp 1621523292
transform 1 0 54372 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1597_
timestamp 1621523292
transform 1 0 53728 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2286_
timestamp 1621523292
transform 1 0 55016 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_54_571
timestamp 1621523292
transform 1 0 53636 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_575
timestamp 1621523292
transform 1 0 54004 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_582
timestamp 1621523292
transform 1 0 54648 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1621523292
transform 1 0 56212 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output227
timestamp 1621523292
transform 1 0 56672 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1621523292
transform 1 0 57224 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_595
timestamp 1621523292
transform 1 0 55844 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_600
timestamp 1621523292
transform 1 0 56304 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_608
timestamp 1621523292
transform 1 0 57040 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_2  _2289_
timestamp 1621523292
transform 1 0 57408 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1621523292
transform -1 0 58880 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_621
timestamp 1621523292
transform 1 0 58236 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1621523292
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1621523292
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1621523292
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1621523292
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1621523292
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1621523292
transform 1 0 6348 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_51
timestamp 1621523292
transform 1 0 5796 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_58
timestamp 1621523292
transform 1 0 6440 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_70
timestamp 1621523292
transform 1 0 7544 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_82
timestamp 1621523292
transform 1 0 8648 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_94
timestamp 1621523292
transform 1 0 9752 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_106
timestamp 1621523292
transform 1 0 10856 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1483_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 13156 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1621523292
transform 1 0 11592 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_115
timestamp 1621523292
transform 1 0 11684 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_127
timestamp 1621523292
transform 1 0 12788 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1500_
timestamp 1621523292
transform 1 0 14628 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_138
timestamp 1621523292
transform 1 0 13800 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_146
timestamp 1621523292
transform 1 0 14536 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_150
timestamp 1621523292
transform 1 0 14904 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1621523292
transform 1 0 16836 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_wb_clk_i
timestamp 1621523292
transform 1 0 15272 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_157
timestamp 1621523292
transform 1 0 15548 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1621523292
transform 1 0 16652 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_172
timestamp 1621523292
transform 1 0 16928 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1501_
timestamp 1621523292
transform 1 0 17940 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_180
timestamp 1621523292
transform 1 0 17664 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_186
timestamp 1621523292
transform 1 0 18216 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1621523292
transform 1 0 19412 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1503_
timestamp 1621523292
transform 1 0 20792 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_55_198
timestamp 1621523292
transform 1 0 19320 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_202
timestamp 1621523292
transform 1 0 19688 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_217
timestamp 1621523292
transform 1 0 21068 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1087_
timestamp 1621523292
transform 1 0 22908 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1621523292
transform 1 0 21436 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1621523292
transform 1 0 22080 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_224
timestamp 1621523292
transform 1 0 21712 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_229
timestamp 1621523292
transform 1 0 22172 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1621523292
transform 1 0 23920 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1748_
timestamp 1621523292
transform 1 0 24932 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_55_244
timestamp 1621523292
transform 1 0 23552 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_251
timestamp 1621523292
transform 1 0 24196 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1621523292
transform 1 0 26128 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_268
timestamp 1621523292
transform 1 0 25760 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_275
timestamp 1621523292
transform 1 0 26404 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_283
timestamp 1621523292
transform 1 0 27140 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1621523292
transform 1 0 27324 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_286
timestamp 1621523292
transform 1 0 27416 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_298
timestamp 1621523292
transform 1 0 28520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2391_
timestamp 1621523292
transform 1 0 30544 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_55_310
timestamp 1621523292
transform 1 0 29624 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_318
timestamp 1621523292
transform 1 0 30360 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1912_
timestamp 1621523292
transform 1 0 33028 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1621523292
transform 1 0 32568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_336
timestamp 1621523292
transform 1 0 32016 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_343
timestamp 1621523292
transform 1 0 32660 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2393_
timestamp 1621523292
transform 1 0 33856 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_55_350
timestamp 1621523292
transform 1 0 33304 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_372
timestamp 1621523292
transform 1 0 35328 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_384
timestamp 1621523292
transform 1 0 36432 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1621523292
transform 1 0 37812 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_396
timestamp 1621523292
transform 1 0 37536 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_400
timestamp 1621523292
transform 1 0 37904 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_412
timestamp 1621523292
transform 1 0 39008 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_424
timestamp 1621523292
transform 1 0 40112 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_436
timestamp 1621523292
transform 1 0 41216 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1621523292
transform 1 0 43056 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_448
timestamp 1621523292
transform 1 0 42320 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_457
timestamp 1621523292
transform 1 0 43148 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_469
timestamp 1621523292
transform 1 0 44252 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_481
timestamp 1621523292
transform 1 0 45356 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_493
timestamp 1621523292
transform 1 0 46460 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1621523292
transform 1 0 48300 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1621523292
transform 1 0 47564 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_514
timestamp 1621523292
transform 1 0 48392 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_526
timestamp 1621523292
transform 1 0 49496 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_538
timestamp 1621523292
transform 1 0 50600 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1621523292
transform 1 0 51704 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_562
timestamp 1621523292
transform 1 0 52808 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1596_
timestamp 1621523292
transform 1 0 54372 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1621523292
transform 1 0 53544 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_571
timestamp 1621523292
transform 1 0 53636 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_582
timestamp 1621523292
transform 1 0 54648 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1590_
timestamp 1621523292
transform 1 0 55476 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  _2292_
timestamp 1621523292
transform 1 0 56120 0 1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1621523292
transform 1 0 55936 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_590
timestamp 1621523292
transform 1 0 55384 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_594
timestamp 1621523292
transform 1 0 55752 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_611
timestamp 1621523292
transform 1 0 57316 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1621523292
transform -1 0 58880 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output189
timestamp 1621523292
transform 1 0 57868 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1621523292
transform 1 0 58236 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1621523292
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1621523292
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1621523292
transform 1 0 1656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_18
timestamp 1621523292
transform 1 0 2760 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1621523292
transform 1 0 3772 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_26
timestamp 1621523292
transform 1 0 3496 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_30
timestamp 1621523292
transform 1 0 3864 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_42
timestamp 1621523292
transform 1 0 4968 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_54
timestamp 1621523292
transform 1 0 6072 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1621523292
transform 1 0 9016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_66
timestamp 1621523292
transform 1 0 7176 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_78
timestamp 1621523292
transform 1 0 8280 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1621523292
transform 1 0 9108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1621523292
transform 1 0 10212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_111
timestamp 1621523292
transform 1 0 11316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_123
timestamp 1621523292
transform 1 0 12420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1621523292
transform 1 0 14260 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_135
timestamp 1621523292
transform 1 0 13524 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_144
timestamp 1621523292
transform 1 0 14352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_156
timestamp 1621523292
transform 1 0 15456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_168
timestamp 1621523292
transform 1 0 16560 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_180
timestamp 1621523292
transform 1 0 17664 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_192
timestamp 1621523292
transform 1 0 18768 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2539_
timestamp 1621523292
transform 1 0 19964 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1621523292
transform 1 0 19504 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_201
timestamp 1621523292
transform 1 0 19596 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1083_
timestamp 1621523292
transform 1 0 21804 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1202_
timestamp 1621523292
transform 1 0 22816 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_56_221
timestamp 1621523292
transform 1 0 21436 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_232
timestamp 1621523292
transform 1 0 22448 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1506_
timestamp 1621523292
transform 1 0 23828 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _1745_
timestamp 1621523292
transform 1 0 25208 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1621523292
transform 1 0 24748 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_243
timestamp 1621523292
transform 1 0 23460 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_250
timestamp 1621523292
transform 1 0 24104 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_256
timestamp 1621523292
transform 1 0 24656 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_258
timestamp 1621523292
transform 1 0 24840 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_271
timestamp 1621523292
transform 1 0 26036 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_283
timestamp 1621523292
transform 1 0 27140 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_295
timestamp 1621523292
transform 1 0 28244 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1621523292
transform 1 0 29992 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_307
timestamp 1621523292
transform 1 0 29348 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_313
timestamp 1621523292
transform 1 0 29900 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_315
timestamp 1621523292
transform 1 0 30084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_327
timestamp 1621523292
transform 1 0 31188 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1914_
timestamp 1621523292
transform 1 0 31556 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _1916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 32844 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_335
timestamp 1621523292
transform 1 0 31924 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_343
timestamp 1621523292
transform 1 0 32660 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1923_
timestamp 1621523292
transform 1 0 34040 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1621523292
transform 1 0 35236 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_354
timestamp 1621523292
transform 1 0 33672 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_367
timestamp 1621523292
transform 1 0 34868 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1925_
timestamp 1621523292
transform 1 0 35696 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_372
timestamp 1621523292
transform 1 0 35328 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_382
timestamp 1621523292
transform 1 0 36248 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_394
timestamp 1621523292
transform 1 0 37352 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_406
timestamp 1621523292
transform 1 0 38456 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1621523292
transform 1 0 40480 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_418
timestamp 1621523292
transform 1 0 39560 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_426
timestamp 1621523292
transform 1 0 40296 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_429
timestamp 1621523292
transform 1 0 40572 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_441
timestamp 1621523292
transform 1 0 41676 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_453
timestamp 1621523292
transform 1 0 42780 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_465
timestamp 1621523292
transform 1 0 43884 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_477
timestamp 1621523292
transform 1 0 44988 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1621523292
transform 1 0 45724 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_486
timestamp 1621523292
transform 1 0 45816 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_498
timestamp 1621523292
transform 1 0 46920 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_510
timestamp 1621523292
transform 1 0 48024 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_522
timestamp 1621523292
transform 1 0 49128 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1621523292
transform 1 0 50968 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_534
timestamp 1621523292
transform 1 0 50232 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_543
timestamp 1621523292
transform 1 0 51060 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_555
timestamp 1621523292
transform 1 0 52164 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_567
timestamp 1621523292
transform 1 0 53268 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1599_
timestamp 1621523292
transform 1 0 53636 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2284_
timestamp 1621523292
transform 1 0 54280 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_56_574
timestamp 1621523292
transform 1 0 53912 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_587
timestamp 1621523292
transform 1 0 55108 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1595_
timestamp 1621523292
transform 1 0 55568 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_2  _2288_
timestamp 1621523292
transform 1 0 57132 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1621523292
transform 1 0 56212 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_591
timestamp 1621523292
transform 1 0 55476 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_595
timestamp 1621523292
transform 1 0 55844 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_600
timestamp 1621523292
transform 1 0 56304 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_608
timestamp 1621523292
transform 1 0 57040 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1621523292
transform -1 0 58880 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_618
timestamp 1621523292
transform 1 0 57960 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_624
timestamp 1621523292
transform 1 0 58512 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1621523292
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1621523292
transform 1 0 1380 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_6
timestamp 1621523292
transform 1 0 1656 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_18
timestamp 1621523292
transform 1 0 2760 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_30
timestamp 1621523292
transform 1 0 3864 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1621523292
transform 1 0 4968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1621523292
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_54
timestamp 1621523292
transform 1 0 6072 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_58
timestamp 1621523292
transform 1 0 6440 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_70
timestamp 1621523292
transform 1 0 7544 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_82
timestamp 1621523292
transform 1 0 8648 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1621523292
transform 1 0 9752 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_106
timestamp 1621523292
transform 1 0 10856 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1621523292
transform 1 0 11592 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_115
timestamp 1621523292
transform 1 0 11684 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_127
timestamp 1621523292
transform 1 0 12788 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_139
timestamp 1621523292
transform 1 0 13892 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_151
timestamp 1621523292
transform 1 0 14996 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1621523292
transform 1 0 16836 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_163
timestamp 1621523292
transform 1 0 16100 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_172
timestamp 1621523292
transform 1 0 16928 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1621523292
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1621523292
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1505_
timestamp 1621523292
transform 1 0 20608 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_208
timestamp 1621523292
transform 1 0 20240 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_215
timestamp 1621523292
transform 1 0 20884 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1621523292
transform 1 0 21252 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1621523292
transform 1 0 22632 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1621523292
transform 1 0 22080 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_222
timestamp 1621523292
transform 1 0 21528 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_229
timestamp 1621523292
transform 1 0 22172 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_233
timestamp 1621523292
transform 1 0 22540 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1621523292
transform 1 0 22908 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2472_
timestamp 1621523292
transform 1 0 23460 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_57_259
timestamp 1621523292
transform 1 0 24932 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1746_
timestamp 1621523292
transform 1 0 25300 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_57_272
timestamp 1621523292
transform 1 0 26128 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1621523292
transform 1 0 27324 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_284
timestamp 1621523292
transform 1 0 27232 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_286
timestamp 1621523292
transform 1 0 27416 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_298
timestamp 1621523292
transform 1 0 28520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _1910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 31188 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_57_310
timestamp 1621523292
transform 1 0 29624 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_322
timestamp 1621523292
transform 1 0 30728 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_326
timestamp 1621523292
transform 1 0 31096 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1913_
timestamp 1621523292
transform 1 0 33028 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1621523292
transform 1 0 32568 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_332
timestamp 1621523292
transform 1 0 31648 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_340
timestamp 1621523292
transform 1 0 32384 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_343
timestamp 1621523292
transform 1 0 32660 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2394_
timestamp 1621523292
transform 1 0 33948 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_57_350
timestamp 1621523292
transform 1 0 33304 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_356
timestamp 1621523292
transform 1 0 33856 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1922_
timestamp 1621523292
transform 1 0 35788 0 1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1621523292
transform 1 0 35420 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_382
timestamp 1621523292
transform 1 0 36248 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1621523292
transform 1 0 37812 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_394
timestamp 1621523292
transform 1 0 37352 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_398
timestamp 1621523292
transform 1 0 37720 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_400
timestamp 1621523292
transform 1 0 37904 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_412
timestamp 1621523292
transform 1 0 39008 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_424
timestamp 1621523292
transform 1 0 40112 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_436
timestamp 1621523292
transform 1 0 41216 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1621523292
transform 1 0 43056 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_448
timestamp 1621523292
transform 1 0 42320 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_457
timestamp 1621523292
transform 1 0 43148 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_469
timestamp 1621523292
transform 1 0 44252 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_481
timestamp 1621523292
transform 1 0 45356 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_493
timestamp 1621523292
transform 1 0 46460 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1621523292
transform 1 0 48300 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_505
timestamp 1621523292
transform 1 0 47564 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_514
timestamp 1621523292
transform 1 0 48392 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_526
timestamp 1621523292
transform 1 0 49496 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_538
timestamp 1621523292
transform 1 0 50600 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_550
timestamp 1621523292
transform 1 0 51704 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_562
timestamp 1621523292
transform 1 0 52808 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_2  _2287_
timestamp 1621523292
transform 1 0 54280 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1621523292
transform 1 0 53544 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1621523292
transform 1 0 54096 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_571
timestamp 1621523292
transform 1 0 53636 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_575
timestamp 1621523292
transform 1 0 54004 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_587
timestamp 1621523292
transform 1 0 55108 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _2285_
timestamp 1621523292
transform 1 0 55568 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output228
timestamp 1621523292
transform 1 0 56764 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_591
timestamp 1621523292
transform 1 0 55476 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_601
timestamp 1621523292
transform 1 0 56396 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_609
timestamp 1621523292
transform 1 0 57132 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2314_
timestamp 1621523292
transform 1 0 57500 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1621523292
transform -1 0 58880 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1621523292
transform 1 0 58236 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1621523292
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1621523292
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1621523292
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1621523292
transform 1 0 3772 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1621523292
transform 1 0 3588 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_30
timestamp 1621523292
transform 1 0 3864 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_42
timestamp 1621523292
transform 1 0 4968 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_54
timestamp 1621523292
transform 1 0 6072 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1621523292
transform 1 0 9016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_66
timestamp 1621523292
transform 1 0 7176 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_78
timestamp 1621523292
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_87
timestamp 1621523292
transform 1 0 9108 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_99
timestamp 1621523292
transform 1 0 10212 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_111
timestamp 1621523292
transform 1 0 11316 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_123
timestamp 1621523292
transform 1 0 12420 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1621523292
transform 1 0 14260 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1621523292
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_144
timestamp 1621523292
transform 1 0 14352 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_156
timestamp 1621523292
transform 1 0 15456 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_168
timestamp 1621523292
transform 1 0 16560 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_180
timestamp 1621523292
transform 1 0 17664 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_192
timestamp 1621523292
transform 1 0 18768 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2473_
timestamp 1621523292
transform 1 0 20976 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1621523292
transform 1 0 19504 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_201
timestamp 1621523292
transform 1 0 19596 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_213
timestamp 1621523292
transform 1 0 20700 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1203_
timestamp 1621523292
transform 1 0 22816 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_58_232
timestamp 1621523292
transform 1 0 22448 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1621523292
transform 1 0 24748 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_243
timestamp 1621523292
transform 1 0 23460 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_255
timestamp 1621523292
transform 1 0 24564 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_258
timestamp 1621523292
transform 1 0 24840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_270
timestamp 1621523292
transform 1 0 25944 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_282
timestamp 1621523292
transform 1 0 27048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_294
timestamp 1621523292
transform 1 0 28152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2390_
timestamp 1621523292
transform 1 0 30452 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1621523292
transform 1 0 29992 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_306
timestamp 1621523292
transform 1 0 29256 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_315
timestamp 1621523292
transform 1 0 30084 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2395_
timestamp 1621523292
transform 1 0 32292 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_58_335
timestamp 1621523292
transform 1 0 31924 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1924_
timestamp 1621523292
transform 1 0 34132 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1621523292
transform 1 0 35236 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_355
timestamp 1621523292
transform 1 0 33764 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_362
timestamp 1621523292
transform 1 0 34408 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_370
timestamp 1621523292
transform 1 0 35144 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1921_
timestamp 1621523292
transform 1 0 35696 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_372
timestamp 1621523292
transform 1 0 35328 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_379
timestamp 1621523292
transform 1 0 35972 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_391
timestamp 1621523292
transform 1 0 37076 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_403
timestamp 1621523292
transform 1 0 38180 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1621523292
transform 1 0 40480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_415
timestamp 1621523292
transform 1 0 39284 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_427
timestamp 1621523292
transform 1 0 40388 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_429
timestamp 1621523292
transform 1 0 40572 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_441
timestamp 1621523292
transform 1 0 41676 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_453
timestamp 1621523292
transform 1 0 42780 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_465
timestamp 1621523292
transform 1 0 43884 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_477
timestamp 1621523292
transform 1 0 44988 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1621523292
transform 1 0 45724 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_486
timestamp 1621523292
transform 1 0 45816 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_498
timestamp 1621523292
transform 1 0 46920 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_510
timestamp 1621523292
transform 1 0 48024 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_522
timestamp 1621523292
transform 1 0 49128 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1621523292
transform 1 0 50968 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_534
timestamp 1621523292
transform 1 0 50232 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_543
timestamp 1621523292
transform 1 0 51060 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_555
timestamp 1621523292
transform 1 0 52164 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_567
timestamp 1621523292
transform 1 0 53268 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1621523292
transform 1 0 54924 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_579
timestamp 1621523292
transform 1 0 54372 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_588
timestamp 1621523292
transform 1 0 55200 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1621523292
transform 1 0 56856 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1598_
timestamp 1621523292
transform 1 0 55568 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1621523292
transform 1 0 56212 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_595
timestamp 1621523292
transform 1 0 55844 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_600
timestamp 1621523292
transform 1 0 56304 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_609
timestamp 1621523292
transform 1 0 57132 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2315_
timestamp 1621523292
transform 1 0 57500 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1621523292
transform -1 0 58880 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_621
timestamp 1621523292
transform 1 0 58236 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1621523292
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1621523292
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1621523292
transform 1 0 1380 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_6
timestamp 1621523292
transform 1 0 1656 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_18
timestamp 1621523292
transform 1 0 2760 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1621523292
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1621523292
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1621523292
transform 1 0 3772 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_30
timestamp 1621523292
transform 1 0 3864 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_42
timestamp 1621523292
transform 1 0 4968 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1621523292
transform 1 0 3588 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_30
timestamp 1621523292
transform 1 0 3864 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_42
timestamp 1621523292
transform 1 0 4968 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1621523292
transform 1 0 6348 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_54
timestamp 1621523292
transform 1 0 6072 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_58
timestamp 1621523292
transform 1 0 6440 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_54
timestamp 1621523292
transform 1 0 6072 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1621523292
transform 1 0 9016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_70
timestamp 1621523292
transform 1 0 7544 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_82
timestamp 1621523292
transform 1 0 8648 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_66
timestamp 1621523292
transform 1 0 7176 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_78
timestamp 1621523292
transform 1 0 8280 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_87
timestamp 1621523292
transform 1 0 9108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_94
timestamp 1621523292
transform 1 0 9752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_106
timestamp 1621523292
transform 1 0 10856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_99
timestamp 1621523292
transform 1 0 10212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1621523292
transform 1 0 11592 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_115
timestamp 1621523292
transform 1 0 11684 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_127
timestamp 1621523292
transform 1 0 12788 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_111
timestamp 1621523292
transform 1 0 11316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_123
timestamp 1621523292
transform 1 0 12420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1621523292
transform 1 0 14260 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_139
timestamp 1621523292
transform 1 0 13892 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1621523292
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_135
timestamp 1621523292
transform 1 0 13524 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_144
timestamp 1621523292
transform 1 0 14352 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1621523292
transform 1 0 16836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_163
timestamp 1621523292
transform 1 0 16100 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_172
timestamp 1621523292
transform 1 0 16928 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_156
timestamp 1621523292
transform 1 0 15456 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_168
timestamp 1621523292
transform 1 0 16560 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 17664 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_183
timestamp 1621523292
transform 1 0 17940 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_195
timestamp 1621523292
transform 1 0 19044 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_180
timestamp 1621523292
transform 1 0 17664 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_192
timestamp 1621523292
transform 1 0 18768 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1621523292
transform 1 0 19504 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_wb_clk_i
timestamp 1621523292
transform 1 0 19964 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_207
timestamp 1621523292
transform 1 0 20148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_201
timestamp 1621523292
transform 1 0 19596 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_208
timestamp 1621523292
transform 1 0 20240 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1621523292
transform 1 0 22080 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_wb_clk_i
timestamp 1621523292
transform 1 0 22540 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_219
timestamp 1621523292
transform 1 0 21252 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_227
timestamp 1621523292
transform 1 0 21988 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_229
timestamp 1621523292
transform 1 0 22172 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_236
timestamp 1621523292
transform 1 0 22816 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_220
timestamp 1621523292
transform 1 0 21344 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_232
timestamp 1621523292
transform 1 0 22448 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1621523292
transform 1 0 24748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_248
timestamp 1621523292
transform 1 0 23920 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_260
timestamp 1621523292
transform 1 0 25024 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_244
timestamp 1621523292
transform 1 0 23552 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_256
timestamp 1621523292
transform 1 0 24656 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1621523292
transform 1 0 24840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_272
timestamp 1621523292
transform 1 0 26128 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_270
timestamp 1621523292
transform 1 0 25944 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_282
timestamp 1621523292
transform 1 0 27048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1621523292
transform 1 0 27324 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_284
timestamp 1621523292
transform 1 0 27232 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_286
timestamp 1621523292
transform 1 0 27416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_298
timestamp 1621523292
transform 1 0 28520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_294
timestamp 1621523292
transform 1 0 28152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1911_
timestamp 1621523292
transform 1 0 30820 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2389_
timestamp 1621523292
transform 1 0 30452 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1621523292
transform 1 0 29992 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_310
timestamp 1621523292
transform 1 0 29624 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_322
timestamp 1621523292
transform 1 0 30728 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_306
timestamp 1621523292
transform 1 0 29256 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_315
timestamp 1621523292
transform 1 0 30084 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_335
timestamp 1621523292
transform 1 0 31924 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_336
timestamp 1621523292
transform 1 0 32016 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_329
timestamp 1621523292
transform 1 0 31372 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1909_
timestamp 1621523292
transform 1 0 31740 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_345
timestamp 1621523292
transform 1 0 32844 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_343
timestamp 1621523292
transform 1 0 32660 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1621523292
transform 1 0 32568 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1932_
timestamp 1621523292
transform 1 0 32292 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1928_
timestamp 1621523292
transform 1 0 33028 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__or3_4  _1930_
timestamp 1621523292
transform 1 0 33212 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1926_
timestamp 1621523292
transform 1 0 34040 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1927_
timestamp 1621523292
transform 1 0 34684 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1929_
timestamp 1621523292
transform 1 0 34408 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1621523292
transform 1 0 35236 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1621523292
transform 1 0 33672 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1621523292
transform 1 0 34316 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_368
timestamp 1621523292
transform 1 0 34960 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_358
timestamp 1621523292
transform 1 0 34040 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_365
timestamp 1621523292
transform 1 0 34684 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_380
timestamp 1621523292
transform 1 0 36064 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_392
timestamp 1621523292
transform 1 0 37168 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1621523292
transform 1 0 35328 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_384
timestamp 1621523292
transform 1 0 36432 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1621523292
transform 1 0 37812 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_398
timestamp 1621523292
transform 1 0 37720 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_400
timestamp 1621523292
transform 1 0 37904 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_412
timestamp 1621523292
transform 1 0 39008 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_396
timestamp 1621523292
transform 1 0 37536 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_408
timestamp 1621523292
transform 1 0 38640 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1621523292
transform 1 0 40480 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_424
timestamp 1621523292
transform 1 0 40112 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_436
timestamp 1621523292
transform 1 0 41216 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_420
timestamp 1621523292
transform 1 0 39744 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_429
timestamp 1621523292
transform 1 0 40572 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1621523292
transform 1 0 43056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_448
timestamp 1621523292
transform 1 0 42320 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_457
timestamp 1621523292
transform 1 0 43148 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_441
timestamp 1621523292
transform 1 0 41676 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_453
timestamp 1621523292
transform 1 0 42780 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_469
timestamp 1621523292
transform 1 0 44252 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_465
timestamp 1621523292
transform 1 0 43884 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_477
timestamp 1621523292
transform 1 0 44988 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1621523292
transform 1 0 45724 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_481
timestamp 1621523292
transform 1 0 45356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_493
timestamp 1621523292
transform 1 0 46460 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_486
timestamp 1621523292
transform 1 0 45816 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_498
timestamp 1621523292
transform 1 0 46920 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1621523292
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1621523292
transform 1 0 47564 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_514
timestamp 1621523292
transform 1 0 48392 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_510
timestamp 1621523292
transform 1 0 48024 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_522
timestamp 1621523292
transform 1 0 49128 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1621523292
transform 1 0 50968 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_526
timestamp 1621523292
transform 1 0 49496 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_538
timestamp 1621523292
transform 1 0 50600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_534
timestamp 1621523292
transform 1 0 50232 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_543
timestamp 1621523292
transform 1 0 51060 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1621523292
transform 1 0 51704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_562
timestamp 1621523292
transform 1 0 52808 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_555
timestamp 1621523292
transform 1 0 52164 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_567
timestamp 1621523292
transform 1 0 53268 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1621523292
transform 1 0 53544 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1621523292
transform 1 0 55292 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_571
timestamp 1621523292
transform 1 0 53636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_583
timestamp 1621523292
transform 1 0 54740 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_579
timestamp 1621523292
transform 1 0 54372 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_591
timestamp 1621523292
transform 1 0 55476 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_592
timestamp 1621523292
transform 1 0 55568 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2166_
timestamp 1621523292
transform 1 0 55936 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_600
timestamp 1621523292
transform 1 0 56304 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_606
timestamp 1621523292
transform 1 0 56856 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_599
timestamp 1621523292
transform 1 0 56212 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1621523292
transform 1 0 56212 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2165_
timestamp 1621523292
transform 1 0 56580 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_60_608
timestamp 1621523292
transform 1 0 57040 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _1563_
timestamp 1621523292
transform 1 0 57224 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1561_
timestamp 1621523292
transform 1 0 57224 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1621523292
transform -1 0 58880 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1621523292
transform -1 0 58880 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output190
timestamp 1621523292
transform 1 0 57868 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output229
timestamp 1621523292
transform 1 0 57868 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_613
timestamp 1621523292
transform 1 0 57500 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_621
timestamp 1621523292
transform 1 0 58236 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1621523292
transform 1 0 57500 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1621523292
transform 1 0 58236 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1621523292
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1621523292
transform 1 0 1380 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_6
timestamp 1621523292
transform 1 0 1656 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_18
timestamp 1621523292
transform 1 0 2760 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_30
timestamp 1621523292
transform 1 0 3864 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_42
timestamp 1621523292
transform 1 0 4968 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1621523292
transform 1 0 6348 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_54
timestamp 1621523292
transform 1 0 6072 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_58
timestamp 1621523292
transform 1 0 6440 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_70
timestamp 1621523292
transform 1 0 7544 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_82
timestamp 1621523292
transform 1 0 8648 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_94
timestamp 1621523292
transform 1 0 9752 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_106
timestamp 1621523292
transform 1 0 10856 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1621523292
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_115
timestamp 1621523292
transform 1 0 11684 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_127
timestamp 1621523292
transform 1 0 12788 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_139
timestamp 1621523292
transform 1 0 13892 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_151
timestamp 1621523292
transform 1 0 14996 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1621523292
transform 1 0 16836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_163
timestamp 1621523292
transform 1 0 16100 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_172
timestamp 1621523292
transform 1 0 16928 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1997_
timestamp 1621523292
transform 1 0 17480 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_wb_clk_i
timestamp 1621523292
transform 1 0 18124 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_181
timestamp 1621523292
transform 1 0 17756 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_188
timestamp 1621523292
transform 1 0 18400 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_200
timestamp 1621523292
transform 1 0 19504 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_212
timestamp 1621523292
transform 1 0 20608 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1621523292
transform 1 0 22080 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_224
timestamp 1621523292
transform 1 0 21712 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_229
timestamp 1621523292
transform 1 0 22172 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_241
timestamp 1621523292
transform 1 0 23276 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_253
timestamp 1621523292
transform 1 0 24380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_265
timestamp 1621523292
transform 1 0 25484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_277
timestamp 1621523292
transform 1 0 26588 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1621523292
transform 1 0 27324 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1621523292
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_298
timestamp 1621523292
transform 1 0 28520 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1908_
timestamp 1621523292
transform 1 0 30728 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_310
timestamp 1621523292
transform 1 0 29624 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1907_
timestamp 1621523292
transform 1 0 31648 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2396_
timestamp 1621523292
transform 1 0 33120 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1621523292
transform 1 0 32568 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_328
timestamp 1621523292
transform 1 0 31280 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_335
timestamp 1621523292
transform 1 0 31924 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_341
timestamp 1621523292
transform 1 0 32476 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_343
timestamp 1621523292
transform 1 0 32660 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_347
timestamp 1621523292
transform 1 0 33028 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _1933_
timestamp 1621523292
transform 1 0 34960 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_364
timestamp 1621523292
transform 1 0 34592 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_371
timestamp 1621523292
transform 1 0 35236 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_383
timestamp 1621523292
transform 1 0 36340 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1621523292
transform 1 0 37812 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1621523292
transform 1 0 37444 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_400
timestamp 1621523292
transform 1 0 37904 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_412
timestamp 1621523292
transform 1 0 39008 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_424
timestamp 1621523292
transform 1 0 40112 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_436
timestamp 1621523292
transform 1 0 41216 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1621523292
transform 1 0 43056 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_448
timestamp 1621523292
transform 1 0 42320 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_457
timestamp 1621523292
transform 1 0 43148 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_469
timestamp 1621523292
transform 1 0 44252 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_481
timestamp 1621523292
transform 1 0 45356 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_493
timestamp 1621523292
transform 1 0 46460 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1621523292
transform 1 0 48300 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_505
timestamp 1621523292
transform 1 0 47564 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_514
timestamp 1621523292
transform 1 0 48392 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_526
timestamp 1621523292
transform 1 0 49496 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_538
timestamp 1621523292
transform 1 0 50600 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_550
timestamp 1621523292
transform 1 0 51704 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_562
timestamp 1621523292
transform 1 0 52808 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1621523292
transform 1 0 53544 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_571
timestamp 1621523292
transform 1 0 53636 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_583
timestamp 1621523292
transform 1 0 54740 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2167_
timestamp 1621523292
transform 1 0 56856 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1621523292
transform 1 0 56212 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_595
timestamp 1621523292
transform 1 0 55844 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_602
timestamp 1621523292
transform 1 0 56488 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_609
timestamp 1621523292
transform 1 0 57132 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2316_
timestamp 1621523292
transform 1 0 57500 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1621523292
transform -1 0 58880 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_621
timestamp 1621523292
transform 1 0 58236 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1621523292
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1621523292
transform 1 0 1380 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_6
timestamp 1621523292
transform 1 0 1656 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_18
timestamp 1621523292
transform 1 0 2760 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1621523292
transform 1 0 3772 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_26
timestamp 1621523292
transform 1 0 3496 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_30
timestamp 1621523292
transform 1 0 3864 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_42
timestamp 1621523292
transform 1 0 4968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_54
timestamp 1621523292
transform 1 0 6072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1621523292
transform 1 0 9016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_66
timestamp 1621523292
transform 1 0 7176 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_78
timestamp 1621523292
transform 1 0 8280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_87
timestamp 1621523292
transform 1 0 9108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_99
timestamp 1621523292
transform 1 0 10212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_111
timestamp 1621523292
transform 1 0 11316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_123
timestamp 1621523292
transform 1 0 12420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1621523292
transform 1 0 14260 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_135
timestamp 1621523292
transform 1 0 13524 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_144
timestamp 1621523292
transform 1 0 14352 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2421_
timestamp 1621523292
transform 1 0 15640 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_62_156
timestamp 1621523292
transform 1 0 15456 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_174
timestamp 1621523292
transform 1 0 17112 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1996_
timestamp 1621523292
transform 1 0 17480 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1999_
timestamp 1621523292
transform 1 0 18400 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_184
timestamp 1621523292
transform 1 0 18032 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_194
timestamp 1621523292
transform 1 0 18952 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1621523292
transform 1 0 19504 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_201
timestamp 1621523292
transform 1 0 19596 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_213
timestamp 1621523292
transform 1 0 20700 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1621523292
transform 1 0 21804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1621523292
transform 1 0 22908 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1621523292
transform 1 0 24748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_249
timestamp 1621523292
transform 1 0 24012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1621523292
transform 1 0 24840 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_270
timestamp 1621523292
transform 1 0 25944 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_282
timestamp 1621523292
transform 1 0 27048 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2387_
timestamp 1621523292
transform 1 0 27232 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1621523292
transform 1 0 28704 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1906_
timestamp 1621523292
transform 1 0 30452 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1621523292
transform 1 0 29992 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_312
timestamp 1621523292
transform 1 0 29808 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_315
timestamp 1621523292
transform 1 0 30084 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_322
timestamp 1621523292
transform 1 0 30728 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _1935_
timestamp 1621523292
transform 1 0 32200 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1937_
timestamp 1621523292
transform 1 0 33212 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_334
timestamp 1621523292
transform 1 0 31832 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_345
timestamp 1621523292
transform 1 0 32844 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1931_
timestamp 1621523292
transform 1 0 34132 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1621523292
transform 1 0 35236 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_355
timestamp 1621523292
transform 1 0 33764 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_362
timestamp 1621523292
transform 1 0 34408 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_370
timestamp 1621523292
transform 1 0 35144 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_372
timestamp 1621523292
transform 1 0 35328 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_384
timestamp 1621523292
transform 1 0 36432 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_396
timestamp 1621523292
transform 1 0 37536 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_408
timestamp 1621523292
transform 1 0 38640 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1621523292
transform 1 0 40480 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_420
timestamp 1621523292
transform 1 0 39744 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_429
timestamp 1621523292
transform 1 0 40572 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_441
timestamp 1621523292
transform 1 0 41676 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_453
timestamp 1621523292
transform 1 0 42780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_465
timestamp 1621523292
transform 1 0 43884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1621523292
transform 1 0 44988 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1621523292
transform 1 0 45724 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_486
timestamp 1621523292
transform 1 0 45816 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_498
timestamp 1621523292
transform 1 0 46920 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_510
timestamp 1621523292
transform 1 0 48024 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_522
timestamp 1621523292
transform 1 0 49128 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1621523292
transform 1 0 50968 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_534
timestamp 1621523292
transform 1 0 50232 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_543
timestamp 1621523292
transform 1 0 51060 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_555
timestamp 1621523292
transform 1 0 52164 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_567
timestamp 1621523292
transform 1 0 53268 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_579
timestamp 1621523292
transform 1 0 54372 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1560_
timestamp 1621523292
transform 1 0 57224 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1621523292
transform 1 0 56212 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_591
timestamp 1621523292
transform 1 0 55476 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_600
timestamp 1621523292
transform 1 0 56304 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_608
timestamp 1621523292
transform 1 0 57040 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1621523292
transform -1 0 58880 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output191
timestamp 1621523292
transform 1 0 57868 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1621523292
transform 1 0 57500 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1621523292
transform 1 0 58236 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1621523292
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1621523292
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1621523292
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1621523292
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1621523292
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1621523292
transform 1 0 6348 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_51
timestamp 1621523292
transform 1 0 5796 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_58
timestamp 1621523292
transform 1 0 6440 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_70
timestamp 1621523292
transform 1 0 7544 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_82
timestamp 1621523292
transform 1 0 8648 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_94
timestamp 1621523292
transform 1 0 9752 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_106
timestamp 1621523292
transform 1 0 10856 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1621523292
transform 1 0 11592 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_115
timestamp 1621523292
transform 1 0 11684 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_127
timestamp 1621523292
transform 1 0 12788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2420_
timestamp 1621523292
transform 1 0 13892 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1992_
timestamp 1621523292
transform 1 0 15732 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1621523292
transform 1 0 16836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_155
timestamp 1621523292
transform 1 0 15364 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_162
timestamp 1621523292
transform 1 0 16008 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_170
timestamp 1621523292
transform 1 0 16744 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_172
timestamp 1621523292
transform 1 0 16928 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2422_
timestamp 1621523292
transform 1 0 17572 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_63_178
timestamp 1621523292
transform 1 0 17480 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_195
timestamp 1621523292
transform 1 0 19044 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_207
timestamp 1621523292
transform 1 0 20148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1621523292
transform 1 0 22080 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_219
timestamp 1621523292
transform 1 0 21252 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_227
timestamp 1621523292
transform 1 0 21988 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_229
timestamp 1621523292
transform 1 0 22172 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_241
timestamp 1621523292
transform 1 0 23276 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_253
timestamp 1621523292
transform 1 0 24380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_265
timestamp 1621523292
transform 1 0 25484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_277
timestamp 1621523292
transform 1 0 26588 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1902_
timestamp 1621523292
transform 1 0 27876 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2388_
timestamp 1621523292
transform 1 0 28980 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1621523292
transform 1 0 27324 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_286
timestamp 1621523292
transform 1 0 27416 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_290
timestamp 1621523292
transform 1 0 27784 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_297
timestamp 1621523292
transform 1 0 28428 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1905_
timestamp 1621523292
transform 1 0 30820 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_319
timestamp 1621523292
transform 1 0 30452 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1934_
timestamp 1621523292
transform 1 0 31924 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1938_
timestamp 1621523292
transform 1 0 33120 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1621523292
transform 1 0 32568 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1621523292
transform 1 0 31372 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_338
timestamp 1621523292
transform 1 0 32200 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_343
timestamp 1621523292
transform 1 0 32660 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_347
timestamp 1621523292
transform 1 0 33028 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_357
timestamp 1621523292
transform 1 0 33948 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_369
timestamp 1621523292
transform 1 0 35052 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_381
timestamp 1621523292
transform 1 0 36156 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_393
timestamp 1621523292
transform 1 0 37260 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1621523292
transform 1 0 37812 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_400
timestamp 1621523292
transform 1 0 37904 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_412
timestamp 1621523292
transform 1 0 39008 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_424
timestamp 1621523292
transform 1 0 40112 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_436
timestamp 1621523292
transform 1 0 41216 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1621523292
transform 1 0 43056 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_448
timestamp 1621523292
transform 1 0 42320 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_457
timestamp 1621523292
transform 1 0 43148 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_469
timestamp 1621523292
transform 1 0 44252 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_481
timestamp 1621523292
transform 1 0 45356 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_493
timestamp 1621523292
transform 1 0 46460 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1621523292
transform 1 0 48300 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_505
timestamp 1621523292
transform 1 0 47564 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_514
timestamp 1621523292
transform 1 0 48392 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_526
timestamp 1621523292
transform 1 0 49496 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_538
timestamp 1621523292
transform 1 0 50600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_550
timestamp 1621523292
transform 1 0 51704 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_562
timestamp 1621523292
transform 1 0 52808 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1621523292
transform 1 0 53544 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_571
timestamp 1621523292
transform 1 0 53636 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_583
timestamp 1621523292
transform 1 0 54740 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2168_
timestamp 1621523292
transform 1 0 56120 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output230
timestamp 1621523292
transform 1 0 56764 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_595
timestamp 1621523292
transform 1 0 55844 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_601
timestamp 1621523292
transform 1 0 56396 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_609
timestamp 1621523292
transform 1 0 57132 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2317_
timestamp 1621523292
transform 1 0 57500 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1621523292
transform -1 0 58880 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_621
timestamp 1621523292
transform 1 0 58236 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1621523292
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 1621523292
transform 1 0 1380 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_6
timestamp 1621523292
transform 1 0 1656 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_18
timestamp 1621523292
transform 1 0 2760 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1621523292
transform 1 0 3772 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_26
timestamp 1621523292
transform 1 0 3496 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_30
timestamp 1621523292
transform 1 0 3864 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_42
timestamp 1621523292
transform 1 0 4968 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_54
timestamp 1621523292
transform 1 0 6072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1621523292
transform 1 0 9016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_66
timestamp 1621523292
transform 1 0 7176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_78
timestamp 1621523292
transform 1 0 8280 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_87
timestamp 1621523292
transform 1 0 9108 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_99
timestamp 1621523292
transform 1 0 10212 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_111
timestamp 1621523292
transform 1 0 11316 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_123
timestamp 1621523292
transform 1 0 12420 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1993_
timestamp 1621523292
transform 1 0 14720 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1621523292
transform 1 0 14260 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_135
timestamp 1621523292
transform 1 0 13524 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_144
timestamp 1621523292
transform 1 0 14352 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1991_
timestamp 1621523292
transform 1 0 15640 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1994_
timestamp 1621523292
transform 1 0 16284 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1995_
timestamp 1621523292
transform 1 0 16928 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_154
timestamp 1621523292
transform 1 0 15272 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_161
timestamp 1621523292
transform 1 0 15916 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_168
timestamp 1621523292
transform 1 0 16560 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1998_
timestamp 1621523292
transform 1 0 18032 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2000_
timestamp 1621523292
transform 1 0 18676 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_175
timestamp 1621523292
transform 1 0 17204 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_183
timestamp 1621523292
transform 1 0 17940 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_187
timestamp 1621523292
transform 1 0 18308 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_194
timestamp 1621523292
transform 1 0 18952 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2005_
timestamp 1621523292
transform 1 0 19964 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1621523292
transform 1 0 19504 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_wb_clk_i
timestamp 1621523292
transform 1 0 20608 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_201
timestamp 1621523292
transform 1 0 19596 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1621523292
transform 1 0 20240 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1621523292
transform 1 0 20884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_227
timestamp 1621523292
transform 1 0 21988 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1621523292
transform 1 0 23092 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1621523292
transform 1 0 24748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_251
timestamp 1621523292
transform 1 0 24196 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_258
timestamp 1621523292
transform 1 0 24840 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_270
timestamp 1621523292
transform 1 0 25944 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_282
timestamp 1621523292
transform 1 0 27048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1621523292
transform 1 0 28336 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1903_
timestamp 1621523292
transform 1 0 28980 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_294
timestamp 1621523292
transform 1 0 28152 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1621523292
transform 1 0 28612 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1904_
timestamp 1621523292
transform 1 0 30452 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2397_
timestamp 1621523292
transform 1 0 31096 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1621523292
transform 1 0 29992 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_306
timestamp 1621523292
transform 1 0 29256 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_315
timestamp 1621523292
transform 1 0 30084 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_322
timestamp 1621523292
transform 1 0 30728 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_342
timestamp 1621523292
transform 1 0 32568 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2398_
timestamp 1621523292
transform 1 0 33396 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1621523292
transform 1 0 35236 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_350
timestamp 1621523292
transform 1 0 33304 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_367
timestamp 1621523292
transform 1 0 34868 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_372
timestamp 1621523292
transform 1 0 35328 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_384
timestamp 1621523292
transform 1 0 36432 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_396
timestamp 1621523292
transform 1 0 37536 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_408
timestamp 1621523292
transform 1 0 38640 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1621523292
transform 1 0 40480 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_420
timestamp 1621523292
transform 1 0 39744 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_429
timestamp 1621523292
transform 1 0 40572 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_441
timestamp 1621523292
transform 1 0 41676 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_453
timestamp 1621523292
transform 1 0 42780 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_465
timestamp 1621523292
transform 1 0 43884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_477
timestamp 1621523292
transform 1 0 44988 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1621523292
transform 1 0 45724 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_486
timestamp 1621523292
transform 1 0 45816 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_498
timestamp 1621523292
transform 1 0 46920 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_510
timestamp 1621523292
transform 1 0 48024 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_522
timestamp 1621523292
transform 1 0 49128 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1621523292
transform 1 0 50968 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_534
timestamp 1621523292
transform 1 0 50232 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_543
timestamp 1621523292
transform 1 0 51060 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_555
timestamp 1621523292
transform 1 0 52164 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_567
timestamp 1621523292
transform 1 0 53268 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_579
timestamp 1621523292
transform 1 0 54372 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1558_
timestamp 1621523292
transform 1 0 57224 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1621523292
transform 1 0 56212 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_591
timestamp 1621523292
transform 1 0 55476 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_600
timestamp 1621523292
transform 1 0 56304 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_608
timestamp 1621523292
transform 1 0 57040 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1621523292
transform -1 0 58880 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output192
timestamp 1621523292
transform 1 0 57868 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_613
timestamp 1621523292
transform 1 0 57500 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_621
timestamp 1621523292
transform 1 0 58236 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1621523292
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1621523292
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1621523292
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1621523292
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1621523292
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1621523292
transform 1 0 6348 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_51
timestamp 1621523292
transform 1 0 5796 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_58
timestamp 1621523292
transform 1 0 6440 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_70
timestamp 1621523292
transform 1 0 7544 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_82
timestamp 1621523292
transform 1 0 8648 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_94
timestamp 1621523292
transform 1 0 9752 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_106
timestamp 1621523292
transform 1 0 10856 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1621523292
transform 1 0 11592 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_115
timestamp 1621523292
transform 1 0 11684 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_127
timestamp 1621523292
transform 1 0 12788 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2419_
timestamp 1621523292
transform 1 0 13708 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_65_135
timestamp 1621523292
transform 1 0 13524 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _1989_
timestamp 1621523292
transform 1 0 15548 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1621523292
transform 1 0 16836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_wb_clk_i
timestamp 1621523292
transform 1 0 16192 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_153
timestamp 1621523292
transform 1 0 15180 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_160
timestamp 1621523292
transform 1 0 15824 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_167
timestamp 1621523292
transform 1 0 16468 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_172
timestamp 1621523292
transform 1 0 16928 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _2001_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 17296 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2003_
timestamp 1621523292
transform 1 0 18400 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_184
timestamp 1621523292
transform 1 0 18032 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_192
timestamp 1621523292
transform 1 0 18768 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 19688 0 1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_65_200
timestamp 1621523292
transform 1 0 19504 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1621523292
transform 1 0 22080 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_222
timestamp 1621523292
transform 1 0 21528 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_229
timestamp 1621523292
transform 1 0 22172 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_241
timestamp 1621523292
transform 1 0 23276 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_253
timestamp 1621523292
transform 1 0 24380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_265
timestamp 1621523292
transform 1 0 25484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_277
timestamp 1621523292
transform 1 0 26588 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1897_
timestamp 1621523292
transform 1 0 27784 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1900_
timestamp 1621523292
transform 1 0 28888 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1621523292
transform 1 0 27324 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_286
timestamp 1621523292
transform 1 0 27416 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_298
timestamp 1621523292
transform 1 0 28520 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_305
timestamp 1621523292
transform 1 0 29164 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_317
timestamp 1621523292
transform 1 0 30268 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2b_1  _1939_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 33120 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1621523292
transform 1 0 32568 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_329
timestamp 1621523292
transform 1 0 31372 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_341
timestamp 1621523292
transform 1 0 32476 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_343
timestamp 1621523292
transform 1 0 32660 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_347
timestamp 1621523292
transform 1 0 33028 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1936_
timestamp 1621523292
transform 1 0 34408 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1940_
timestamp 1621523292
transform 1 0 35052 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_353
timestamp 1621523292
transform 1 0 33580 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_361
timestamp 1621523292
transform 1 0 34316 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_365
timestamp 1621523292
transform 1 0 34684 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_372
timestamp 1621523292
transform 1 0 35328 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_384
timestamp 1621523292
transform 1 0 36432 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1621523292
transform 1 0 37812 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_396
timestamp 1621523292
transform 1 0 37536 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_400
timestamp 1621523292
transform 1 0 37904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_412
timestamp 1621523292
transform 1 0 39008 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_424
timestamp 1621523292
transform 1 0 40112 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_436
timestamp 1621523292
transform 1 0 41216 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1621523292
transform 1 0 43056 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_448
timestamp 1621523292
transform 1 0 42320 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_457
timestamp 1621523292
transform 1 0 43148 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_469
timestamp 1621523292
transform 1 0 44252 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_481
timestamp 1621523292
transform 1 0 45356 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_493
timestamp 1621523292
transform 1 0 46460 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1621523292
transform 1 0 48300 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_505
timestamp 1621523292
transform 1 0 47564 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_514
timestamp 1621523292
transform 1 0 48392 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_526
timestamp 1621523292
transform 1 0 49496 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_538
timestamp 1621523292
transform 1 0 50600 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_550
timestamp 1621523292
transform 1 0 51704 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_562
timestamp 1621523292
transform 1 0 52808 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1621523292
transform 1 0 53544 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_571
timestamp 1621523292
transform 1 0 53636 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_583
timestamp 1621523292
transform 1 0 54740 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1559_
timestamp 1621523292
transform 1 0 57224 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1621523292
transform 1 0 56580 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_595
timestamp 1621523292
transform 1 0 55844 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_606
timestamp 1621523292
transform 1 0 56856 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1621523292
transform -1 0 58880 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output231
timestamp 1621523292
transform 1 0 57868 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_613
timestamp 1621523292
transform 1 0 57500 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1621523292
transform 1 0 58236 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1621523292
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1621523292
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1621523292
transform 1 0 1380 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1621523292
transform 1 0 1380 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_6
timestamp 1621523292
transform 1 0 1656 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_18
timestamp 1621523292
transform 1 0 2760 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_6
timestamp 1621523292
transform 1 0 1656 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_18
timestamp 1621523292
transform 1 0 2760 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1621523292
transform 1 0 3772 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_26
timestamp 1621523292
transform 1 0 3496 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_30
timestamp 1621523292
transform 1 0 3864 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_42
timestamp 1621523292
transform 1 0 4968 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_30
timestamp 1621523292
transform 1 0 3864 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_42
timestamp 1621523292
transform 1 0 4968 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1621523292
transform 1 0 6348 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_54
timestamp 1621523292
transform 1 0 6072 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_54
timestamp 1621523292
transform 1 0 6072 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_58
timestamp 1621523292
transform 1 0 6440 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1621523292
transform 1 0 9016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_66
timestamp 1621523292
transform 1 0 7176 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_78
timestamp 1621523292
transform 1 0 8280 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_87
timestamp 1621523292
transform 1 0 9108 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_70
timestamp 1621523292
transform 1 0 7544 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_82
timestamp 1621523292
transform 1 0 8648 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_99
timestamp 1621523292
transform 1 0 10212 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_94
timestamp 1621523292
transform 1 0 9752 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_106
timestamp 1621523292
transform 1 0 10856 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1718_
timestamp 1621523292
transform 1 0 12420 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2415_
timestamp 1621523292
transform 1 0 11868 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1621523292
transform 1 0 11592 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_111
timestamp 1621523292
transform 1 0 11316 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_115
timestamp 1621523292
transform 1 0 11684 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_126
timestamp 1621523292
transform 1 0 12696 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1984_
timestamp 1621523292
transform 1 0 13340 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1986_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 14720 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1990_
timestamp 1621523292
transform 1 0 14720 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1621523292
transform 1 0 14260 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_133
timestamp 1621523292
transform 1 0 13340 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1621523292
transform 1 0 14076 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_144
timestamp 1621523292
transform 1 0 14352 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_132
timestamp 1621523292
transform 1 0 13248 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_136
timestamp 1621523292
transform 1 0 13616 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1987_
timestamp 1621523292
transform 1 0 15548 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2423_
timestamp 1621523292
transform 1 0 15916 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1621523292
transform 1 0 16836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_154
timestamp 1621523292
transform 1 0 15272 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_160
timestamp 1621523292
transform 1 0 15824 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_153
timestamp 1621523292
transform 1 0 15180 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_161
timestamp 1621523292
transform 1 0 15916 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1621523292
transform 1 0 16652 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_172
timestamp 1621523292
transform 1 0 16928 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2002_
timestamp 1621523292
transform 1 0 18032 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2004_
timestamp 1621523292
transform 1 0 18860 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2424_
timestamp 1621523292
transform 1 0 17664 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_66_177
timestamp 1621523292
transform 1 0 17388 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_183
timestamp 1621523292
transform 1 0 17940 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_189
timestamp 1621523292
transform 1 0 18492 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_196
timestamp 1621523292
transform 1 0 19136 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_196
timestamp 1621523292
transform 1 0 19136 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2006_
timestamp 1621523292
transform 1 0 19504 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2007_
timestamp 1621523292
transform 1 0 20424 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2425_
timestamp 1621523292
transform 1 0 19964 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1621523292
transform 1 0 19504 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_201
timestamp 1621523292
transform 1 0 19596 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_206
timestamp 1621523292
transform 1 0 20056 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_213
timestamp 1621523292
transform 1 0 20700 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1621523292
transform 1 0 22080 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_221
timestamp 1621523292
transform 1 0 21436 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_233
timestamp 1621523292
transform 1 0 22540 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_225
timestamp 1621523292
transform 1 0 21804 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_229
timestamp 1621523292
transform 1 0 22172 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2384_
timestamp 1621523292
transform 1 0 24472 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1621523292
transform 1 0 24748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_245
timestamp 1621523292
transform 1 0 23644 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_258
timestamp 1621523292
transform 1 0 24840 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_241
timestamp 1621523292
transform 1 0 23276 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_253
timestamp 1621523292
transform 1 0 24380 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1894_
timestamp 1621523292
transform 1 0 25852 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1895_
timestamp 1621523292
transform 1 0 26312 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2385_
timestamp 1621523292
transform 1 0 26496 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_66_266
timestamp 1621523292
transform 1 0 25576 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_272
timestamp 1621523292
transform 1 0 26128 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_270
timestamp 1621523292
transform 1 0 25944 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_280
timestamp 1621523292
transform 1 0 26864 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1898_
timestamp 1621523292
transform 1 0 28336 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1899_
timestamp 1621523292
transform 1 0 29164 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2386_
timestamp 1621523292
transform 1 0 28336 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1621523292
transform 1 0 27324 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_292
timestamp 1621523292
transform 1 0 27968 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_301
timestamp 1621523292
transform 1 0 28796 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_284
timestamp 1621523292
transform 1 0 27232 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_286
timestamp 1621523292
transform 1 0 27416 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_294
timestamp 1621523292
transform 1 0 28152 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2400_
timestamp 1621523292
transform 1 0 30912 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1621523292
transform 1 0 29992 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1621523292
transform 1 0 29532 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_313
timestamp 1621523292
transform 1 0 29900 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_315
timestamp 1621523292
transform 1 0 30084 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_323
timestamp 1621523292
transform 1 0 30820 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_312
timestamp 1621523292
transform 1 0 29808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_324
timestamp 1621523292
transform 1 0 30912 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1941_
timestamp 1621523292
transform 1 0 33028 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1944_
timestamp 1621523292
transform 1 0 32752 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1945_
timestamp 1621523292
transform 1 0 31648 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1621523292
transform 1 0 32568 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_340
timestamp 1621523292
transform 1 0 32384 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_338
timestamp 1621523292
transform 1 0 32200 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_343
timestamp 1621523292
transform 1 0 32660 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1942_
timestamp 1621523292
transform 1 0 33948 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2399_
timestamp 1621523292
transform 1 0 33672 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1621523292
transform 1 0 35236 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_353
timestamp 1621523292
transform 1 0 33580 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_361
timestamp 1621523292
transform 1 0 34316 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_369
timestamp 1621523292
transform 1 0 35052 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_350
timestamp 1621523292
transform 1 0 33304 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_370
timestamp 1621523292
transform 1 0 35144 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_372
timestamp 1621523292
transform 1 0 35328 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_384
timestamp 1621523292
transform 1 0 36432 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_382
timestamp 1621523292
transform 1 0 36248 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1621523292
transform 1 0 37812 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_396
timestamp 1621523292
transform 1 0 37536 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_408
timestamp 1621523292
transform 1 0 38640 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_394
timestamp 1621523292
transform 1 0 37352 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_398
timestamp 1621523292
transform 1 0 37720 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_400
timestamp 1621523292
transform 1 0 37904 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_412
timestamp 1621523292
transform 1 0 39008 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1621523292
transform 1 0 40480 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_420
timestamp 1621523292
transform 1 0 39744 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_429
timestamp 1621523292
transform 1 0 40572 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_424
timestamp 1621523292
transform 1 0 40112 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_436
timestamp 1621523292
transform 1 0 41216 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1621523292
transform 1 0 43056 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_441
timestamp 1621523292
transform 1 0 41676 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_453
timestamp 1621523292
transform 1 0 42780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_448
timestamp 1621523292
transform 1 0 42320 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_457
timestamp 1621523292
transform 1 0 43148 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_465
timestamp 1621523292
transform 1 0 43884 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_477
timestamp 1621523292
transform 1 0 44988 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_469
timestamp 1621523292
transform 1 0 44252 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1621523292
transform 1 0 45724 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_486
timestamp 1621523292
transform 1 0 45816 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_498
timestamp 1621523292
transform 1 0 46920 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_481
timestamp 1621523292
transform 1 0 45356 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_493
timestamp 1621523292
transform 1 0 46460 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1621523292
transform 1 0 48300 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_510
timestamp 1621523292
transform 1 0 48024 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_522
timestamp 1621523292
transform 1 0 49128 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_505
timestamp 1621523292
transform 1 0 47564 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_514
timestamp 1621523292
transform 1 0 48392 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1621523292
transform 1 0 50968 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_534
timestamp 1621523292
transform 1 0 50232 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_543
timestamp 1621523292
transform 1 0 51060 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_526
timestamp 1621523292
transform 1 0 49496 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_538
timestamp 1621523292
transform 1 0 50600 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_555
timestamp 1621523292
transform 1 0 52164 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_567
timestamp 1621523292
transform 1 0 53268 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_550
timestamp 1621523292
transform 1 0 51704 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_562
timestamp 1621523292
transform 1 0 52808 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1621523292
transform 1 0 53544 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_579
timestamp 1621523292
transform 1 0 54372 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_571
timestamp 1621523292
transform 1 0 53636 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_583
timestamp 1621523292
transform 1 0 54740 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2169_
timestamp 1621523292
transform 1 0 56856 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1621523292
transform 1 0 56212 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_591
timestamp 1621523292
transform 1 0 55476 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_600
timestamp 1621523292
transform 1 0 56304 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_609
timestamp 1621523292
transform 1 0 57132 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_595
timestamp 1621523292
transform 1 0 55844 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_607
timestamp 1621523292
transform 1 0 56948 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2318_
timestamp 1621523292
transform 1 0 57500 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1621523292
transform -1 0 58880 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1621523292
transform -1 0 58880 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output193
timestamp 1621523292
transform 1 0 57868 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_621
timestamp 1621523292
transform 1 0 58236 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_615
timestamp 1621523292
transform 1 0 57684 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1621523292
transform 1 0 58236 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1621523292
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1621523292
transform 1 0 1380 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1621523292
transform 1 0 2484 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1621523292
transform 1 0 3772 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_27
timestamp 1621523292
transform 1 0 3588 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_30
timestamp 1621523292
transform 1 0 3864 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_42
timestamp 1621523292
transform 1 0 4968 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_54
timestamp 1621523292
transform 1 0 6072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1621523292
transform 1 0 9016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_66
timestamp 1621523292
transform 1 0 7176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_78
timestamp 1621523292
transform 1 0 8280 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_87
timestamp 1621523292
transform 1 0 9108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_99
timestamp 1621523292
transform 1 0 10212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2416_
timestamp 1621523292
transform 1 0 11500 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_68_111
timestamp 1621523292
transform 1 0 11316 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_129
timestamp 1621523292
transform 1 0 12972 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1621523292
transform 1 0 13340 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1621523292
transform 1 0 14260 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_136
timestamp 1621523292
transform 1 0 13616 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_142
timestamp 1621523292
transform 1 0 14168 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_144
timestamp 1621523292
transform 1 0 14352 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_152
timestamp 1621523292
transform 1 0 15088 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2418_
timestamp 1621523292
transform 1 0 15180 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_68_169
timestamp 1621523292
transform 1 0 16652 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_wb_clk_i
timestamp 1621523292
transform 1 0 17296 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_175
timestamp 1621523292
transform 1 0 17204 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_179
timestamp 1621523292
transform 1 0 17572 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_191
timestamp 1621523292
transform 1 0 18676 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2010_
timestamp 1621523292
transform 1 0 20148 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2011_
timestamp 1621523292
transform 1 0 20792 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1621523292
transform 1 0 19504 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_199
timestamp 1621523292
transform 1 0 19412 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_201
timestamp 1621523292
transform 1 0 19596 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_210
timestamp 1621523292
transform 1 0 20424 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_217
timestamp 1621523292
transform 1 0 21068 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_229
timestamp 1621523292
transform 1 0 22172 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1621523292
transform 1 0 24748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_241
timestamp 1621523292
transform 1 0 23276 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1621523292
transform 1 0 24380 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_258
timestamp 1621523292
transform 1 0 24840 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2383_
timestamp 1621523292
transform 1 0 25484 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_68_264
timestamp 1621523292
transform 1 0 25392 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_281
timestamp 1621523292
transform 1 0 26956 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1896_
timestamp 1621523292
transform 1 0 27324 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2033_
timestamp 1621523292
transform 1 0 28060 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_288
timestamp 1621523292
transform 1 0 27600 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_292
timestamp 1621523292
transform 1 0 27968 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_296
timestamp 1621523292
transform 1 0 28336 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1947_
timestamp 1621523292
transform 1 0 31188 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1621523292
transform 1 0 29992 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_308
timestamp 1621523292
transform 1 0 29440 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_315
timestamp 1621523292
transform 1 0 30084 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1943_
timestamp 1621523292
transform 1 0 31832 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_2  _1951_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 32476 0 -1 39712
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_68_330
timestamp 1621523292
transform 1 0 31464 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_337
timestamp 1621523292
transform 1 0 32108 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1621523292
transform 1 0 35236 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_351
timestamp 1621523292
transform 1 0 33396 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_363
timestamp 1621523292
transform 1 0 34500 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_372
timestamp 1621523292
transform 1 0 35328 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_384
timestamp 1621523292
transform 1 0 36432 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_396
timestamp 1621523292
transform 1 0 37536 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_408
timestamp 1621523292
transform 1 0 38640 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1621523292
transform 1 0 40480 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_420
timestamp 1621523292
transform 1 0 39744 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_429
timestamp 1621523292
transform 1 0 40572 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_441
timestamp 1621523292
transform 1 0 41676 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_453
timestamp 1621523292
transform 1 0 42780 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_465
timestamp 1621523292
transform 1 0 43884 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_477
timestamp 1621523292
transform 1 0 44988 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1621523292
transform 1 0 45724 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_486
timestamp 1621523292
transform 1 0 45816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_498
timestamp 1621523292
transform 1 0 46920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_510
timestamp 1621523292
transform 1 0 48024 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_522
timestamp 1621523292
transform 1 0 49128 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1621523292
transform 1 0 50968 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_534
timestamp 1621523292
transform 1 0 50232 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_543
timestamp 1621523292
transform 1 0 51060 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_555
timestamp 1621523292
transform 1 0 52164 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_567
timestamp 1621523292
transform 1 0 53268 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_579
timestamp 1621523292
transform 1 0 54372 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1621523292
transform 1 0 56212 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_591
timestamp 1621523292
transform 1 0 55476 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_600
timestamp 1621523292
transform 1 0 56304 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1621523292
transform -1 0 58880 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1621523292
transform 1 0 57960 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_612
timestamp 1621523292
transform 1 0 57408 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_621
timestamp 1621523292
transform 1 0 58236 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1621523292
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1621523292
transform 1 0 1380 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_6
timestamp 1621523292
transform 1 0 1656 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_18
timestamp 1621523292
transform 1 0 2760 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_30
timestamp 1621523292
transform 1 0 3864 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_42
timestamp 1621523292
transform 1 0 4968 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1621523292
transform 1 0 6348 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_54
timestamp 1621523292
transform 1 0 6072 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_58
timestamp 1621523292
transform 1 0 6440 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_70
timestamp 1621523292
transform 1 0 7544 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_82
timestamp 1621523292
transform 1 0 8648 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_94
timestamp 1621523292
transform 1 0 9752 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_106
timestamp 1621523292
transform 1 0 10856 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1983_
timestamp 1621523292
transform 1 0 12236 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1621523292
transform 1 0 11592 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_115
timestamp 1621523292
transform 1 0 11684 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_127
timestamp 1621523292
transform 1 0 12788 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2417_
timestamp 1621523292
transform 1 0 13340 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_149
timestamp 1621523292
transform 1 0 14812 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1985_
timestamp 1621523292
transform 1 0 15180 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1621523292
transform 1 0 16836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_161
timestamp 1621523292
transform 1 0 15916 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_169
timestamp 1621523292
transform 1 0 16652 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_172
timestamp 1621523292
transform 1 0 16928 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2426_
timestamp 1621523292
transform 1 0 18308 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_69_184
timestamp 1621523292
transform 1 0 18032 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2427_
timestamp 1621523292
transform 1 0 20148 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_203
timestamp 1621523292
transform 1 0 19780 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1621523292
transform 1 0 22080 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_223
timestamp 1621523292
transform 1 0 21620 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_227
timestamp 1621523292
transform 1 0 21988 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_229
timestamp 1621523292
transform 1 0 22172 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_241
timestamp 1621523292
transform 1 0 23276 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_253
timestamp 1621523292
transform 1 0 24380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1717_
timestamp 1621523292
transform 1 0 25944 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_265
timestamp 1621523292
transform 1 0 25484 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_269
timestamp 1621523292
transform 1 0 25852 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_273
timestamp 1621523292
transform 1 0 26220 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2436_
timestamp 1621523292
transform 1 0 27784 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1621523292
transform 1 0 27324 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_286
timestamp 1621523292
transform 1 0 27416 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2037_
timestamp 1621523292
transform 1 0 29624 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2401_
timestamp 1621523292
transform 1 0 30452 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_69_306
timestamp 1621523292
transform 1 0 29256 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_313
timestamp 1621523292
transform 1 0 29900 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2402_
timestamp 1621523292
transform 1 0 33028 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1621523292
transform 1 0 32568 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_335
timestamp 1621523292
transform 1 0 31924 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_341
timestamp 1621523292
transform 1 0 32476 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_343
timestamp 1621523292
transform 1 0 32660 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1949_
timestamp 1621523292
transform 1 0 34868 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_363
timestamp 1621523292
transform 1 0 34500 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_370
timestamp 1621523292
transform 1 0 35144 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_382
timestamp 1621523292
transform 1 0 36248 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1621523292
transform 1 0 37812 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_394
timestamp 1621523292
transform 1 0 37352 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_398
timestamp 1621523292
transform 1 0 37720 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_400
timestamp 1621523292
transform 1 0 37904 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_412
timestamp 1621523292
transform 1 0 39008 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_424
timestamp 1621523292
transform 1 0 40112 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_436
timestamp 1621523292
transform 1 0 41216 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1621523292
transform 1 0 43056 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_448
timestamp 1621523292
transform 1 0 42320 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_457
timestamp 1621523292
transform 1 0 43148 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_469
timestamp 1621523292
transform 1 0 44252 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_481
timestamp 1621523292
transform 1 0 45356 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_493
timestamp 1621523292
transform 1 0 46460 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1621523292
transform 1 0 48300 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1621523292
transform 1 0 47564 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_514
timestamp 1621523292
transform 1 0 48392 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_526
timestamp 1621523292
transform 1 0 49496 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_538
timestamp 1621523292
transform 1 0 50600 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_550
timestamp 1621523292
transform 1 0 51704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_562
timestamp 1621523292
transform 1 0 52808 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1621523292
transform 1 0 53544 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_571
timestamp 1621523292
transform 1 0 53636 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_583
timestamp 1621523292
transform 1 0 54740 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2170_
timestamp 1621523292
transform 1 0 57224 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_595
timestamp 1621523292
transform 1 0 55844 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_607
timestamp 1621523292
transform 1 0 56948 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1621523292
transform -1 0 58880 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output232
timestamp 1621523292
transform 1 0 57868 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_613
timestamp 1621523292
transform 1 0 57500 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_621
timestamp 1621523292
transform 1 0 58236 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1621523292
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1621523292
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1621523292
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1621523292
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_27
timestamp 1621523292
transform 1 0 3588 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_30
timestamp 1621523292
transform 1 0 3864 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_42
timestamp 1621523292
transform 1 0 4968 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_54
timestamp 1621523292
transform 1 0 6072 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1621523292
transform 1 0 9016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_66
timestamp 1621523292
transform 1 0 7176 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_78
timestamp 1621523292
transform 1 0 8280 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_87
timestamp 1621523292
transform 1 0 9108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_99
timestamp 1621523292
transform 1 0 10212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_111
timestamp 1621523292
transform 1 0 11316 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_123
timestamp 1621523292
transform 1 0 12420 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1988_
timestamp 1621523292
transform 1 0 15088 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1621523292
transform 1 0 14260 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_135
timestamp 1621523292
transform 1 0 13524 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_144
timestamp 1621523292
transform 1 0 14352 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_155
timestamp 1621523292
transform 1 0 15364 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_167
timestamp 1621523292
transform 1 0 16468 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _2009_
timestamp 1621523292
transform 1 0 18584 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_179
timestamp 1621523292
transform 1 0 17572 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_187
timestamp 1621523292
transform 1 0 18308 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_196
timestamp 1621523292
transform 1 0 19136 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2008_
timestamp 1621523292
transform 1 0 19964 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2012_
timestamp 1621523292
transform 1 0 20608 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1621523292
transform 1 0 19504 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_201
timestamp 1621523292
transform 1 0 19596 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_208
timestamp 1621523292
transform 1 0 20240 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_218
timestamp 1621523292
transform 1 0 21160 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2013_
timestamp 1621523292
transform 1 0 21528 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2014_
timestamp 1621523292
transform 1 0 22172 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_225
timestamp 1621523292
transform 1 0 21804 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_232
timestamp 1621523292
transform 1 0 22448 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _2025_
timestamp 1621523292
transform 1 0 24012 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1621523292
transform 1 0 24748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_244
timestamp 1621523292
transform 1 0 23552 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_248
timestamp 1621523292
transform 1 0 23920 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_252
timestamp 1621523292
transform 1 0 24288 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_256
timestamp 1621523292
transform 1 0 24656 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_258
timestamp 1621523292
transform 1 0 24840 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _2028_
timestamp 1621523292
transform 1 0 25576 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2031_
timestamp 1621523292
transform 1 0 26864 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_271
timestamp 1621523292
transform 1 0 26036 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_279
timestamp 1621523292
transform 1 0 26772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_283
timestamp 1621523292
transform 1 0 27140 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2035_
timestamp 1621523292
transform 1 0 27508 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _2038_
timestamp 1621523292
transform 1 0 28980 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_70_293
timestamp 1621523292
transform 1 0 28060 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_301
timestamp 1621523292
transform 1 0 28796 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _2036_
timestamp 1621523292
transform 1 0 30452 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1621523292
transform 1 0 29992 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_310
timestamp 1621523292
transform 1 0 29624 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_315
timestamp 1621523292
transform 1 0 30084 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_322
timestamp 1621523292
transform 1 0 30728 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1948_
timestamp 1621523292
transform 1 0 31280 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1952_
timestamp 1621523292
transform 1 0 32568 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_70_335
timestamp 1621523292
transform 1 0 31924 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_341
timestamp 1621523292
transform 1 0 32476 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_348
timestamp 1621523292
transform 1 0 33120 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1950_
timestamp 1621523292
transform 1 0 33488 0 -1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1621523292
transform 1 0 35236 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_357
timestamp 1621523292
transform 1 0 33948 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_369
timestamp 1621523292
transform 1 0 35052 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_372
timestamp 1621523292
transform 1 0 35328 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_384
timestamp 1621523292
transform 1 0 36432 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_396
timestamp 1621523292
transform 1 0 37536 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_408
timestamp 1621523292
transform 1 0 38640 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1621523292
transform 1 0 40480 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_420
timestamp 1621523292
transform 1 0 39744 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_429
timestamp 1621523292
transform 1 0 40572 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_441
timestamp 1621523292
transform 1 0 41676 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_453
timestamp 1621523292
transform 1 0 42780 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_465
timestamp 1621523292
transform 1 0 43884 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_477
timestamp 1621523292
transform 1 0 44988 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1621523292
transform 1 0 45724 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_486
timestamp 1621523292
transform 1 0 45816 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_498
timestamp 1621523292
transform 1 0 46920 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_510
timestamp 1621523292
transform 1 0 48024 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_522
timestamp 1621523292
transform 1 0 49128 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1621523292
transform 1 0 50968 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_534
timestamp 1621523292
transform 1 0 50232 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_543
timestamp 1621523292
transform 1 0 51060 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_555
timestamp 1621523292
transform 1 0 52164 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_567
timestamp 1621523292
transform 1 0 53268 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_579
timestamp 1621523292
transform 1 0 54372 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1557_
timestamp 1621523292
transform 1 0 56856 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1621523292
transform 1 0 56212 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_591
timestamp 1621523292
transform 1 0 55476 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_70_600
timestamp 1621523292
transform 1 0 56304 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_609
timestamp 1621523292
transform 1 0 57132 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2319_
timestamp 1621523292
transform 1 0 57500 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1621523292
transform -1 0 58880 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1621523292
transform 1 0 58236 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1621523292
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1621523292
transform 1 0 1380 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_6
timestamp 1621523292
transform 1 0 1656 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1621523292
transform 1 0 2760 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1621523292
transform 1 0 3864 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1621523292
transform 1 0 4968 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1621523292
transform 1 0 6348 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_54
timestamp 1621523292
transform 1 0 6072 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_58
timestamp 1621523292
transform 1 0 6440 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_70
timestamp 1621523292
transform 1 0 7544 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_82
timestamp 1621523292
transform 1 0 8648 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_94
timestamp 1621523292
transform 1 0 9752 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_106
timestamp 1621523292
transform 1 0 10856 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1621523292
transform 1 0 11592 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_115
timestamp 1621523292
transform 1 0 11684 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_127
timestamp 1621523292
transform 1 0 12788 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_139
timestamp 1621523292
transform 1 0 13892 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_151
timestamp 1621523292
transform 1 0 14996 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1621523292
transform 1 0 16836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_163
timestamp 1621523292
transform 1 0 16100 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_172
timestamp 1621523292
transform 1 0 16928 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1621523292
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_196
timestamp 1621523292
transform 1 0 19136 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _2015_
timestamp 1621523292
transform 1 0 21160 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_208
timestamp 1621523292
transform 1 0 20240 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_216
timestamp 1621523292
transform 1 0 20976 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2433_
timestamp 1621523292
transform 1 0 23092 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1621523292
transform 1 0 22080 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_224
timestamp 1621523292
transform 1 0 21712 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_229
timestamp 1621523292
transform 1 0 22172 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_237
timestamp 1621523292
transform 1 0 22908 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2434_
timestamp 1621523292
transform 1 0 24932 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_255
timestamp 1621523292
transform 1 0 24564 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_275
timestamp 1621523292
transform 1 0 26404 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_283
timestamp 1621523292
transform 1 0 27140 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_1  _2032_
timestamp 1621523292
transform 1 0 27784 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2437_
timestamp 1621523292
transform 1 0 28796 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1621523292
transform 1 0 27324 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_286
timestamp 1621523292
transform 1 0 27416 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_294
timestamp 1621523292
transform 1 0 28152 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_300
timestamp 1621523292
transform 1 0 28704 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _2040_
timestamp 1621523292
transform 1 0 30636 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_317
timestamp 1621523292
transform 1 0 30268 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_327
timestamp 1621523292
transform 1 0 31188 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1946_
timestamp 1621523292
transform 1 0 31832 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1953_
timestamp 1621523292
transform 1 0 33028 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1621523292
transform 1 0 32568 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_333
timestamp 1621523292
transform 1 0 31740 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_337
timestamp 1621523292
transform 1 0 32108 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_341
timestamp 1621523292
transform 1 0 32476 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_343
timestamp 1621523292
transform 1 0 32660 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_350
timestamp 1621523292
transform 1 0 33304 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_362
timestamp 1621523292
transform 1 0 34408 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_374
timestamp 1621523292
transform 1 0 35512 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_386
timestamp 1621523292
transform 1 0 36616 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1621523292
transform 1 0 37812 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_398
timestamp 1621523292
transform 1 0 37720 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_400
timestamp 1621523292
transform 1 0 37904 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_412
timestamp 1621523292
transform 1 0 39008 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_424
timestamp 1621523292
transform 1 0 40112 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_436
timestamp 1621523292
transform 1 0 41216 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1621523292
transform 1 0 43056 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_448
timestamp 1621523292
transform 1 0 42320 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_457
timestamp 1621523292
transform 1 0 43148 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_469
timestamp 1621523292
transform 1 0 44252 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_481
timestamp 1621523292
transform 1 0 45356 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_493
timestamp 1621523292
transform 1 0 46460 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1621523292
transform 1 0 48300 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1621523292
transform 1 0 47564 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_514
timestamp 1621523292
transform 1 0 48392 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_526
timestamp 1621523292
transform 1 0 49496 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_538
timestamp 1621523292
transform 1 0 50600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_550
timestamp 1621523292
transform 1 0 51704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_562
timestamp 1621523292
transform 1 0 52808 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1621523292
transform 1 0 53544 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_571
timestamp 1621523292
transform 1 0 53636 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_583
timestamp 1621523292
transform 1 0 54740 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1621523292
transform 1 0 56488 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output233
timestamp 1621523292
transform 1 0 57132 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_595
timestamp 1621523292
transform 1 0 55844 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_601
timestamp 1621523292
transform 1 0 56396 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_605
timestamp 1621523292
transform 1 0 56764 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1621523292
transform -1 0 58880 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output194
timestamp 1621523292
transform 1 0 57868 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_613
timestamp 1621523292
transform 1 0 57500 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_621
timestamp 1621523292
transform 1 0 58236 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1621523292
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1621523292
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1621523292
transform 1 0 1380 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1621523292
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1621523292
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_6
timestamp 1621523292
transform 1 0 1656 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_18
timestamp 1621523292
transform 1 0 2760 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1621523292
transform 1 0 3772 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_27
timestamp 1621523292
transform 1 0 3588 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_30
timestamp 1621523292
transform 1 0 3864 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_42
timestamp 1621523292
transform 1 0 4968 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_30
timestamp 1621523292
transform 1 0 3864 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_42
timestamp 1621523292
transform 1 0 4968 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1621523292
transform 1 0 6348 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_54
timestamp 1621523292
transform 1 0 6072 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_54
timestamp 1621523292
transform 1 0 6072 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_58
timestamp 1621523292
transform 1 0 6440 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1621523292
transform 1 0 9016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_66
timestamp 1621523292
transform 1 0 7176 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_78
timestamp 1621523292
transform 1 0 8280 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_87
timestamp 1621523292
transform 1 0 9108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_70
timestamp 1621523292
transform 1 0 7544 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_82
timestamp 1621523292
transform 1 0 8648 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_99
timestamp 1621523292
transform 1 0 10212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_94
timestamp 1621523292
transform 1 0 9752 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_106
timestamp 1621523292
transform 1 0 10856 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1621523292
transform 1 0 11592 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_111
timestamp 1621523292
transform 1 0 11316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_123
timestamp 1621523292
transform 1 0 12420 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_115
timestamp 1621523292
transform 1 0 11684 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_127
timestamp 1621523292
transform 1 0 12788 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1621523292
transform 1 0 14260 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_135
timestamp 1621523292
transform 1 0 13524 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_144
timestamp 1621523292
transform 1 0 14352 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_139
timestamp 1621523292
transform 1 0 13892 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_151
timestamp 1621523292
transform 1 0 14996 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1621523292
transform 1 0 16836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_156
timestamp 1621523292
transform 1 0 15456 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_168
timestamp 1621523292
transform 1 0 16560 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_163
timestamp 1621523292
transform 1 0 16100 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_172
timestamp 1621523292
transform 1 0 16928 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_180
timestamp 1621523292
transform 1 0 17664 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_192
timestamp 1621523292
transform 1 0 18768 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_184
timestamp 1621523292
transform 1 0 18032 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_196
timestamp 1621523292
transform 1 0 19136 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2016_
timestamp 1621523292
transform 1 0 20792 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2429_
timestamp 1621523292
transform 1 0 19504 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1621523292
transform 1 0 19504 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_201
timestamp 1621523292
transform 1 0 19596 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_213
timestamp 1621523292
transform 1 0 20700 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_217
timestamp 1621523292
transform 1 0 21068 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_216
timestamp 1621523292
transform 1 0 20976 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2019_
timestamp 1621523292
transform 1 0 21344 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2428_
timestamp 1621523292
transform 1 0 21436 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1621523292
transform 1 0 22080 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_237
timestamp 1621523292
transform 1 0 22908 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_224
timestamp 1621523292
transform 1 0 21712 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_229
timestamp 1621523292
transform 1 0 22172 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_241
timestamp 1621523292
transform 1 0 23276 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2026_
timestamp 1621523292
transform 1 0 23644 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2023_
timestamp 1621523292
transform 1 0 23552 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_248
timestamp 1621523292
transform 1 0 23920 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_251
timestamp 1621523292
transform 1 0 24196 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2024_
timestamp 1621523292
transform 1 0 24288 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_255
timestamp 1621523292
transform 1 0 24564 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_258
timestamp 1621523292
transform 1 0 24840 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1621523292
transform 1 0 24748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2027_
timestamp 1621523292
transform 1 0 24932 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_262
timestamp 1621523292
transform 1 0 25208 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_262
timestamp 1621523292
transform 1 0 25208 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _2029_
timestamp 1621523292
transform 1 0 25300 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2051_
timestamp 1621523292
transform 1 0 26496 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2435_
timestamp 1621523292
transform 1 0 26312 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_wb_clk_i
timestamp 1621523292
transform 1 0 25852 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_269
timestamp 1621523292
transform 1 0 25852 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_273
timestamp 1621523292
transform 1 0 26220 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_268
timestamp 1621523292
transform 1 0 25760 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_272
timestamp 1621523292
transform 1 0 26128 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_279
timestamp 1621523292
transform 1 0 26772 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _2034_
timestamp 1621523292
transform 1 0 28152 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _2042_
timestamp 1621523292
transform 1 0 27876 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2438_
timestamp 1621523292
transform 1 0 29072 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1621523292
transform 1 0 27324 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_290
timestamp 1621523292
transform 1 0 27784 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_303
timestamp 1621523292
transform 1 0 28980 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_286
timestamp 1621523292
transform 1 0 27416 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_290
timestamp 1621523292
transform 1 0 27784 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_300
timestamp 1621523292
transform 1 0 28704 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2030_
timestamp 1621523292
transform 1 0 29348 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2403_
timestamp 1621523292
transform 1 0 30636 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1621523292
transform 1 0 29992 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_310
timestamp 1621523292
transform 1 0 29624 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_315
timestamp 1621523292
transform 1 0 30084 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_320
timestamp 1621523292
transform 1 0 30544 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1954_
timestamp 1621523292
transform 1 0 31464 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1955_
timestamp 1621523292
transform 1 0 32476 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2404_
timestamp 1621523292
transform 1 0 33028 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1621523292
transform 1 0 32568 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_337
timestamp 1621523292
transform 1 0 32108 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_346
timestamp 1621523292
transform 1 0 32936 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_328
timestamp 1621523292
transform 1 0 31280 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_338
timestamp 1621523292
transform 1 0 32200 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_343
timestamp 1621523292
transform 1 0 32660 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1956_
timestamp 1621523292
transform 1 0 33304 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1621523292
transform 1 0 35236 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_354
timestamp 1621523292
transform 1 0 33672 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_366
timestamp 1621523292
transform 1 0 34776 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_370
timestamp 1621523292
transform 1 0 35144 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_363
timestamp 1621523292
transform 1 0 34500 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_372
timestamp 1621523292
transform 1 0 35328 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_384
timestamp 1621523292
transform 1 0 36432 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_375
timestamp 1621523292
transform 1 0 35604 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_387
timestamp 1621523292
transform 1 0 36708 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1621523292
transform 1 0 37812 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_396
timestamp 1621523292
transform 1 0 37536 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_408
timestamp 1621523292
transform 1 0 38640 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_400
timestamp 1621523292
transform 1 0 37904 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_412
timestamp 1621523292
transform 1 0 39008 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1621523292
transform 1 0 40480 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_420
timestamp 1621523292
transform 1 0 39744 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_429
timestamp 1621523292
transform 1 0 40572 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_424
timestamp 1621523292
transform 1 0 40112 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_436
timestamp 1621523292
transform 1 0 41216 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1621523292
transform 1 0 43056 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_441
timestamp 1621523292
transform 1 0 41676 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_453
timestamp 1621523292
transform 1 0 42780 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_448
timestamp 1621523292
transform 1 0 42320 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_457
timestamp 1621523292
transform 1 0 43148 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_465
timestamp 1621523292
transform 1 0 43884 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_477
timestamp 1621523292
transform 1 0 44988 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_469
timestamp 1621523292
transform 1 0 44252 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1621523292
transform 1 0 45724 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_486
timestamp 1621523292
transform 1 0 45816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_498
timestamp 1621523292
transform 1 0 46920 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_481
timestamp 1621523292
transform 1 0 45356 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_493
timestamp 1621523292
transform 1 0 46460 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1621523292
transform 1 0 48300 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_510
timestamp 1621523292
transform 1 0 48024 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_522
timestamp 1621523292
transform 1 0 49128 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1621523292
transform 1 0 47564 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_514
timestamp 1621523292
transform 1 0 48392 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1621523292
transform 1 0 50968 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_534
timestamp 1621523292
transform 1 0 50232 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_543
timestamp 1621523292
transform 1 0 51060 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_526
timestamp 1621523292
transform 1 0 49496 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_538
timestamp 1621523292
transform 1 0 50600 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_555
timestamp 1621523292
transform 1 0 52164 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_567
timestamp 1621523292
transform 1 0 53268 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_550
timestamp 1621523292
transform 1 0 51704 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_562
timestamp 1621523292
transform 1 0 52808 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1621523292
transform 1 0 53544 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_579
timestamp 1621523292
transform 1 0 54372 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_571
timestamp 1621523292
transform 1 0 53636 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_583
timestamp 1621523292
transform 1 0 54740 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1556_
timestamp 1621523292
transform 1 0 56856 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2171_
timestamp 1621523292
transform 1 0 57224 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1621523292
transform 1 0 56212 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1621523292
transform 1 0 56580 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_591
timestamp 1621523292
transform 1 0 55476 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_72_600
timestamp 1621523292
transform 1 0 56304 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_609
timestamp 1621523292
transform 1 0 57132 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_595
timestamp 1621523292
transform 1 0 55844 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_606
timestamp 1621523292
transform 1 0 56856 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2320_
timestamp 1621523292
transform 1 0 57500 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1621523292
transform -1 0 58880 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1621523292
transform -1 0 58880 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output195
timestamp 1621523292
transform 1 0 57868 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1621523292
transform 1 0 58236 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_613
timestamp 1621523292
transform 1 0 57500 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_621
timestamp 1621523292
transform 1 0 58236 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1621523292
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1621523292
transform 1 0 1380 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_6
timestamp 1621523292
transform 1 0 1656 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_18
timestamp 1621523292
transform 1 0 2760 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1621523292
transform 1 0 3772 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_26
timestamp 1621523292
transform 1 0 3496 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_30
timestamp 1621523292
transform 1 0 3864 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_42
timestamp 1621523292
transform 1 0 4968 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_54
timestamp 1621523292
transform 1 0 6072 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1621523292
transform 1 0 9016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_66
timestamp 1621523292
transform 1 0 7176 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_78
timestamp 1621523292
transform 1 0 8280 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_87
timestamp 1621523292
transform 1 0 9108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_99
timestamp 1621523292
transform 1 0 10212 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_111
timestamp 1621523292
transform 1 0 11316 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_123
timestamp 1621523292
transform 1 0 12420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1621523292
transform 1 0 14260 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_135
timestamp 1621523292
transform 1 0 13524 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_144
timestamp 1621523292
transform 1 0 14352 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_156
timestamp 1621523292
transform 1 0 15456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_168
timestamp 1621523292
transform 1 0 16560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_180
timestamp 1621523292
transform 1 0 17664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_192
timestamp 1621523292
transform 1 0 18768 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _2017_
timestamp 1621523292
transform 1 0 20240 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1621523292
transform 1 0 19504 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_201
timestamp 1621523292
transform 1 0 19596 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_207
timestamp 1621523292
transform 1 0 20148 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_216
timestamp 1621523292
transform 1 0 20976 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2431_
timestamp 1621523292
transform 1 0 21896 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_74_224
timestamp 1621523292
transform 1 0 21712 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__and3_1  _2022_
timestamp 1621523292
transform 1 0 23736 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2441_
timestamp 1621523292
transform 1 0 25208 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1621523292
transform 1 0 24748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_242
timestamp 1621523292
transform 1 0 23368 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_251
timestamp 1621523292
transform 1 0 24196 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_258
timestamp 1621523292
transform 1 0 24840 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1621523292
transform 1 0 27048 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_278
timestamp 1621523292
transform 1 0 26680 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2041_
timestamp 1621523292
transform 1 0 29164 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2049_
timestamp 1621523292
transform 1 0 27968 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_285
timestamp 1621523292
transform 1 0 27324 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_291
timestamp 1621523292
transform 1 0 27876 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_298
timestamp 1621523292
transform 1 0 28520 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_304
timestamp 1621523292
transform 1 0 29072 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1621523292
transform 1 0 30452 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1621523292
transform 1 0 29992 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_wb_clk_i
timestamp 1621523292
transform 1 0 31096 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_310
timestamp 1621523292
transform 1 0 29624 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_315
timestamp 1621523292
transform 1 0 30084 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_322
timestamp 1621523292
transform 1 0 30728 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1957_
timestamp 1621523292
transform 1 0 32476 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_wb_clk_i
timestamp 1621523292
transform 1 0 31740 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_329
timestamp 1621523292
transform 1 0 31372 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_336
timestamp 1621523292
transform 1 0 32016 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_340
timestamp 1621523292
transform 1 0 32384 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_344
timestamp 1621523292
transform 1 0 32752 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1621523292
transform 1 0 35236 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_356
timestamp 1621523292
transform 1 0 33856 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_368
timestamp 1621523292
transform 1 0 34960 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_372
timestamp 1621523292
transform 1 0 35328 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_384
timestamp 1621523292
transform 1 0 36432 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_396
timestamp 1621523292
transform 1 0 37536 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_408
timestamp 1621523292
transform 1 0 38640 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1621523292
transform 1 0 40480 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_420
timestamp 1621523292
transform 1 0 39744 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_429
timestamp 1621523292
transform 1 0 40572 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_441
timestamp 1621523292
transform 1 0 41676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_453
timestamp 1621523292
transform 1 0 42780 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_465
timestamp 1621523292
transform 1 0 43884 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_477
timestamp 1621523292
transform 1 0 44988 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1621523292
transform 1 0 45724 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_486
timestamp 1621523292
transform 1 0 45816 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_498
timestamp 1621523292
transform 1 0 46920 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_510
timestamp 1621523292
transform 1 0 48024 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_522
timestamp 1621523292
transform 1 0 49128 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1621523292
transform 1 0 50968 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_534
timestamp 1621523292
transform 1 0 50232 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_543
timestamp 1621523292
transform 1 0 51060 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_555
timestamp 1621523292
transform 1 0 52164 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_567
timestamp 1621523292
transform 1 0 53268 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_579
timestamp 1621523292
transform 1 0 54372 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1621523292
transform 1 0 56212 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output234
timestamp 1621523292
transform 1 0 56764 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_591
timestamp 1621523292
transform 1 0 55476 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_600
timestamp 1621523292
transform 1 0 56304 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_604
timestamp 1621523292
transform 1 0 56672 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_609
timestamp 1621523292
transform 1 0 57132 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2321_
timestamp 1621523292
transform 1 0 57500 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1621523292
transform -1 0 58880 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_621
timestamp 1621523292
transform 1 0 58236 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1621523292
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1621523292
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1621523292
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1621523292
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1621523292
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1621523292
transform 1 0 6348 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_51
timestamp 1621523292
transform 1 0 5796 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_58
timestamp 1621523292
transform 1 0 6440 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_70
timestamp 1621523292
transform 1 0 7544 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_82
timestamp 1621523292
transform 1 0 8648 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_94
timestamp 1621523292
transform 1 0 9752 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_106
timestamp 1621523292
transform 1 0 10856 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1621523292
transform 1 0 11592 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_115
timestamp 1621523292
transform 1 0 11684 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_127
timestamp 1621523292
transform 1 0 12788 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_139
timestamp 1621523292
transform 1 0 13892 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_151
timestamp 1621523292
transform 1 0 14996 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1621523292
transform 1 0 16836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_163
timestamp 1621523292
transform 1 0 16100 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_172
timestamp 1621523292
transform 1 0 16928 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1621523292
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_196
timestamp 1621523292
transform 1 0 19136 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2430_
timestamp 1621523292
transform 1 0 20148 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_75_204
timestamp 1621523292
transform 1 0 19872 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _2021_
timestamp 1621523292
transform 1 0 22540 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1621523292
transform 1 0 22080 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_223
timestamp 1621523292
transform 1 0 21620 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_227
timestamp 1621523292
transform 1 0 21988 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_229
timestamp 1621523292
transform 1 0 22172 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2432_
timestamp 1621523292
transform 1 0 23736 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_241
timestamp 1621523292
transform 1 0 23276 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_245
timestamp 1621523292
transform 1 0 23644 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_262
timestamp 1621523292
transform 1 0 25208 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _2052_
timestamp 1621523292
transform 1 0 25852 0 1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_75_268
timestamp 1621523292
transform 1 0 25760 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_276
timestamp 1621523292
transform 1 0 26496 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2440_
timestamp 1621523292
transform 1 0 27784 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1621523292
transform 1 0 27324 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_284
timestamp 1621523292
transform 1 0 27232 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_286
timestamp 1621523292
transform 1 0 27416 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__nor2b_1  _2043_
timestamp 1621523292
transform 1 0 29624 0 1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2405_
timestamp 1621523292
transform 1 0 30636 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_306
timestamp 1621523292
transform 1 0 29256 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_315
timestamp 1621523292
transform 1 0 30084 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1621523292
transform 1 0 32568 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_337
timestamp 1621523292
transform 1 0 32108 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_341
timestamp 1621523292
transform 1 0 32476 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_343
timestamp 1621523292
transform 1 0 32660 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_355
timestamp 1621523292
transform 1 0 33764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1621523292
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1621523292
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_391
timestamp 1621523292
transform 1 0 37076 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1621523292
transform 1 0 37812 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_400
timestamp 1621523292
transform 1 0 37904 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_412
timestamp 1621523292
transform 1 0 39008 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_424
timestamp 1621523292
transform 1 0 40112 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_436
timestamp 1621523292
transform 1 0 41216 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1621523292
transform 1 0 43056 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_448
timestamp 1621523292
transform 1 0 42320 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_457
timestamp 1621523292
transform 1 0 43148 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_469
timestamp 1621523292
transform 1 0 44252 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_481
timestamp 1621523292
transform 1 0 45356 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_493
timestamp 1621523292
transform 1 0 46460 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1621523292
transform 1 0 48300 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1621523292
transform 1 0 47564 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_514
timestamp 1621523292
transform 1 0 48392 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_526
timestamp 1621523292
transform 1 0 49496 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_538
timestamp 1621523292
transform 1 0 50600 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_550
timestamp 1621523292
transform 1 0 51704 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_562
timestamp 1621523292
transform 1 0 52808 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1621523292
transform 1 0 53544 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_571
timestamp 1621523292
transform 1 0 53636 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_583
timestamp 1621523292
transform 1 0 54740 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1621523292
transform 1 0 57224 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1621523292
transform 1 0 56580 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_595
timestamp 1621523292
transform 1 0 55844 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_75_606
timestamp 1621523292
transform 1 0 56856 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1621523292
transform -1 0 58880 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output196
timestamp 1621523292
transform 1 0 57868 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_613
timestamp 1621523292
transform 1 0 57500 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1621523292
transform 1 0 58236 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1621523292
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1621523292
transform 1 0 1380 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_6
timestamp 1621523292
transform 1 0 1656 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_18
timestamp 1621523292
transform 1 0 2760 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1621523292
transform 1 0 3772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_26
timestamp 1621523292
transform 1 0 3496 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_30
timestamp 1621523292
transform 1 0 3864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_42
timestamp 1621523292
transform 1 0 4968 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_54
timestamp 1621523292
transform 1 0 6072 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1621523292
transform 1 0 9016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_66
timestamp 1621523292
transform 1 0 7176 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_78
timestamp 1621523292
transform 1 0 8280 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_87
timestamp 1621523292
transform 1 0 9108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_99
timestamp 1621523292
transform 1 0 10212 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_111
timestamp 1621523292
transform 1 0 11316 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_123
timestamp 1621523292
transform 1 0 12420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1621523292
transform 1 0 14260 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_135
timestamp 1621523292
transform 1 0 13524 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_144
timestamp 1621523292
transform 1 0 14352 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_156
timestamp 1621523292
transform 1 0 15456 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_168
timestamp 1621523292
transform 1 0 16560 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_180
timestamp 1621523292
transform 1 0 17664 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_192
timestamp 1621523292
transform 1 0 18768 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2018_
timestamp 1621523292
transform 1 0 21068 0 -1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2020_
timestamp 1621523292
transform 1 0 20424 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1621523292
transform 1 0 19504 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_201
timestamp 1621523292
transform 1 0 19596 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_209
timestamp 1621523292
transform 1 0 20332 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_213
timestamp 1621523292
transform 1 0 20700 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_222
timestamp 1621523292
transform 1 0 21528 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_234
timestamp 1621523292
transform 1 0 22632 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1860_
timestamp 1621523292
transform 1 0 23644 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1621523292
transform 1 0 24748 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_wb_clk_i
timestamp 1621523292
transform 1 0 25208 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_76_242
timestamp 1621523292
transform 1 0 23368 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_248
timestamp 1621523292
transform 1 0 23920 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_256
timestamp 1621523292
transform 1 0 24656 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_258
timestamp 1621523292
transform 1 0 24840 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2054_
timestamp 1621523292
transform 1 0 26128 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_76_265
timestamp 1621523292
transform 1 0 25484 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_271
timestamp 1621523292
transform 1 0 26036 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_278
timestamp 1621523292
transform 1 0 26680 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2047_
timestamp 1621523292
transform 1 0 27416 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _2048_
timestamp 1621523292
transform 1 0 28060 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_76_289
timestamp 1621523292
transform 1 0 27692 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_302
timestamp 1621523292
transform 1 0 28888 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2044_
timestamp 1621523292
transform 1 0 30452 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2046_
timestamp 1621523292
transform 1 0 29256 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1621523292
transform 1 0 29992 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_310
timestamp 1621523292
transform 1 0 29624 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_315
timestamp 1621523292
transform 1 0 30084 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_322
timestamp 1621523292
transform 1 0 30728 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1958_
timestamp 1621523292
transform 1 0 31372 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2406_
timestamp 1621523292
transform 1 0 32568 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_76_328
timestamp 1621523292
transform 1 0 31280 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_337
timestamp 1621523292
transform 1 0 32108 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_341
timestamp 1621523292
transform 1 0 32476 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1621523292
transform 1 0 35236 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_358
timestamp 1621523292
transform 1 0 34040 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_370
timestamp 1621523292
transform 1 0 35144 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_372
timestamp 1621523292
transform 1 0 35328 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_384
timestamp 1621523292
transform 1 0 36432 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_396
timestamp 1621523292
transform 1 0 37536 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_408
timestamp 1621523292
transform 1 0 38640 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1621523292
transform 1 0 40480 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_420
timestamp 1621523292
transform 1 0 39744 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_429
timestamp 1621523292
transform 1 0 40572 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_441
timestamp 1621523292
transform 1 0 41676 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_453
timestamp 1621523292
transform 1 0 42780 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_465
timestamp 1621523292
transform 1 0 43884 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_477
timestamp 1621523292
transform 1 0 44988 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1621523292
transform 1 0 45724 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_486
timestamp 1621523292
transform 1 0 45816 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_498
timestamp 1621523292
transform 1 0 46920 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_510
timestamp 1621523292
transform 1 0 48024 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_522
timestamp 1621523292
transform 1 0 49128 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1621523292
transform 1 0 50968 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_534
timestamp 1621523292
transform 1 0 50232 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_543
timestamp 1621523292
transform 1 0 51060 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_555
timestamp 1621523292
transform 1 0 52164 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_567
timestamp 1621523292
transform 1 0 53268 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_579
timestamp 1621523292
transform 1 0 54372 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2172_
timestamp 1621523292
transform 1 0 57224 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1621523292
transform 1 0 56212 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_591
timestamp 1621523292
transform 1 0 55476 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_76_600
timestamp 1621523292
transform 1 0 56304 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_608
timestamp 1621523292
transform 1 0 57040 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1621523292
transform -1 0 58880 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output235
timestamp 1621523292
transform 1 0 57868 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_613
timestamp 1621523292
transform 1 0 57500 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_621
timestamp 1621523292
transform 1 0 58236 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1621523292
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1621523292
transform 1 0 1380 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1621523292
transform 1 0 2484 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1621523292
transform 1 0 3588 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1621523292
transform 1 0 4692 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1621523292
transform 1 0 6348 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_51
timestamp 1621523292
transform 1 0 5796 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_58
timestamp 1621523292
transform 1 0 6440 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_70
timestamp 1621523292
transform 1 0 7544 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_82
timestamp 1621523292
transform 1 0 8648 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_94
timestamp 1621523292
transform 1 0 9752 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_106
timestamp 1621523292
transform 1 0 10856 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1621523292
transform 1 0 11592 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_115
timestamp 1621523292
transform 1 0 11684 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_127
timestamp 1621523292
transform 1 0 12788 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_139
timestamp 1621523292
transform 1 0 13892 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_151
timestamp 1621523292
transform 1 0 14996 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1621523292
transform 1 0 16836 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_163
timestamp 1621523292
transform 1 0 16100 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_77_172
timestamp 1621523292
transform 1 0 16928 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1845_
timestamp 1621523292
transform 1 0 17664 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1847_
timestamp 1621523292
transform 1 0 18492 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_183
timestamp 1621523292
transform 1 0 17940 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_192
timestamp 1621523292
transform 1 0 18768 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1850_
timestamp 1621523292
transform 1 0 20332 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1851_
timestamp 1621523292
transform 1 0 20976 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_204
timestamp 1621523292
transform 1 0 19872 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_208
timestamp 1621523292
transform 1 0 20240 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_212
timestamp 1621523292
transform 1 0 20608 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2369_
timestamp 1621523292
transform 1 0 22540 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1621523292
transform 1 0 22080 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_219
timestamp 1621523292
transform 1 0 21252 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_227
timestamp 1621523292
transform 1 0 21988 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_229
timestamp 1621523292
transform 1 0 22172 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2370_
timestamp 1621523292
transform 1 0 24380 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_77_249
timestamp 1621523292
transform 1 0 24012 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2055_
timestamp 1621523292
transform 1 0 26496 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_77_269
timestamp 1621523292
transform 1 0 25852 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_275
timestamp 1621523292
transform 1 0 26404 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_281
timestamp 1621523292
transform 1 0 26956 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _2056_
timestamp 1621523292
transform 1 0 27968 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1621523292
transform 1 0 27324 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_286
timestamp 1621523292
transform 1 0 27416 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_301
timestamp 1621523292
transform 1 0 28796 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_305
timestamp 1621523292
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2439_
timestamp 1621523292
transform 1 0 29256 0 1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_77_322
timestamp 1621523292
transform 1 0 30728 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1959_
timestamp 1621523292
transform 1 0 31740 0 1 44064
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1961_
timestamp 1621523292
transform 1 0 33028 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1621523292
transform 1 0 32568 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_330
timestamp 1621523292
transform 1 0 31464 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_338
timestamp 1621523292
transform 1 0 32200 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_343
timestamp 1621523292
transform 1 0 32660 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_350
timestamp 1621523292
transform 1 0 33304 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_362
timestamp 1621523292
transform 1 0 34408 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_374
timestamp 1621523292
transform 1 0 35512 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_386
timestamp 1621523292
transform 1 0 36616 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1621523292
transform 1 0 37812 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_398
timestamp 1621523292
transform 1 0 37720 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_400
timestamp 1621523292
transform 1 0 37904 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_412
timestamp 1621523292
transform 1 0 39008 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_424
timestamp 1621523292
transform 1 0 40112 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_436
timestamp 1621523292
transform 1 0 41216 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1621523292
transform 1 0 43056 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_448
timestamp 1621523292
transform 1 0 42320 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_457
timestamp 1621523292
transform 1 0 43148 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_469
timestamp 1621523292
transform 1 0 44252 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_481
timestamp 1621523292
transform 1 0 45356 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_493
timestamp 1621523292
transform 1 0 46460 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1621523292
transform 1 0 48300 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_505
timestamp 1621523292
transform 1 0 47564 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_77_514
timestamp 1621523292
transform 1 0 48392 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_526
timestamp 1621523292
transform 1 0 49496 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_538
timestamp 1621523292
transform 1 0 50600 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_550
timestamp 1621523292
transform 1 0 51704 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_562
timestamp 1621523292
transform 1 0 52808 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1621523292
transform 1 0 53544 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_571
timestamp 1621523292
transform 1 0 53636 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_583
timestamp 1621523292
transform 1 0 54740 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1554_
timestamp 1621523292
transform 1 0 56856 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2173_
timestamp 1621523292
transform 1 0 56212 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_595
timestamp 1621523292
transform 1 0 55844 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_602
timestamp 1621523292
transform 1 0 56488 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_609
timestamp 1621523292
transform 1 0 57132 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2322_
timestamp 1621523292
transform 1 0 57500 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1621523292
transform -1 0 58880 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1621523292
transform 1 0 58236 0 1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1621523292
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1621523292
transform 1 0 1380 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_6
timestamp 1621523292
transform 1 0 1656 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_18
timestamp 1621523292
transform 1 0 2760 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1621523292
transform 1 0 3772 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_26
timestamp 1621523292
transform 1 0 3496 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_30
timestamp 1621523292
transform 1 0 3864 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_42
timestamp 1621523292
transform 1 0 4968 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_54
timestamp 1621523292
transform 1 0 6072 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1621523292
transform 1 0 9016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_66
timestamp 1621523292
transform 1 0 7176 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_78
timestamp 1621523292
transform 1 0 8280 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_87
timestamp 1621523292
transform 1 0 9108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_99
timestamp 1621523292
transform 1 0 10212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_111
timestamp 1621523292
transform 1 0 11316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_123
timestamp 1621523292
transform 1 0 12420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1621523292
transform 1 0 14260 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_135
timestamp 1621523292
transform 1 0 13524 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_144
timestamp 1621523292
transform 1 0 14352 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2364_
timestamp 1621523292
transform 1 0 16744 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_78_156
timestamp 1621523292
transform 1 0 15456 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_168
timestamp 1621523292
transform 1 0 16560 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _1849_
timestamp 1621523292
transform 1 0 18584 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_186
timestamp 1621523292
transform 1 0 18216 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_196
timestamp 1621523292
transform 1 0 19136 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2366_
timestamp 1621523292
transform 1 0 20240 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1621523292
transform 1 0 19504 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_201
timestamp 1621523292
transform 1 0 19596 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_207
timestamp 1621523292
transform 1 0 20148 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1859_
timestamp 1621523292
transform 1 0 22540 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_78_224
timestamp 1621523292
transform 1 0 21712 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_232
timestamp 1621523292
transform 1 0 22448 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_239
timestamp 1621523292
transform 1 0 23092 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1862_
timestamp 1621523292
transform 1 0 23828 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1621523292
transform 1 0 24748 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_253
timestamp 1621523292
transform 1 0 24380 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_258
timestamp 1621523292
transform 1 0 24840 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_262
timestamp 1621523292
transform 1 0 25208 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2053_
timestamp 1621523292
transform 1 0 27140 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2442_
timestamp 1621523292
transform 1 0 25300 0 -1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_78_279
timestamp 1621523292
transform 1 0 26772 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2045_
timestamp 1621523292
transform 1 0 29072 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2061_
timestamp 1621523292
transform 1 0 27784 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_wb_clk_i
timestamp 1621523292
transform 1 0 28428 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_286
timestamp 1621523292
transform 1 0 27416 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_293
timestamp 1621523292
transform 1 0 28060 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_300
timestamp 1621523292
transform 1 0 28704 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1962_
timestamp 1621523292
transform 1 0 30452 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1621523292
transform 1 0 29992 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_307
timestamp 1621523292
transform 1 0 29348 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_313
timestamp 1621523292
transform 1 0 29900 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_315
timestamp 1621523292
transform 1 0 30084 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_327
timestamp 1621523292
transform 1 0 31188 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1960_
timestamp 1621523292
transform 1 0 32016 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_335
timestamp 1621523292
transform 1 0 31924 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_340
timestamp 1621523292
transform 1 0 32384 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1621523292
transform 1 0 35236 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_352
timestamp 1621523292
transform 1 0 33488 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_364
timestamp 1621523292
transform 1 0 34592 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_370
timestamp 1621523292
transform 1 0 35144 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_372
timestamp 1621523292
transform 1 0 35328 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_384
timestamp 1621523292
transform 1 0 36432 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_396
timestamp 1621523292
transform 1 0 37536 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_408
timestamp 1621523292
transform 1 0 38640 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1621523292
transform 1 0 40480 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_420
timestamp 1621523292
transform 1 0 39744 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_429
timestamp 1621523292
transform 1 0 40572 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_441
timestamp 1621523292
transform 1 0 41676 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_453
timestamp 1621523292
transform 1 0 42780 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_465
timestamp 1621523292
transform 1 0 43884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_477
timestamp 1621523292
transform 1 0 44988 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1621523292
transform 1 0 45724 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_486
timestamp 1621523292
transform 1 0 45816 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_498
timestamp 1621523292
transform 1 0 46920 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_510
timestamp 1621523292
transform 1 0 48024 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_522
timestamp 1621523292
transform 1 0 49128 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1621523292
transform 1 0 50968 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_534
timestamp 1621523292
transform 1 0 50232 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_543
timestamp 1621523292
transform 1 0 51060 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_555
timestamp 1621523292
transform 1 0 52164 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_567
timestamp 1621523292
transform 1 0 53268 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_579
timestamp 1621523292
transform 1 0 54372 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1552_
timestamp 1621523292
transform 1 0 57224 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1621523292
transform 1 0 56212 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_591
timestamp 1621523292
transform 1 0 55476 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_78_600
timestamp 1621523292
transform 1 0 56304 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_608
timestamp 1621523292
transform 1 0 57040 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1621523292
transform -1 0 58880 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output197
timestamp 1621523292
transform 1 0 57868 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_613
timestamp 1621523292
transform 1 0 57500 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_621
timestamp 1621523292
transform 1 0 58236 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1621523292
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1621523292
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 1621523292
transform 1 0 1380 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_6
timestamp 1621523292
transform 1 0 1656 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_18
timestamp 1621523292
transform 1 0 2760 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1621523292
transform 1 0 1380 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1621523292
transform 1 0 2484 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1621523292
transform 1 0 3772 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_30
timestamp 1621523292
transform 1 0 3864 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_42
timestamp 1621523292
transform 1 0 4968 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_27
timestamp 1621523292
transform 1 0 3588 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_30
timestamp 1621523292
transform 1 0 3864 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_42
timestamp 1621523292
transform 1 0 4968 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1621523292
transform 1 0 6348 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_54
timestamp 1621523292
transform 1 0 6072 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_58
timestamp 1621523292
transform 1 0 6440 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_54
timestamp 1621523292
transform 1 0 6072 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1621523292
transform 1 0 9016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_70
timestamp 1621523292
transform 1 0 7544 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_82
timestamp 1621523292
transform 1 0 8648 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_66
timestamp 1621523292
transform 1 0 7176 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_78
timestamp 1621523292
transform 1 0 8280 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_87
timestamp 1621523292
transform 1 0 9108 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_94
timestamp 1621523292
transform 1 0 9752 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_106
timestamp 1621523292
transform 1 0 10856 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_99
timestamp 1621523292
transform 1 0 10212 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1621523292
transform 1 0 11592 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_115
timestamp 1621523292
transform 1 0 11684 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_127
timestamp 1621523292
transform 1 0 12788 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_111
timestamp 1621523292
transform 1 0 11316 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_123
timestamp 1621523292
transform 1 0 12420 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1716_
timestamp 1621523292
transform 1 0 14720 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2359_
timestamp 1621523292
transform 1 0 13984 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1621523292
transform 1 0 14260 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_139
timestamp 1621523292
transform 1 0 13892 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_135
timestamp 1621523292
transform 1 0 13524 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_144
timestamp 1621523292
transform 1 0 14352 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_151
timestamp 1621523292
transform 1 0 14996 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2363_
timestamp 1621523292
transform 1 0 15732 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1621523292
transform 1 0 16836 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_156
timestamp 1621523292
transform 1 0 15456 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_168
timestamp 1621523292
transform 1 0 16560 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_172
timestamp 1621523292
transform 1 0 16928 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_185
timestamp 1621523292
transform 1 0 18124 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_175
timestamp 1621523292
transform 1 0 17204 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_183
timestamp 1621523292
transform 1 0 17940 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_176
timestamp 1621523292
transform 1 0 17296 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1846_
timestamp 1621523292
transform 1 0 17388 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1843_
timestamp 1621523292
transform 1 0 17572 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_192
timestamp 1621523292
transform 1 0 18768 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_189
timestamp 1621523292
transform 1 0 18492 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1844_
timestamp 1621523292
transform 1 0 18492 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2365_
timestamp 1621523292
transform 1 0 18584 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1848_
timestamp 1621523292
transform 1 0 19964 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1852_
timestamp 1621523292
transform 1 0 20700 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1621523292
transform 1 0 19504 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_wb_clk_i
timestamp 1621523292
transform 1 0 20608 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_206
timestamp 1621523292
transform 1 0 20056 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_212
timestamp 1621523292
transform 1 0 20608 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_201
timestamp 1621523292
transform 1 0 19596 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_208
timestamp 1621523292
transform 1 0 20240 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_215
timestamp 1621523292
transform 1 0 20884 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1854_
timestamp 1621523292
transform 1 0 21436 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1856_
timestamp 1621523292
transform 1 0 22540 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2368_
timestamp 1621523292
transform 1 0 22724 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1621523292
transform 1 0 22080 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_219
timestamp 1621523292
transform 1 0 21252 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_227
timestamp 1621523292
transform 1 0 21988 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_229
timestamp 1621523292
transform 1 0 22172 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_237
timestamp 1621523292
transform 1 0 22908 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_229
timestamp 1621523292
transform 1 0 22172 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_80_251
timestamp 1621523292
transform 1 0 24196 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_79_244
timestamp 1621523292
transform 1 0 23552 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1858_
timestamp 1621523292
transform 1 0 23276 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_258
timestamp 1621523292
transform 1 0 24840 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_256
timestamp 1621523292
transform 1 0 24656 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_252
timestamp 1621523292
transform 1 0 24288 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1621523292
transform 1 0 24748 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1863_
timestamp 1621523292
transform 1 0 25024 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1861_
timestamp 1621523292
transform 1 0 24380 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2371_
timestamp 1621523292
transform 1 0 25208 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1864_
timestamp 1621523292
transform 1 0 27048 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__nor2b_1  _2057_
timestamp 1621523292
transform 1 0 26036 0 1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_79_263
timestamp 1621523292
transform 1 0 25300 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_79_276
timestamp 1621523292
transform 1 0 26496 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_278
timestamp 1621523292
transform 1 0 26680 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_285
timestamp 1621523292
transform 1 0 27324 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_294
timestamp 1621523292
transform 1 0 28152 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_286
timestamp 1621523292
transform 1 0 27416 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_284
timestamp 1621523292
transform 1 0 27232 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1621523292
transform 1 0 27324 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _2060_
timestamp 1621523292
transform 1 0 27784 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_305
timestamp 1621523292
transform 1 0 29164 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_302
timestamp 1621523292
transform 1 0 28888 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_298
timestamp 1621523292
transform 1 0 28520 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2058_
timestamp 1621523292
transform 1 0 28612 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2443_
timestamp 1621523292
transform 1 0 27692 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2407_
timestamp 1621523292
transform 1 0 29256 0 1 45152
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2408_
timestamp 1621523292
transform 1 0 31096 0 -1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1621523292
transform 1 0 29992 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_wb_clk_i
timestamp 1621523292
transform 1 0 30452 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_79_322
timestamp 1621523292
transform 1 0 30728 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_313
timestamp 1621523292
transform 1 0 29900 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_315
timestamp 1621523292
transform 1 0 30084 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_322
timestamp 1621523292
transform 1 0 30728 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1963_
timestamp 1621523292
transform 1 0 31280 0 1 45152
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1965_
timestamp 1621523292
transform 1 0 33028 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1621523292
transform 1 0 32568 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_333
timestamp 1621523292
transform 1 0 31740 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_341
timestamp 1621523292
transform 1 0 32476 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_343
timestamp 1621523292
transform 1 0 32660 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_342
timestamp 1621523292
transform 1 0 32568 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1792_
timestamp 1621523292
transform 1 0 33396 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1621523292
transform 1 0 35236 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_350
timestamp 1621523292
transform 1 0 33304 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_362
timestamp 1621523292
transform 1 0 34408 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_350
timestamp 1621523292
transform 1 0 33304 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_354
timestamp 1621523292
transform 1 0 33672 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_366
timestamp 1621523292
transform 1 0 34776 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_370
timestamp 1621523292
transform 1 0 35144 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_374
timestamp 1621523292
transform 1 0 35512 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_386
timestamp 1621523292
transform 1 0 36616 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_372
timestamp 1621523292
transform 1 0 35328 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_384
timestamp 1621523292
transform 1 0 36432 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1621523292
transform 1 0 37812 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_79_398
timestamp 1621523292
transform 1 0 37720 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_400
timestamp 1621523292
transform 1 0 37904 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_412
timestamp 1621523292
transform 1 0 39008 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_396
timestamp 1621523292
transform 1 0 37536 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_408
timestamp 1621523292
transform 1 0 38640 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1621523292
transform 1 0 40480 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_424
timestamp 1621523292
transform 1 0 40112 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_436
timestamp 1621523292
transform 1 0 41216 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_420
timestamp 1621523292
transform 1 0 39744 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_429
timestamp 1621523292
transform 1 0 40572 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1621523292
transform 1 0 43056 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_448
timestamp 1621523292
transform 1 0 42320 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_457
timestamp 1621523292
transform 1 0 43148 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_441
timestamp 1621523292
transform 1 0 41676 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_453
timestamp 1621523292
transform 1 0 42780 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_469
timestamp 1621523292
transform 1 0 44252 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_465
timestamp 1621523292
transform 1 0 43884 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_477
timestamp 1621523292
transform 1 0 44988 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1621523292
transform 1 0 45724 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_481
timestamp 1621523292
transform 1 0 45356 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_493
timestamp 1621523292
transform 1 0 46460 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_486
timestamp 1621523292
transform 1 0 45816 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_498
timestamp 1621523292
transform 1 0 46920 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1621523292
transform 1 0 48300 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_505
timestamp 1621523292
transform 1 0 47564 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_514
timestamp 1621523292
transform 1 0 48392 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_510
timestamp 1621523292
transform 1 0 48024 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_522
timestamp 1621523292
transform 1 0 49128 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1621523292
transform 1 0 50968 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_526
timestamp 1621523292
transform 1 0 49496 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_538
timestamp 1621523292
transform 1 0 50600 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_534
timestamp 1621523292
transform 1 0 50232 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_543
timestamp 1621523292
transform 1 0 51060 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_550
timestamp 1621523292
transform 1 0 51704 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_562
timestamp 1621523292
transform 1 0 52808 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_555
timestamp 1621523292
transform 1 0 52164 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_567
timestamp 1621523292
transform 1 0 53268 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1621523292
transform 1 0 53544 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_571
timestamp 1621523292
transform 1 0 53636 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_583
timestamp 1621523292
transform 1 0 54740 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_579
timestamp 1621523292
transform 1 0 54372 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1621523292
transform 1 0 57224 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2174_
timestamp 1621523292
transform 1 0 56856 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1621523292
transform 1 0 56212 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1621523292
transform 1 0 56580 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_595
timestamp 1621523292
transform 1 0 55844 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_606
timestamp 1621523292
transform 1 0 56856 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_591
timestamp 1621523292
transform 1 0 55476 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_600
timestamp 1621523292
transform 1 0 56304 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_609
timestamp 1621523292
transform 1 0 57132 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2323_
timestamp 1621523292
transform 1 0 57500 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1621523292
transform -1 0 58880 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1621523292
transform -1 0 58880 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output236
timestamp 1621523292
transform 1 0 57868 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_613
timestamp 1621523292
transform 1 0 57500 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_621
timestamp 1621523292
transform 1 0 58236 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1621523292
transform 1 0 58236 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1621523292
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1621523292
transform 1 0 1380 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_6
timestamp 1621523292
transform 1 0 1656 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_18
timestamp 1621523292
transform 1 0 2760 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1621523292
transform 1 0 3864 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1621523292
transform 1 0 4968 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1621523292
transform 1 0 6348 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_54
timestamp 1621523292
transform 1 0 6072 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_58
timestamp 1621523292
transform 1 0 6440 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_70
timestamp 1621523292
transform 1 0 7544 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_82
timestamp 1621523292
transform 1 0 8648 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_94
timestamp 1621523292
transform 1 0 9752 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_106
timestamp 1621523292
transform 1 0 10856 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1621523292
transform 1 0 11592 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_115
timestamp 1621523292
transform 1 0 11684 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_127
timestamp 1621523292
transform 1 0 12788 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2360_
timestamp 1621523292
transform 1 0 13432 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_133
timestamp 1621523292
transform 1 0 13340 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_150
timestamp 1621523292
transform 1 0 14904 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1835_
timestamp 1621523292
transform 1 0 15272 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1837_
timestamp 1621523292
transform 1 0 15916 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1621523292
transform 1 0 16836 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_157
timestamp 1621523292
transform 1 0 15548 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_164
timestamp 1621523292
transform 1 0 16192 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_170
timestamp 1621523292
transform 1 0 16744 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_172
timestamp 1621523292
transform 1 0 16928 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2344_
timestamp 1621523292
transform 1 0 17572 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_81_178
timestamp 1621523292
transform 1 0 17480 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_195
timestamp 1621523292
transform 1 0 19044 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2343_
timestamp 1621523292
transform 1 0 19412 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_81_215
timestamp 1621523292
transform 1 0 20884 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1853_
timestamp 1621523292
transform 1 0 21436 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1855_
timestamp 1621523292
transform 1 0 22540 0 1 46240
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1621523292
transform 1 0 22080 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_224
timestamp 1621523292
transform 1 0 21712 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_229
timestamp 1621523292
transform 1 0 22172 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_238
timestamp 1621523292
transform 1 0 23000 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1857_
timestamp 1621523292
transform 1 0 23368 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1865_
timestamp 1621523292
transform 1 0 24564 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_245
timestamp 1621523292
transform 1 0 23644 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_253
timestamp 1621523292
transform 1 0 24380 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_261
timestamp 1621523292
transform 1 0 25116 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2444_
timestamp 1621523292
transform 1 0 25484 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_81_281
timestamp 1621523292
transform 1 0 26956 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2059_
timestamp 1621523292
transform 1 0 27784 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2410_
timestamp 1621523292
transform 1 0 28888 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1621523292
transform 1 0 27324 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_286
timestamp 1621523292
transform 1 0 27416 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_293
timestamp 1621523292
transform 1 0 28060 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_301
timestamp 1621523292
transform 1 0 28796 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_1  _1964_
timestamp 1621523292
transform 1 0 31188 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_318
timestamp 1621523292
transform 1 0 30360 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_326
timestamp 1621523292
transform 1 0 31096 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1966_
timestamp 1621523292
transform 1 0 31924 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2335_
timestamp 1621523292
transform 1 0 33028 0 1 46240
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1621523292
transform 1 0 32568 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_331
timestamp 1621523292
transform 1 0 31556 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_338
timestamp 1621523292
transform 1 0 32200 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_343
timestamp 1621523292
transform 1 0 32660 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_363
timestamp 1621523292
transform 1 0 34500 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_375
timestamp 1621523292
transform 1 0 35604 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_387
timestamp 1621523292
transform 1 0 36708 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1621523292
transform 1 0 37812 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_400
timestamp 1621523292
transform 1 0 37904 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_412
timestamp 1621523292
transform 1 0 39008 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_424
timestamp 1621523292
transform 1 0 40112 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_436
timestamp 1621523292
transform 1 0 41216 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1621523292
transform 1 0 43056 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_448
timestamp 1621523292
transform 1 0 42320 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_457
timestamp 1621523292
transform 1 0 43148 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_469
timestamp 1621523292
transform 1 0 44252 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_481
timestamp 1621523292
transform 1 0 45356 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_493
timestamp 1621523292
transform 1 0 46460 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1621523292
transform 1 0 48300 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_505
timestamp 1621523292
transform 1 0 47564 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_81_514
timestamp 1621523292
transform 1 0 48392 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_526
timestamp 1621523292
transform 1 0 49496 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_538
timestamp 1621523292
transform 1 0 50600 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_550
timestamp 1621523292
transform 1 0 51704 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_562
timestamp 1621523292
transform 1 0 52808 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1621523292
transform 1 0 53544 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_571
timestamp 1621523292
transform 1 0 53636 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_583
timestamp 1621523292
transform 1 0 54740 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_595
timestamp 1621523292
transform 1 0 55844 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_607
timestamp 1621523292
transform 1 0 56948 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1621523292
transform -1 0 58880 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output198
timestamp 1621523292
transform 1 0 57868 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_615
timestamp 1621523292
transform 1 0 57684 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_621
timestamp 1621523292
transform 1 0 58236 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1621523292
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1621523292
transform 1 0 1380 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1621523292
transform 1 0 2484 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1621523292
transform 1 0 3772 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_27
timestamp 1621523292
transform 1 0 3588 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_30
timestamp 1621523292
transform 1 0 3864 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_42
timestamp 1621523292
transform 1 0 4968 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_54
timestamp 1621523292
transform 1 0 6072 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1621523292
transform 1 0 9016 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_66
timestamp 1621523292
transform 1 0 7176 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_78
timestamp 1621523292
transform 1 0 8280 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_87
timestamp 1621523292
transform 1 0 9108 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_99
timestamp 1621523292
transform 1 0 10212 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_111
timestamp 1621523292
transform 1 0 11316 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_123
timestamp 1621523292
transform 1 0 12420 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1836_
timestamp 1621523292
transform 1 0 14720 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1621523292
transform 1 0 14260 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_135
timestamp 1621523292
transform 1 0 13524 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_82_144
timestamp 1621523292
transform 1 0 14352 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1840_
timestamp 1621523292
transform 1 0 16100 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1842_
timestamp 1621523292
transform 1 0 16836 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_154
timestamp 1621523292
transform 1 0 15272 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_162
timestamp 1621523292
transform 1 0 16008 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_167
timestamp 1621523292
transform 1 0 16468 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_174
timestamp 1621523292
transform 1 0 17112 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1795_
timestamp 1621523292
transform 1 0 18584 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_186
timestamp 1621523292
transform 1 0 18216 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_196
timestamp 1621523292
transform 1 0 19136 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1793_
timestamp 1621523292
transform 1 0 19964 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2367_
timestamp 1621523292
transform 1 0 20884 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1621523292
transform 1 0 19504 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_201
timestamp 1621523292
transform 1 0 19596 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_208
timestamp 1621523292
transform 1 0 20240 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_214
timestamp 1621523292
transform 1 0 20792 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_wb_clk_i
timestamp 1621523292
transform 1 0 22724 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_231
timestamp 1621523292
transform 1 0 22356 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_238
timestamp 1621523292
transform 1 0 23000 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1866_
timestamp 1621523292
transform 1 0 24104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1868_
timestamp 1621523292
transform 1 0 25208 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1621523292
transform 1 0 24748 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_wb_clk_i
timestamp 1621523292
transform 1 0 23460 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_242
timestamp 1621523292
transform 1 0 23368 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_246
timestamp 1621523292
transform 1 0 23736 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_253
timestamp 1621523292
transform 1 0 24380 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_258
timestamp 1621523292
transform 1 0 24840 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2063_
timestamp 1621523292
transform 1 0 26588 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_82_268
timestamp 1621523292
transform 1 0 25760 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_276
timestamp 1621523292
transform 1 0 26496 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_283
timestamp 1621523292
transform 1 0 27140 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_2  _2069_
timestamp 1621523292
transform 1 0 27692 0 -1 47328
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_82_299
timestamp 1621523292
transform 1 0 28612 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1967_
timestamp 1621523292
transform 1 0 31004 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1969_
timestamp 1621523292
transform 1 0 29348 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1621523292
transform 1 0 29992 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_310
timestamp 1621523292
transform 1 0 29624 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_315
timestamp 1621523292
transform 1 0 30084 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_323
timestamp 1621523292
transform 1 0 30820 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  _2336_
timestamp 1621523292
transform 1 0 32292 0 -1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_82_331
timestamp 1621523292
transform 1 0 31556 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2082_
timestamp 1621523292
transform 1 0 34132 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1621523292
transform 1 0 35236 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_355
timestamp 1621523292
transform 1 0 33764 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_362
timestamp 1621523292
transform 1 0 34408 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_370
timestamp 1621523292
transform 1 0 35144 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_372
timestamp 1621523292
transform 1 0 35328 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_384
timestamp 1621523292
transform 1 0 36432 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_396
timestamp 1621523292
transform 1 0 37536 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_408
timestamp 1621523292
transform 1 0 38640 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1621523292
transform 1 0 40480 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_420
timestamp 1621523292
transform 1 0 39744 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_429
timestamp 1621523292
transform 1 0 40572 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_441
timestamp 1621523292
transform 1 0 41676 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_453
timestamp 1621523292
transform 1 0 42780 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_465
timestamp 1621523292
transform 1 0 43884 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_477
timestamp 1621523292
transform 1 0 44988 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1621523292
transform 1 0 45724 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_486
timestamp 1621523292
transform 1 0 45816 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_498
timestamp 1621523292
transform 1 0 46920 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_510
timestamp 1621523292
transform 1 0 48024 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_522
timestamp 1621523292
transform 1 0 49128 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1621523292
transform 1 0 50968 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_534
timestamp 1621523292
transform 1 0 50232 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_543
timestamp 1621523292
transform 1 0 51060 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_555
timestamp 1621523292
transform 1 0 52164 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_567
timestamp 1621523292
transform 1 0 53268 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_579
timestamp 1621523292
transform 1 0 54372 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1621523292
transform 1 0 56212 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1621523292
transform 1 0 56856 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_591
timestamp 1621523292
transform 1 0 55476 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_82_600
timestamp 1621523292
transform 1 0 56304 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_609
timestamp 1621523292
transform 1 0 57132 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1546_
timestamp 1621523292
transform 1 0 57500 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1621523292
transform -1 0 58880 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_616
timestamp 1621523292
transform 1 0 57776 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_624
timestamp 1621523292
transform 1 0 58512 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1621523292
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1621523292
transform 1 0 1380 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_6
timestamp 1621523292
transform 1 0 1656 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_18
timestamp 1621523292
transform 1 0 2760 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_30
timestamp 1621523292
transform 1 0 3864 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_42
timestamp 1621523292
transform 1 0 4968 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1621523292
transform 1 0 6348 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_54
timestamp 1621523292
transform 1 0 6072 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_58
timestamp 1621523292
transform 1 0 6440 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_70
timestamp 1621523292
transform 1 0 7544 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_82
timestamp 1621523292
transform 1 0 8648 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_94
timestamp 1621523292
transform 1 0 9752 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_106
timestamp 1621523292
transform 1 0 10856 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1621523292
transform 1 0 11592 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_115
timestamp 1621523292
transform 1 0 11684 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_127
timestamp 1621523292
transform 1 0 12788 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2361_
timestamp 1621523292
transform 1 0 14352 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_139
timestamp 1621523292
transform 1 0 13892 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_143
timestamp 1621523292
transform 1 0 14260 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1621523292
transform 1 0 16836 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_160
timestamp 1621523292
transform 1 0 15824 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_168
timestamp 1621523292
transform 1 0 16560 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_172
timestamp 1621523292
transform 1 0 16928 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1794_
timestamp 1621523292
transform 1 0 19136 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2362_
timestamp 1621523292
transform 1 0 17296 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_83_192
timestamp 1621523292
transform 1 0 18768 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1796_
timestamp 1621523292
transform 1 0 20884 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1799_
timestamp 1621523292
transform 1 0 20148 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_199
timestamp 1621523292
transform 1 0 19412 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_211
timestamp 1621523292
transform 1 0 20516 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_218
timestamp 1621523292
transform 1 0 21160 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1621523292
transform 1 0 22080 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_226
timestamp 1621523292
transform 1 0 21896 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_229
timestamp 1621523292
transform 1 0 22172 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2372_
timestamp 1621523292
transform 1 0 23920 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_83_241
timestamp 1621523292
transform 1 0 23276 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_247
timestamp 1621523292
transform 1 0 23828 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _2066_
timestamp 1621523292
transform 1 0 26312 0 1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_83_264
timestamp 1621523292
transform 1 0 25392 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_272
timestamp 1621523292
transform 1 0 26128 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_281
timestamp 1621523292
transform 1 0 26956 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _2062_
timestamp 1621523292
transform 1 0 27784 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1621523292
transform 1 0 27324 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_286
timestamp 1621523292
transform 1 0 27416 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_299
timestamp 1621523292
transform 1 0 28612 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1970_
timestamp 1621523292
transform 1 0 29532 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2409_
timestamp 1621523292
transform 1 0 30636 0 1 47328
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_83_307
timestamp 1621523292
transform 1 0 29348 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_83_315
timestamp 1621523292
transform 1 0 30084 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2083_
timestamp 1621523292
transform 1 0 33120 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1621523292
transform 1 0 32568 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_337
timestamp 1621523292
transform 1 0 32108 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_341
timestamp 1621523292
transform 1 0 32476 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_343
timestamp 1621523292
transform 1 0 32660 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_347
timestamp 1621523292
transform 1 0 33028 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_354
timestamp 1621523292
transform 1 0 33672 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_366
timestamp 1621523292
transform 1 0 34776 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_378
timestamp 1621523292
transform 1 0 35880 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_390
timestamp 1621523292
transform 1 0 36984 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1621523292
transform 1 0 37812 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_398
timestamp 1621523292
transform 1 0 37720 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_400
timestamp 1621523292
transform 1 0 37904 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_412
timestamp 1621523292
transform 1 0 39008 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_424
timestamp 1621523292
transform 1 0 40112 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_436
timestamp 1621523292
transform 1 0 41216 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1621523292
transform 1 0 43056 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_448
timestamp 1621523292
transform 1 0 42320 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_457
timestamp 1621523292
transform 1 0 43148 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_469
timestamp 1621523292
transform 1 0 44252 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_481
timestamp 1621523292
transform 1 0 45356 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_493
timestamp 1621523292
transform 1 0 46460 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1621523292
transform 1 0 48300 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_505
timestamp 1621523292
transform 1 0 47564 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_514
timestamp 1621523292
transform 1 0 48392 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_526
timestamp 1621523292
transform 1 0 49496 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_538
timestamp 1621523292
transform 1 0 50600 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_550
timestamp 1621523292
transform 1 0 51704 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_562
timestamp 1621523292
transform 1 0 52808 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1621523292
transform 1 0 53544 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_571
timestamp 1621523292
transform 1 0 53636 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_583
timestamp 1621523292
transform 1 0 54740 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1551_
timestamp 1621523292
transform 1 0 57224 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_595
timestamp 1621523292
transform 1 0 55844 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_607
timestamp 1621523292
transform 1 0 56948 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1621523292
transform -1 0 58880 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output238
timestamp 1621523292
transform 1 0 57868 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_613
timestamp 1621523292
transform 1 0 57500 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_621
timestamp 1621523292
transform 1 0 58236 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1621523292
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1621523292
transform 1 0 1380 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_6
timestamp 1621523292
transform 1 0 1656 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_18
timestamp 1621523292
transform 1 0 2760 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1621523292
transform 1 0 3772 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_26
timestamp 1621523292
transform 1 0 3496 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_30
timestamp 1621523292
transform 1 0 3864 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_42
timestamp 1621523292
transform 1 0 4968 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_54
timestamp 1621523292
transform 1 0 6072 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1621523292
transform 1 0 9016 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_66
timestamp 1621523292
transform 1 0 7176 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_78
timestamp 1621523292
transform 1 0 8280 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_87
timestamp 1621523292
transform 1 0 9108 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_99
timestamp 1621523292
transform 1 0 10212 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_111
timestamp 1621523292
transform 1 0 11316 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_123
timestamp 1621523292
transform 1 0 12420 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _1838_
timestamp 1621523292
transform 1 0 14996 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1621523292
transform 1 0 14260 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_135
timestamp 1621523292
transform 1 0 13524 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_84_144
timestamp 1621523292
transform 1 0 14352 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_150
timestamp 1621523292
transform 1 0 14904 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 1621523292
transform 1 0 16192 0 -1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1841_
timestamp 1621523292
transform 1 0 17020 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_159
timestamp 1621523292
transform 1 0 15732 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_163
timestamp 1621523292
transform 1 0 16100 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_169
timestamp 1621523292
transform 1 0 16652 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1797_
timestamp 1621523292
transform 1 0 18400 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_176
timestamp 1621523292
transform 1 0 17296 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_196
timestamp 1621523292
transform 1 0 19136 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2346_
timestamp 1621523292
transform 1 0 20516 0 -1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1621523292
transform 1 0 19504 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_201
timestamp 1621523292
transform 1 0 19596 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_209
timestamp 1621523292
transform 1 0 20332 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_227
timestamp 1621523292
transform 1 0 21988 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_239
timestamp 1621523292
transform 1 0 23092 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1867_
timestamp 1621523292
transform 1 0 24104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1621523292
transform 1 0 24748 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_wb_clk_i
timestamp 1621523292
transform 1 0 23460 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_246
timestamp 1621523292
transform 1 0 23736 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_253
timestamp 1621523292
transform 1 0 24380 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_258
timestamp 1621523292
transform 1 0 24840 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2445_
timestamp 1621523292
transform 1 0 25576 0 -1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_84_282
timestamp 1621523292
transform 1 0 27048 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2068_
timestamp 1621523292
transform 1 0 28612 0 -1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2070_
timestamp 1621523292
transform 1 0 27692 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_288
timestamp 1621523292
transform 1 0 27600 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_295
timestamp 1621523292
transform 1 0 28244 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_304
timestamp 1621523292
transform 1 0 29072 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1968_
timestamp 1621523292
transform 1 0 30452 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1621523292
transform 1 0 29992 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_312
timestamp 1621523292
transform 1 0 29808 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_315
timestamp 1621523292
transform 1 0 30084 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_322
timestamp 1621523292
transform 1 0 30728 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1971_
timestamp 1621523292
transform 1 0 32200 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1976_
timestamp 1621523292
transform 1 0 31280 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_wb_clk_i
timestamp 1621523292
transform 1 0 32844 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_334
timestamp 1621523292
transform 1 0 31832 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_341
timestamp 1621523292
transform 1 0 32476 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_348
timestamp 1621523292
transform 1 0 33120 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2084_
timestamp 1621523292
transform 1 0 33580 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2087_
timestamp 1621523292
transform 1 0 34224 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1621523292
transform 1 0 35236 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_352
timestamp 1621523292
transform 1 0 33488 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_356
timestamp 1621523292
transform 1 0 33856 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_364
timestamp 1621523292
transform 1 0 34592 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_370
timestamp 1621523292
transform 1 0 35144 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_372
timestamp 1621523292
transform 1 0 35328 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_384
timestamp 1621523292
transform 1 0 36432 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_396
timestamp 1621523292
transform 1 0 37536 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_408
timestamp 1621523292
transform 1 0 38640 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1621523292
transform 1 0 40480 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_420
timestamp 1621523292
transform 1 0 39744 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_429
timestamp 1621523292
transform 1 0 40572 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_441
timestamp 1621523292
transform 1 0 41676 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_453
timestamp 1621523292
transform 1 0 42780 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_465
timestamp 1621523292
transform 1 0 43884 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_477
timestamp 1621523292
transform 1 0 44988 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1621523292
transform 1 0 45724 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_486
timestamp 1621523292
transform 1 0 45816 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_498
timestamp 1621523292
transform 1 0 46920 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_510
timestamp 1621523292
transform 1 0 48024 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_522
timestamp 1621523292
transform 1 0 49128 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1621523292
transform 1 0 50968 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_534
timestamp 1621523292
transform 1 0 50232 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_84_543
timestamp 1621523292
transform 1 0 51060 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_555
timestamp 1621523292
transform 1 0 52164 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_567
timestamp 1621523292
transform 1 0 53268 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_579
timestamp 1621523292
transform 1 0 54372 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2175_
timestamp 1621523292
transform 1 0 56856 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1621523292
transform 1 0 56212 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_591
timestamp 1621523292
transform 1 0 55476 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_84_600
timestamp 1621523292
transform 1 0 56304 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_609
timestamp 1621523292
transform 1 0 57132 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2324_
timestamp 1621523292
transform 1 0 57500 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1621523292
transform -1 0 58880 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_621
timestamp 1621523292
transform 1 0 58236 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1621523292
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1621523292
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1621523292
transform 1 0 1380 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1621523292
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1621523292
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_6
timestamp 1621523292
transform 1 0 1656 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 1621523292
transform 1 0 2760 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1621523292
transform 1 0 3772 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1621523292
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1621523292
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_26
timestamp 1621523292
transform 1 0 3496 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_30
timestamp 1621523292
transform 1 0 3864 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_42
timestamp 1621523292
transform 1 0 4968 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1621523292
transform 1 0 6348 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_51
timestamp 1621523292
transform 1 0 5796 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_58
timestamp 1621523292
transform 1 0 6440 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_54
timestamp 1621523292
transform 1 0 6072 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1621523292
transform 1 0 9016 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_70
timestamp 1621523292
transform 1 0 7544 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_82
timestamp 1621523292
transform 1 0 8648 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_66
timestamp 1621523292
transform 1 0 7176 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_78
timestamp 1621523292
transform 1 0 8280 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_87
timestamp 1621523292
transform 1 0 9108 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_94
timestamp 1621523292
transform 1 0 9752 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_106
timestamp 1621523292
transform 1 0 10856 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_99
timestamp 1621523292
transform 1 0 10212 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1621523292
transform 1 0 11592 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_115
timestamp 1621523292
transform 1 0 11684 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_127
timestamp 1621523292
transform 1 0 12788 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_111
timestamp 1621523292
transform 1 0 11316 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_123
timestamp 1621523292
transform 1 0 12420 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1621523292
transform 1 0 14260 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_139
timestamp 1621523292
transform 1 0 13892 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_151
timestamp 1621523292
transform 1 0 14996 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_135
timestamp 1621523292
transform 1 0 13524 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_144
timestamp 1621523292
transform 1 0 14352 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1621523292
transform 1 0 16836 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_163
timestamp 1621523292
transform 1 0 16100 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_172
timestamp 1621523292
transform 1 0 16928 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_156
timestamp 1621523292
transform 1 0 15456 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_168
timestamp 1621523292
transform 1 0 16560 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2345_
timestamp 1621523292
transform 1 0 18124 0 1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_85_184
timestamp 1621523292
transform 1 0 18032 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_180
timestamp 1621523292
transform 1 0 17664 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_192
timestamp 1621523292
transform 1 0 18768 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1798_
timestamp 1621523292
transform 1 0 20240 0 1 48416
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1800_
timestamp 1621523292
transform 1 0 21068 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1621523292
transform 1 0 19504 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_201
timestamp 1621523292
transform 1 0 19596 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_207
timestamp 1621523292
transform 1 0 20148 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_213
timestamp 1621523292
transform 1 0 20700 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_201
timestamp 1621523292
transform 1 0 19596 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_213
timestamp 1621523292
transform 1 0 20700 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1804_
timestamp 1621523292
transform 1 0 22356 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1805_
timestamp 1621523292
transform 1 0 21436 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1621523292
transform 1 0 22080 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_220
timestamp 1621523292
transform 1 0 21344 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_229
timestamp 1621523292
transform 1 0 22172 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_227
timestamp 1621523292
transform 1 0 21988 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_234
timestamp 1621523292
transform 1 0 22632 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_246
timestamp 1621523292
transform 1 0 23736 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_86_258
timestamp 1621523292
transform 1 0 24840 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_86_254
timestamp 1621523292
transform 1 0 24472 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_261
timestamp 1621523292
transform 1 0 25116 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_257
timestamp 1621523292
transform 1 0 24748 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_253
timestamp 1621523292
transform 1 0 24380 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1621523292
transform 1 0 24748 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _1870_
timestamp 1621523292
transform 1 0 25208 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1869_
timestamp 1621523292
transform 1 0 24840 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_241
timestamp 1621523292
transform 1 0 23276 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_1  _1871_
timestamp 1621523292
transform 1 0 26312 0 -1 49504
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1872_
timestamp 1621523292
transform 1 0 25484 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2065_
timestamp 1621523292
transform 1 0 26680 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_85_269
timestamp 1621523292
transform 1 0 25852 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_277
timestamp 1621523292
transform 1 0 26588 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_281
timestamp 1621523292
transform 1 0 26956 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_270
timestamp 1621523292
transform 1 0 25944 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_279
timestamp 1621523292
transform 1 0 26772 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_285
timestamp 1621523292
transform 1 0 27324 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_293
timestamp 1621523292
transform 1 0 28060 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_286
timestamp 1621523292
transform 1 0 27416 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1621523292
transform 1 0 27324 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2064_
timestamp 1621523292
transform 1 0 27784 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_86_302
timestamp 1621523292
transform 1 0 28888 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_300
timestamp 1621523292
transform 1 0 28704 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2067_
timestamp 1621523292
transform 1 0 28428 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2446_
timestamp 1621523292
transform 1 0 27416 0 -1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2411_
timestamp 1621523292
transform 1 0 29072 0 1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_1  _1973_
timestamp 1621523292
transform 1 0 30912 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2071_
timestamp 1621523292
transform 1 0 29256 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2412_
timestamp 1621523292
transform 1 0 31004 0 -1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1621523292
transform 1 0 29992 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_320
timestamp 1621523292
transform 1 0 30544 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_309
timestamp 1621523292
transform 1 0 29532 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_313
timestamp 1621523292
transform 1 0 29900 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_315
timestamp 1621523292
transform 1 0 30084 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_323
timestamp 1621523292
transform 1 0 30820 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1974_
timestamp 1621523292
transform 1 0 31832 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2337_
timestamp 1621523292
transform 1 0 33028 0 1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1621523292
transform 1 0 32568 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_330
timestamp 1621523292
transform 1 0 31464 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_337
timestamp 1621523292
transform 1 0 32108 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_341
timestamp 1621523292
transform 1 0 32476 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_343
timestamp 1621523292
transform 1 0 32660 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_341
timestamp 1621523292
transform 1 0 32476 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_349
timestamp 1621523292
transform 1 0 33212 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _2085_
timestamp 1621523292
transform 1 0 33304 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _2086_
timestamp 1621523292
transform 1 0 34408 0 -1 49504
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _2338_
timestamp 1621523292
transform 1 0 34868 0 1 48416
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1621523292
transform 1 0 35236 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_363
timestamp 1621523292
transform 1 0 34500 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_358
timestamp 1621523292
transform 1 0 34040 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_367
timestamp 1621523292
transform 1 0 34868 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_383
timestamp 1621523292
transform 1 0 36340 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_372
timestamp 1621523292
transform 1 0 35328 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_384
timestamp 1621523292
transform 1 0 36432 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1621523292
transform 1 0 37812 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_395
timestamp 1621523292
transform 1 0 37444 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_400
timestamp 1621523292
transform 1 0 37904 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_412
timestamp 1621523292
transform 1 0 39008 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_396
timestamp 1621523292
transform 1 0 37536 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_408
timestamp 1621523292
transform 1 0 38640 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1621523292
transform 1 0 40480 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_424
timestamp 1621523292
transform 1 0 40112 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_436
timestamp 1621523292
transform 1 0 41216 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_420
timestamp 1621523292
transform 1 0 39744 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_429
timestamp 1621523292
transform 1 0 40572 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1621523292
transform 1 0 43056 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_448
timestamp 1621523292
transform 1 0 42320 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_457
timestamp 1621523292
transform 1 0 43148 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_441
timestamp 1621523292
transform 1 0 41676 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_453
timestamp 1621523292
transform 1 0 42780 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_469
timestamp 1621523292
transform 1 0 44252 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_465
timestamp 1621523292
transform 1 0 43884 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_477
timestamp 1621523292
transform 1 0 44988 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1621523292
transform 1 0 45724 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_481
timestamp 1621523292
transform 1 0 45356 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_493
timestamp 1621523292
transform 1 0 46460 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_486
timestamp 1621523292
transform 1 0 45816 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_498
timestamp 1621523292
transform 1 0 46920 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1621523292
transform 1 0 48300 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_505
timestamp 1621523292
transform 1 0 47564 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_85_514
timestamp 1621523292
transform 1 0 48392 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_510
timestamp 1621523292
transform 1 0 48024 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_522
timestamp 1621523292
transform 1 0 49128 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1621523292
transform 1 0 50968 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_526
timestamp 1621523292
transform 1 0 49496 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_538
timestamp 1621523292
transform 1 0 50600 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_534
timestamp 1621523292
transform 1 0 50232 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_543
timestamp 1621523292
transform 1 0 51060 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_550
timestamp 1621523292
transform 1 0 51704 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_562
timestamp 1621523292
transform 1 0 52808 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_555
timestamp 1621523292
transform 1 0 52164 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_567
timestamp 1621523292
transform 1 0 53268 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1621523292
transform 1 0 53544 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_571
timestamp 1621523292
transform 1 0 53636 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_583
timestamp 1621523292
transform 1 0 54740 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_579
timestamp 1621523292
transform 1 0 54372 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_591
timestamp 1621523292
transform 1 0 55476 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_85_595
timestamp 1621523292
transform 1 0 55844 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_604
timestamp 1621523292
transform 1 0 56672 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_600
timestamp 1621523292
transform 1 0 56304 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_606
timestamp 1621523292
transform 1 0 56856 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output239
timestamp 1621523292
transform 1 0 56764 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1621523292
transform 1 0 56580 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1621523292
transform 1 0 56212 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_609
timestamp 1621523292
transform 1 0 57132 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2176_
timestamp 1621523292
transform 1 0 57224 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_1  _2325_
timestamp 1621523292
transform 1 0 57500 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1621523292
transform -1 0 58880 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1621523292
transform -1 0 58880 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output200
timestamp 1621523292
transform 1 0 57868 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_613
timestamp 1621523292
transform 1 0 57500 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1621523292
transform 1 0 58236 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_621
timestamp 1621523292
transform 1 0 58236 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1621523292
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1621523292
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1621523292
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1621523292
transform 1 0 3588 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1621523292
transform 1 0 4692 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1621523292
transform 1 0 6348 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_51
timestamp 1621523292
transform 1 0 5796 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_58
timestamp 1621523292
transform 1 0 6440 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_70
timestamp 1621523292
transform 1 0 7544 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_82
timestamp 1621523292
transform 1 0 8648 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_94
timestamp 1621523292
transform 1 0 9752 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_106
timestamp 1621523292
transform 1 0 10856 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1621523292
transform 1 0 11592 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_115
timestamp 1621523292
transform 1 0 11684 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_127
timestamp 1621523292
transform 1 0 12788 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_139
timestamp 1621523292
transform 1 0 13892 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_151
timestamp 1621523292
transform 1 0 14996 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1621523292
transform 1 0 16836 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_163
timestamp 1621523292
transform 1 0 16100 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_172
timestamp 1621523292
transform 1 0 16928 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_184
timestamp 1621523292
transform 1 0 18032 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_196
timestamp 1621523292
transform 1 0 19136 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2347_
timestamp 1621523292
transform 1 0 19412 0 1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_215
timestamp 1621523292
transform 1 0 20884 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1801_
timestamp 1621523292
transform 1 0 21252 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1803_
timestamp 1621523292
transform 1 0 22540 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1621523292
transform 1 0 22080 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_222
timestamp 1621523292
transform 1 0 21528 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_87_229
timestamp 1621523292
transform 1 0 22172 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_87_236
timestamp 1621523292
transform 1 0 22816 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2373_
timestamp 1621523292
transform 1 0 23552 0 1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_87_260
timestamp 1621523292
transform 1 0 25024 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2374_
timestamp 1621523292
transform 1 0 25484 0 1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_87_264
timestamp 1621523292
transform 1 0 25392 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_281
timestamp 1621523292
transform 1 0 26956 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2447_
timestamp 1621523292
transform 1 0 27784 0 1 49504
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1621523292
transform 1 0 27324 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_286
timestamp 1621523292
transform 1 0 27416 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1972_
timestamp 1621523292
transform 1 0 29992 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1977_
timestamp 1621523292
transform 1 0 31004 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_87_306
timestamp 1621523292
transform 1 0 29256 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_87_317
timestamp 1621523292
transform 1 0 30268 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1975_
timestamp 1621523292
transform 1 0 31648 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1980_
timestamp 1621523292
transform 1 0 33028 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1621523292
transform 1 0 32568 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_328
timestamp 1621523292
transform 1 0 31280 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_335
timestamp 1621523292
transform 1 0 31924 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_341
timestamp 1621523292
transform 1 0 32476 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_343
timestamp 1621523292
transform 1 0 32660 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2088_
timestamp 1621523292
transform 1 0 34500 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_wb_clk_i
timestamp 1621523292
transform 1 0 33672 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_350
timestamp 1621523292
transform 1 0 33304 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_357
timestamp 1621523292
transform 1 0 33948 0 1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_87_366
timestamp 1621523292
transform 1 0 34776 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_378
timestamp 1621523292
transform 1 0 35880 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_390
timestamp 1621523292
transform 1 0 36984 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1621523292
transform 1 0 37812 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_398
timestamp 1621523292
transform 1 0 37720 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_400
timestamp 1621523292
transform 1 0 37904 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_412
timestamp 1621523292
transform 1 0 39008 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_424
timestamp 1621523292
transform 1 0 40112 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_436
timestamp 1621523292
transform 1 0 41216 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1621523292
transform 1 0 43056 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_448
timestamp 1621523292
transform 1 0 42320 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_457
timestamp 1621523292
transform 1 0 43148 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_469
timestamp 1621523292
transform 1 0 44252 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_481
timestamp 1621523292
transform 1 0 45356 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_493
timestamp 1621523292
transform 1 0 46460 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1621523292
transform 1 0 48300 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_505
timestamp 1621523292
transform 1 0 47564 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_87_514
timestamp 1621523292
transform 1 0 48392 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_526
timestamp 1621523292
transform 1 0 49496 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_538
timestamp 1621523292
transform 1 0 50600 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_550
timestamp 1621523292
transform 1 0 51704 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_562
timestamp 1621523292
transform 1 0 52808 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1621523292
transform 1 0 53544 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_571
timestamp 1621523292
transform 1 0 53636 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_583
timestamp 1621523292
transform 1 0 54740 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1621523292
transform 1 0 57224 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_595
timestamp 1621523292
transform 1 0 55844 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_87_607
timestamp 1621523292
transform 1 0 56948 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1621523292
transform -1 0 58880 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output201
timestamp 1621523292
transform 1 0 57868 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_613
timestamp 1621523292
transform 1 0 57500 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_621
timestamp 1621523292
transform 1 0 58236 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1621523292
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1621523292
transform 1 0 1380 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_6
timestamp 1621523292
transform 1 0 1656 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 1621523292
transform 1 0 2760 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1621523292
transform 1 0 3772 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_26
timestamp 1621523292
transform 1 0 3496 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_30
timestamp 1621523292
transform 1 0 3864 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_42
timestamp 1621523292
transform 1 0 4968 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_54
timestamp 1621523292
transform 1 0 6072 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1621523292
transform 1 0 9016 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_66
timestamp 1621523292
transform 1 0 7176 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_78
timestamp 1621523292
transform 1 0 8280 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_87
timestamp 1621523292
transform 1 0 9108 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_99
timestamp 1621523292
transform 1 0 10212 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_111
timestamp 1621523292
transform 1 0 11316 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_123
timestamp 1621523292
transform 1 0 12420 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1621523292
transform 1 0 14260 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_135
timestamp 1621523292
transform 1 0 13524 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_144
timestamp 1621523292
transform 1 0 14352 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_156
timestamp 1621523292
transform 1 0 15456 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_168
timestamp 1621523292
transform 1 0 16560 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_180
timestamp 1621523292
transform 1 0 17664 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_192
timestamp 1621523292
transform 1 0 18768 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1802_
timestamp 1621523292
transform 1 0 20148 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2348_
timestamp 1621523292
transform 1 0 21160 0 -1 50592
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1621523292
transform 1 0 19504 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_88_201
timestamp 1621523292
transform 1 0 19596 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_213
timestamp 1621523292
transform 1 0 20700 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_217
timestamp 1621523292
transform 1 0 21068 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_234
timestamp 1621523292
transform 1 0 22632 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1621523292
transform 1 0 24748 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_wb_clk_i
timestamp 1621523292
transform 1 0 23920 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_246
timestamp 1621523292
transform 1 0 23736 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_88_251
timestamp 1621523292
transform 1 0 24196 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_88_258
timestamp 1621523292
transform 1 0 24840 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1873_
timestamp 1621523292
transform 1 0 25760 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_266
timestamp 1621523292
transform 1 0 25576 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_88_271
timestamp 1621523292
transform 1 0 26036 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_283
timestamp 1621523292
transform 1 0 27140 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2072_
timestamp 1621523292
transform 1 0 28796 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2073_
timestamp 1621523292
transform 1 0 27876 0 -1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_88_297
timestamp 1621523292
transform 1 0 28428 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_304
timestamp 1621523292
transform 1 0 29072 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2413_
timestamp 1621523292
transform 1 0 30452 0 -1 50592
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1621523292
transform 1 0 29992 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_312
timestamp 1621523292
transform 1 0 29808 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_315
timestamp 1621523292
transform 1 0 30084 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 32292 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_88_335
timestamp 1621523292
transform 1 0 31924 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_347
timestamp 1621523292
transform 1 0 33028 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2339_
timestamp 1621523292
transform 1 0 33396 0 -1 50592
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1621523292
transform 1 0 35236 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_367
timestamp 1621523292
transform 1 0 34868 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_372
timestamp 1621523292
transform 1 0 35328 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_384
timestamp 1621523292
transform 1 0 36432 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_396
timestamp 1621523292
transform 1 0 37536 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_408
timestamp 1621523292
transform 1 0 38640 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1621523292
transform 1 0 40480 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_420
timestamp 1621523292
transform 1 0 39744 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_429
timestamp 1621523292
transform 1 0 40572 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_441
timestamp 1621523292
transform 1 0 41676 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_453
timestamp 1621523292
transform 1 0 42780 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_465
timestamp 1621523292
transform 1 0 43884 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_477
timestamp 1621523292
transform 1 0 44988 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1621523292
transform 1 0 45724 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_486
timestamp 1621523292
transform 1 0 45816 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_498
timestamp 1621523292
transform 1 0 46920 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_510
timestamp 1621523292
transform 1 0 48024 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_522
timestamp 1621523292
transform 1 0 49128 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1621523292
transform 1 0 50968 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_534
timestamp 1621523292
transform 1 0 50232 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_543
timestamp 1621523292
transform 1 0 51060 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_555
timestamp 1621523292
transform 1 0 52164 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_567
timestamp 1621523292
transform 1 0 53268 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_579
timestamp 1621523292
transform 1 0 54372 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1621523292
transform 1 0 56212 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1621523292
transform 1 0 57224 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_88_591
timestamp 1621523292
transform 1 0 55476 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_88_600
timestamp 1621523292
transform 1 0 56304 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_608
timestamp 1621523292
transform 1 0 57040 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1621523292
transform -1 0 58880 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output240
timestamp 1621523292
transform 1 0 57868 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_613
timestamp 1621523292
transform 1 0 57500 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_621
timestamp 1621523292
transform 1 0 58236 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1621523292
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1621523292
transform 1 0 1380 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1621523292
transform 1 0 2484 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1621523292
transform 1 0 3588 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1621523292
transform 1 0 4692 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1621523292
transform 1 0 6348 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_51
timestamp 1621523292
transform 1 0 5796 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_89_58
timestamp 1621523292
transform 1 0 6440 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_70
timestamp 1621523292
transform 1 0 7544 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_82
timestamp 1621523292
transform 1 0 8648 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_94
timestamp 1621523292
transform 1 0 9752 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_106
timestamp 1621523292
transform 1 0 10856 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1621523292
transform 1 0 11592 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_115
timestamp 1621523292
transform 1 0 11684 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_127
timestamp 1621523292
transform 1 0 12788 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_139
timestamp 1621523292
transform 1 0 13892 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_151
timestamp 1621523292
transform 1 0 14996 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1621523292
transform 1 0 16836 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_163
timestamp 1621523292
transform 1 0 16100 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_172
timestamp 1621523292
transform 1 0 16928 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_184
timestamp 1621523292
transform 1 0 18032 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_196
timestamp 1621523292
transform 1 0 19136 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1807_
timestamp 1621523292
transform 1 0 20792 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_89_208
timestamp 1621523292
transform 1 0 20240 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_89_217
timestamp 1621523292
transform 1 0 21068 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1806_
timestamp 1621523292
transform 1 0 21436 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1621523292
transform 1 0 22080 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_wb_clk_i
timestamp 1621523292
transform 1 0 22632 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_224
timestamp 1621523292
transform 1 0 21712 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_229
timestamp 1621523292
transform 1 0 22172 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_233
timestamp 1621523292
transform 1 0 22540 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_237
timestamp 1621523292
transform 1 0 22908 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__o2bb2a_1  _1874_
timestamp 1621523292
transform 1 0 25024 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_89_249
timestamp 1621523292
transform 1 0 24012 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_257
timestamp 1621523292
transform 1 0 24748 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1876_
timestamp 1621523292
transform 1 0 26128 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_268
timestamp 1621523292
transform 1 0 25760 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_276
timestamp 1621523292
transform 1 0 26496 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2074_
timestamp 1621523292
transform 1 0 28152 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2075_
timestamp 1621523292
transform 1 0 28796 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1621523292
transform 1 0 27324 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_284
timestamp 1621523292
transform 1 0 27232 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_286
timestamp 1621523292
transform 1 0 27416 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_89_297
timestamp 1621523292
transform 1 0 28428 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_304
timestamp 1621523292
transform 1 0 29072 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2077_
timestamp 1621523292
transform 1 0 29440 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2078_
timestamp 1621523292
transform 1 0 30452 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_311
timestamp 1621523292
transform 1 0 29716 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_89_322
timestamp 1621523292
transform 1 0 30728 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1978_
timestamp 1621523292
transform 1 0 33028 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1979_
timestamp 1621523292
transform 1 0 31372 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1621523292
transform 1 0 32568 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_89_328
timestamp 1621523292
transform 1 0 31280 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_89_335
timestamp 1621523292
transform 1 0 31924 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_341
timestamp 1621523292
transform 1 0 32476 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_343
timestamp 1621523292
transform 1 0 32660 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2089_
timestamp 1621523292
transform 1 0 35052 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2090_
timestamp 1621523292
transform 1 0 34132 0 1 50592
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_89_350
timestamp 1621523292
transform 1 0 33304 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_358
timestamp 1621523292
transform 1 0 34040 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_365
timestamp 1621523292
transform 1 0 34684 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2091_
timestamp 1621523292
transform 1 0 35696 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_372
timestamp 1621523292
transform 1 0 35328 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_379
timestamp 1621523292
transform 1 0 35972 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_391
timestamp 1621523292
transform 1 0 37076 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1621523292
transform 1 0 37812 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_400
timestamp 1621523292
transform 1 0 37904 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_412
timestamp 1621523292
transform 1 0 39008 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_424
timestamp 1621523292
transform 1 0 40112 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_436
timestamp 1621523292
transform 1 0 41216 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1621523292
transform 1 0 43056 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_448
timestamp 1621523292
transform 1 0 42320 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_457
timestamp 1621523292
transform 1 0 43148 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_469
timestamp 1621523292
transform 1 0 44252 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_481
timestamp 1621523292
transform 1 0 45356 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_493
timestamp 1621523292
transform 1 0 46460 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1621523292
transform 1 0 48300 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_505
timestamp 1621523292
transform 1 0 47564 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_514
timestamp 1621523292
transform 1 0 48392 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_526
timestamp 1621523292
transform 1 0 49496 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_538
timestamp 1621523292
transform 1 0 50600 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_550
timestamp 1621523292
transform 1 0 51704 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_562
timestamp 1621523292
transform 1 0 52808 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1621523292
transform 1 0 53544 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_571
timestamp 1621523292
transform 1 0 53636 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_583
timestamp 1621523292
transform 1 0 54740 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1549_
timestamp 1621523292
transform 1 0 56856 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_89_595
timestamp 1621523292
transform 1 0 55844 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_603
timestamp 1621523292
transform 1 0 56580 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_609
timestamp 1621523292
transform 1 0 57132 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2326_
timestamp 1621523292
transform 1 0 57500 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1621523292
transform -1 0 58880 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_621
timestamp 1621523292
transform 1 0 58236 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1621523292
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1621523292
transform 1 0 1380 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_6
timestamp 1621523292
transform 1 0 1656 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_18
timestamp 1621523292
transform 1 0 2760 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1621523292
transform 1 0 3772 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_26
timestamp 1621523292
transform 1 0 3496 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_30
timestamp 1621523292
transform 1 0 3864 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_42
timestamp 1621523292
transform 1 0 4968 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_54
timestamp 1621523292
transform 1 0 6072 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1621523292
transform 1 0 9016 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_66
timestamp 1621523292
transform 1 0 7176 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_78
timestamp 1621523292
transform 1 0 8280 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_87
timestamp 1621523292
transform 1 0 9108 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_99
timestamp 1621523292
transform 1 0 10212 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_111
timestamp 1621523292
transform 1 0 11316 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_123
timestamp 1621523292
transform 1 0 12420 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1621523292
transform 1 0 14260 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_135
timestamp 1621523292
transform 1 0 13524 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_144
timestamp 1621523292
transform 1 0 14352 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_156
timestamp 1621523292
transform 1 0 15456 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_168
timestamp 1621523292
transform 1 0 16560 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_180
timestamp 1621523292
transform 1 0 17664 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_192
timestamp 1621523292
transform 1 0 18768 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2349_
timestamp 1621523292
transform 1 0 20424 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1621523292
transform 1 0 19504 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_201
timestamp 1621523292
transform 1 0 19596 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_209
timestamp 1621523292
transform 1 0 20332 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2377_
timestamp 1621523292
transform 1 0 22264 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_226
timestamp 1621523292
transform 1 0 21896 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1878_
timestamp 1621523292
transform 1 0 24104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1621523292
transform 1 0 24748 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_246
timestamp 1621523292
transform 1 0 23736 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_253
timestamp 1621523292
transform 1 0 24380 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_258
timestamp 1621523292
transform 1 0 24840 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2376_
timestamp 1621523292
transform 1 0 25392 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_280
timestamp 1621523292
transform 1 0 26864 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2079_
timestamp 1621523292
transform 1 0 29072 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2448_
timestamp 1621523292
transform 1 0 27232 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_90_300
timestamp 1621523292
transform 1 0 28704 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1486_
timestamp 1621523292
transform 1 0 30912 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1621523292
transform 1 0 29992 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_310
timestamp 1621523292
transform 1 0 29624 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_315
timestamp 1621523292
transform 1 0 30084 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_323
timestamp 1621523292
transform 1 0 30820 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2414_
timestamp 1621523292
transform 1 0 32016 0 -1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_90_328
timestamp 1621523292
transform 1 0 31280 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2080_
timestamp 1621523292
transform 1 0 33856 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1621523292
transform 1 0 35236 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_352
timestamp 1621523292
transform 1 0 33488 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_359
timestamp 1621523292
transform 1 0 34132 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_372
timestamp 1621523292
transform 1 0 35328 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_384
timestamp 1621523292
transform 1 0 36432 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_396
timestamp 1621523292
transform 1 0 37536 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_408
timestamp 1621523292
transform 1 0 38640 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1621523292
transform 1 0 40480 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_420
timestamp 1621523292
transform 1 0 39744 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_429
timestamp 1621523292
transform 1 0 40572 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_441
timestamp 1621523292
transform 1 0 41676 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_453
timestamp 1621523292
transform 1 0 42780 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_465
timestamp 1621523292
transform 1 0 43884 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_477
timestamp 1621523292
transform 1 0 44988 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1621523292
transform 1 0 45724 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_486
timestamp 1621523292
transform 1 0 45816 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_498
timestamp 1621523292
transform 1 0 46920 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_510
timestamp 1621523292
transform 1 0 48024 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_522
timestamp 1621523292
transform 1 0 49128 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1621523292
transform 1 0 50968 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_534
timestamp 1621523292
transform 1 0 50232 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_90_543
timestamp 1621523292
transform 1 0 51060 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_555
timestamp 1621523292
transform 1 0 52164 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_567
timestamp 1621523292
transform 1 0 53268 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_579
timestamp 1621523292
transform 1 0 54372 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _2177_
timestamp 1621523292
transform 1 0 57224 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1621523292
transform 1 0 56212 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_591
timestamp 1621523292
transform 1 0 55476 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_90_600
timestamp 1621523292
transform 1 0 56304 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_608
timestamp 1621523292
transform 1 0 57040 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1621523292
transform -1 0 58880 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output202
timestamp 1621523292
transform 1 0 57868 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1621523292
transform 1 0 57500 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_621
timestamp 1621523292
transform 1 0 58236 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1621523292
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1621523292
transform 1 0 1380 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_6
timestamp 1621523292
transform 1 0 1656 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_18
timestamp 1621523292
transform 1 0 2760 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_30
timestamp 1621523292
transform 1 0 3864 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_42
timestamp 1621523292
transform 1 0 4968 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1621523292
transform 1 0 6348 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_54
timestamp 1621523292
transform 1 0 6072 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_58
timestamp 1621523292
transform 1 0 6440 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_70
timestamp 1621523292
transform 1 0 7544 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_82
timestamp 1621523292
transform 1 0 8648 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_94
timestamp 1621523292
transform 1 0 9752 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_106
timestamp 1621523292
transform 1 0 10856 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1621523292
transform 1 0 11592 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_115
timestamp 1621523292
transform 1 0 11684 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_127
timestamp 1621523292
transform 1 0 12788 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_139
timestamp 1621523292
transform 1 0 13892 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_151
timestamp 1621523292
transform 1 0 14996 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1621523292
transform 1 0 16836 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_163
timestamp 1621523292
transform 1 0 16100 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_172
timestamp 1621523292
transform 1 0 16928 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_184
timestamp 1621523292
transform 1 0 18032 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_196
timestamp 1621523292
transform 1 0 19136 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1808_
timestamp 1621523292
transform 1 0 21068 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_91_208
timestamp 1621523292
transform 1 0 20240 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_216
timestamp 1621523292
transform 1 0 20976 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1879_
timestamp 1621523292
transform 1 0 22908 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1621523292
transform 1 0 22080 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_223
timestamp 1621523292
transform 1 0 21620 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_227
timestamp 1621523292
transform 1 0 21988 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_229
timestamp 1621523292
transform 1 0 22172 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2375_
timestamp 1621523292
transform 1 0 23920 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_243
timestamp 1621523292
transform 1 0 23460 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_247
timestamp 1621523292
transform 1 0 23828 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__and3_1  _1875_
timestamp 1621523292
transform 1 0 25760 0 1 51680
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_wb_clk_i
timestamp 1621523292
transform 1 0 26588 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_264
timestamp 1621523292
transform 1 0 25392 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_273
timestamp 1621523292
transform 1 0 26220 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_280
timestamp 1621523292
transform 1 0 26864 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2076_
timestamp 1621523292
transform 1 0 27784 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2081_
timestamp 1621523292
transform 1 0 28888 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1621523292
transform 1 0 27324 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_284
timestamp 1621523292
transform 1 0 27232 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_286
timestamp 1621523292
transform 1 0 27416 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_91_296
timestamp 1621523292
transform 1 0 28336 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2450_
timestamp 1621523292
transform 1 0 29992 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_310
timestamp 1621523292
transform 1 0 29624 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1485_
timestamp 1621523292
transform 1 0 31832 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 33028 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1621523292
transform 1 0 32568 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_330
timestamp 1621523292
transform 1 0 31464 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_338
timestamp 1621523292
transform 1 0 32200 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_343
timestamp 1621523292
transform 1 0 32660 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2340_
timestamp 1621523292
transform 1 0 34316 0 1 51680
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_91_356
timestamp 1621523292
transform 1 0 33856 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_360
timestamp 1621523292
transform 1 0 34224 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _2092_
timestamp 1621523292
transform 1 0 36156 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_377
timestamp 1621523292
transform 1 0 35788 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_384
timestamp 1621523292
transform 1 0 36432 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1621523292
transform 1 0 37812 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_396
timestamp 1621523292
transform 1 0 37536 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_400
timestamp 1621523292
transform 1 0 37904 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_412
timestamp 1621523292
transform 1 0 39008 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_424
timestamp 1621523292
transform 1 0 40112 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_436
timestamp 1621523292
transform 1 0 41216 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1621523292
transform 1 0 43056 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_448
timestamp 1621523292
transform 1 0 42320 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_457
timestamp 1621523292
transform 1 0 43148 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_469
timestamp 1621523292
transform 1 0 44252 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_481
timestamp 1621523292
transform 1 0 45356 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_493
timestamp 1621523292
transform 1 0 46460 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1621523292
transform 1 0 48300 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_505
timestamp 1621523292
transform 1 0 47564 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_514
timestamp 1621523292
transform 1 0 48392 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_526
timestamp 1621523292
transform 1 0 49496 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_538
timestamp 1621523292
transform 1 0 50600 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_550
timestamp 1621523292
transform 1 0 51704 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_562
timestamp 1621523292
transform 1 0 52808 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1621523292
transform 1 0 53544 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_571
timestamp 1621523292
transform 1 0 53636 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_583
timestamp 1621523292
transform 1 0 54740 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1621523292
transform 1 0 57224 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1621523292
transform 1 0 56580 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_91_595
timestamp 1621523292
transform 1 0 55844 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_91_606
timestamp 1621523292
transform 1 0 56856 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1621523292
transform -1 0 58880 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output241
timestamp 1621523292
transform 1 0 57868 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_613
timestamp 1621523292
transform 1 0 57500 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_621
timestamp 1621523292
transform 1 0 58236 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1621523292
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1621523292
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1621523292
transform 1 0 1380 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1621523292
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1621523292
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_6
timestamp 1621523292
transform 1 0 1656 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_18
timestamp 1621523292
transform 1 0 2760 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1621523292
transform 1 0 3772 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_27
timestamp 1621523292
transform 1 0 3588 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_30
timestamp 1621523292
transform 1 0 3864 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_42
timestamp 1621523292
transform 1 0 4968 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_30
timestamp 1621523292
transform 1 0 3864 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_42
timestamp 1621523292
transform 1 0 4968 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1621523292
transform 1 0 6348 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_54
timestamp 1621523292
transform 1 0 6072 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_54
timestamp 1621523292
transform 1 0 6072 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_58
timestamp 1621523292
transform 1 0 6440 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1621523292
transform 1 0 9016 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_66
timestamp 1621523292
transform 1 0 7176 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_78
timestamp 1621523292
transform 1 0 8280 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_87
timestamp 1621523292
transform 1 0 9108 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_70
timestamp 1621523292
transform 1 0 7544 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_82
timestamp 1621523292
transform 1 0 8648 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_99
timestamp 1621523292
transform 1 0 10212 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_94
timestamp 1621523292
transform 1 0 9752 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_106
timestamp 1621523292
transform 1 0 10856 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1621523292
transform 1 0 11592 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_111
timestamp 1621523292
transform 1 0 11316 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_123
timestamp 1621523292
transform 1 0 12420 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_115
timestamp 1621523292
transform 1 0 11684 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_127
timestamp 1621523292
transform 1 0 12788 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1621523292
transform 1 0 14260 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_135
timestamp 1621523292
transform 1 0 13524 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_144
timestamp 1621523292
transform 1 0 14352 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_139
timestamp 1621523292
transform 1 0 13892 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_151
timestamp 1621523292
transform 1 0 14996 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1621523292
transform 1 0 16836 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_156
timestamp 1621523292
transform 1 0 15456 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_168
timestamp 1621523292
transform 1 0 16560 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_163
timestamp 1621523292
transform 1 0 16100 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_172
timestamp 1621523292
transform 1 0 16928 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_180
timestamp 1621523292
transform 1 0 17664 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_192
timestamp 1621523292
transform 1 0 18768 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_184
timestamp 1621523292
transform 1 0 18032 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_196
timestamp 1621523292
transform 1 0 19136 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1809_
timestamp 1621523292
transform 1 0 21068 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1621523292
transform 1 0 19504 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_201
timestamp 1621523292
transform 1 0 19596 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_213
timestamp 1621523292
transform 1 0 20700 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_208
timestamp 1621523292
transform 1 0 20240 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_229
timestamp 1621523292
transform 1 0 22172 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_224
timestamp 1621523292
transform 1 0 21712 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_220
timestamp 1621523292
transform 1 0 21344 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_220
timestamp 1621523292
transform 1 0 21344 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1621523292
transform 1 0 22080 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _1811_
timestamp 1621523292
transform 1 0 21712 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1810_
timestamp 1621523292
transform 1 0 21436 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_93_235
timestamp 1621523292
transform 1 0 22724 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_240
timestamp 1621523292
transform 1 0 23184 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_236
timestamp 1621523292
transform 1 0 22816 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_230
timestamp 1621523292
transform 1 0 22264 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1881_
timestamp 1621523292
transform 1 0 22908 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2378_
timestamp 1621523292
transform 1 0 22816 0 1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1880_
timestamp 1621523292
transform 1 0 23552 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2379_
timestamp 1621523292
transform 1 0 24656 0 1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1621523292
transform 1 0 24748 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_247
timestamp 1621523292
transform 1 0 23828 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_255
timestamp 1621523292
transform 1 0 24564 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_258
timestamp 1621523292
transform 1 0 24840 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_252
timestamp 1621523292
transform 1 0 24288 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1877_
timestamp 1621523292
transform 1 0 25668 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1884_
timestamp 1621523292
transform 1 0 26496 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_92_266
timestamp 1621523292
transform 1 0 25576 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_270
timestamp 1621523292
transform 1 0 25944 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_282
timestamp 1621523292
transform 1 0 27048 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_272
timestamp 1621523292
transform 1 0 26128 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_93_279
timestamp 1621523292
transform 1 0 26772 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1889_
timestamp 1621523292
transform 1 0 27876 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1892_
timestamp 1621523292
transform 1 0 29164 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2449_
timestamp 1621523292
transform 1 0 28152 0 -1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1621523292
transform 1 0 27324 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_286
timestamp 1621523292
transform 1 0 27416 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_290
timestamp 1621523292
transform 1 0 27784 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_294
timestamp 1621523292
transform 1 0 28152 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_93_302
timestamp 1621523292
transform 1 0 28888 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_308
timestamp 1621523292
transform 1 0 29440 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_310
timestamp 1621523292
transform 1 0 29624 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1621523292
transform 1 0 29992 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _1890_
timestamp 1621523292
transform 1 0 29808 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_93_315
timestamp 1621523292
transform 1 0 30084 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_319
timestamp 1621523292
transform 1 0 30452 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_315
timestamp 1621523292
transform 1 0 30084 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1621523292
transform 1 0 30544 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1493_
timestamp 1621523292
transform 1 0 30452 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_327
timestamp 1621523292
transform 1 0 31188 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_338
timestamp 1621523292
transform 1 0 32200 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_331
timestamp 1621523292
transform 1 0 31556 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_328
timestamp 1621523292
transform 1 0 31280 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2190_
timestamp 1621523292
transform 1 0 31648 0 -1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1791_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 31648 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_343
timestamp 1621523292
transform 1 0 32660 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_341
timestamp 1621523292
transform 1 0 32476 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1621523292
transform 1 0 32568 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1487_
timestamp 1621523292
transform 1 0 33028 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2486_
timestamp 1621523292
transform 1 0 32844 0 -1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2341_
timestamp 1621523292
transform 1 0 34684 0 1 52768
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1621523292
transform 1 0 35236 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_361
timestamp 1621523292
transform 1 0 34316 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_369
timestamp 1621523292
transform 1 0 35052 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_356
timestamp 1621523292
transform 1 0 33856 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_364
timestamp 1621523292
transform 1 0 34592 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _2093_
timestamp 1621523292
transform 1 0 35696 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2094_
timestamp 1621523292
transform 1 0 36616 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_372
timestamp 1621523292
transform 1 0 35328 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_382
timestamp 1621523292
transform 1 0 36248 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_389
timestamp 1621523292
transform 1 0 36892 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_381
timestamp 1621523292
transform 1 0 36156 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_393
timestamp 1621523292
transform 1 0 37260 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1621523292
transform 1 0 37812 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_401
timestamp 1621523292
transform 1 0 37996 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_413
timestamp 1621523292
transform 1 0 39100 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_400
timestamp 1621523292
transform 1 0 37904 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_412
timestamp 1621523292
transform 1 0 39008 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1621523292
transform 1 0 40480 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_425
timestamp 1621523292
transform 1 0 40204 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_429
timestamp 1621523292
transform 1 0 40572 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_424
timestamp 1621523292
transform 1 0 40112 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_436
timestamp 1621523292
transform 1 0 41216 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1621523292
transform 1 0 43056 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_441
timestamp 1621523292
transform 1 0 41676 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_453
timestamp 1621523292
transform 1 0 42780 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_448
timestamp 1621523292
transform 1 0 42320 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_457
timestamp 1621523292
transform 1 0 43148 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_465
timestamp 1621523292
transform 1 0 43884 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_477
timestamp 1621523292
transform 1 0 44988 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_469
timestamp 1621523292
transform 1 0 44252 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1621523292
transform 1 0 45724 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_486
timestamp 1621523292
transform 1 0 45816 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_498
timestamp 1621523292
transform 1 0 46920 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_481
timestamp 1621523292
transform 1 0 45356 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_493
timestamp 1621523292
transform 1 0 46460 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1621523292
transform 1 0 48300 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_510
timestamp 1621523292
transform 1 0 48024 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_522
timestamp 1621523292
transform 1 0 49128 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_505
timestamp 1621523292
transform 1 0 47564 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_514
timestamp 1621523292
transform 1 0 48392 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1621523292
transform 1 0 50968 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_534
timestamp 1621523292
transform 1 0 50232 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_543
timestamp 1621523292
transform 1 0 51060 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_526
timestamp 1621523292
transform 1 0 49496 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_538
timestamp 1621523292
transform 1 0 50600 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_555
timestamp 1621523292
transform 1 0 52164 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_567
timestamp 1621523292
transform 1 0 53268 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_550
timestamp 1621523292
transform 1 0 51704 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_562
timestamp 1621523292
transform 1 0 52808 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1621523292
transform 1 0 53544 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_579
timestamp 1621523292
transform 1 0 54372 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_571
timestamp 1621523292
transform 1 0 53636 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_583
timestamp 1621523292
transform 1 0 54740 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _1547_
timestamp 1621523292
transform 1 0 57224 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2178_
timestamp 1621523292
transform 1 0 56856 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1621523292
transform 1 0 56212 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1621523292
transform 1 0 56580 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_92_591
timestamp 1621523292
transform 1 0 55476 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_92_600
timestamp 1621523292
transform 1 0 56304 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_609
timestamp 1621523292
transform 1 0 57132 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_93_595
timestamp 1621523292
transform 1 0 55844 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_606
timestamp 1621523292
transform 1 0 56856 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2327_
timestamp 1621523292
transform 1 0 57500 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1621523292
transform -1 0 58880 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1621523292
transform -1 0 58880 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output203
timestamp 1621523292
transform 1 0 57868 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1621523292
transform 1 0 58236 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_613
timestamp 1621523292
transform 1 0 57500 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_621
timestamp 1621523292
transform 1 0 58236 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1621523292
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1621523292
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1621523292
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1621523292
transform 1 0 3772 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_27
timestamp 1621523292
transform 1 0 3588 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_30
timestamp 1621523292
transform 1 0 3864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_42
timestamp 1621523292
transform 1 0 4968 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_54
timestamp 1621523292
transform 1 0 6072 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1621523292
transform 1 0 9016 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_66
timestamp 1621523292
transform 1 0 7176 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_78
timestamp 1621523292
transform 1 0 8280 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_87
timestamp 1621523292
transform 1 0 9108 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_99
timestamp 1621523292
transform 1 0 10212 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_111
timestamp 1621523292
transform 1 0 11316 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_123
timestamp 1621523292
transform 1 0 12420 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1621523292
transform 1 0 14260 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_135
timestamp 1621523292
transform 1 0 13524 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_144
timestamp 1621523292
transform 1 0 14352 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_156
timestamp 1621523292
transform 1 0 15456 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_168
timestamp 1621523292
transform 1 0 16560 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_180
timestamp 1621523292
transform 1 0 17664 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_192
timestamp 1621523292
transform 1 0 18768 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2350_
timestamp 1621523292
transform 1 0 21160 0 -1 53856
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1621523292
transform 1 0 19504 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_201
timestamp 1621523292
transform 1 0 19596 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_213
timestamp 1621523292
transform 1 0 20700 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_217
timestamp 1621523292
transform 1 0 21068 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_234
timestamp 1621523292
transform 1 0 22632 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1882_
timestamp 1621523292
transform 1 0 23460 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1885_
timestamp 1621523292
transform 1 0 25208 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1621523292
transform 1 0 24748 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_242
timestamp 1621523292
transform 1 0 23368 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_249
timestamp 1621523292
transform 1 0 24012 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_258
timestamp 1621523292
transform 1 0 24840 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2380_
timestamp 1621523292
transform 1 0 26312 0 -1 53856
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_94_268
timestamp 1621523292
transform 1 0 25760 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2381_
timestamp 1621523292
transform 1 0 28152 0 -1 53856
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_290
timestamp 1621523292
transform 1 0 27784 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2481_
timestamp 1621523292
transform 1 0 30636 0 -1 53856
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1621523292
transform 1 0 29992 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_310
timestamp 1621523292
transform 1 0 29624 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_315
timestamp 1621523292
transform 1 0 30084 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1484_
timestamp 1621523292
transform 1 0 32476 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2485_
timestamp 1621523292
transform 1 0 33120 0 -1 53856
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_94_337
timestamp 1621523292
transform 1 0 32108 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_344
timestamp 1621523292
transform 1 0 32752 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1621523292
transform 1 0 35236 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_364
timestamp 1621523292
transform 1 0 34592 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_370
timestamp 1621523292
transform 1 0 35144 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_1  _2096_
timestamp 1621523292
transform 1 0 35696 0 -1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_94_372
timestamp 1621523292
transform 1 0 35328 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_382
timestamp 1621523292
transform 1 0 36248 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_394
timestamp 1621523292
transform 1 0 37352 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_406
timestamp 1621523292
transform 1 0 38456 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1621523292
transform 1 0 40480 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_418
timestamp 1621523292
transform 1 0 39560 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_426
timestamp 1621523292
transform 1 0 40296 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_429
timestamp 1621523292
transform 1 0 40572 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_441
timestamp 1621523292
transform 1 0 41676 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_453
timestamp 1621523292
transform 1 0 42780 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_465
timestamp 1621523292
transform 1 0 43884 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_477
timestamp 1621523292
transform 1 0 44988 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1621523292
transform 1 0 45724 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_486
timestamp 1621523292
transform 1 0 45816 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_498
timestamp 1621523292
transform 1 0 46920 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_510
timestamp 1621523292
transform 1 0 48024 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_522
timestamp 1621523292
transform 1 0 49128 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1621523292
transform 1 0 50968 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_534
timestamp 1621523292
transform 1 0 50232 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_94_543
timestamp 1621523292
transform 1 0 51060 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_555
timestamp 1621523292
transform 1 0 52164 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_567
timestamp 1621523292
transform 1 0 53268 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_579
timestamp 1621523292
transform 1 0 54372 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1621523292
transform 1 0 56212 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1621523292
transform 1 0 55568 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output242
timestamp 1621523292
transform 1 0 56764 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_591
timestamp 1621523292
transform 1 0 55476 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_595
timestamp 1621523292
transform 1 0 55844 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_600
timestamp 1621523292
transform 1 0 56304 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_604
timestamp 1621523292
transform 1 0 56672 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_609
timestamp 1621523292
transform 1 0 57132 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2328_
timestamp 1621523292
transform 1 0 57500 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1621523292
transform -1 0 58880 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_621
timestamp 1621523292
transform 1 0 58236 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1621523292
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1621523292
transform 1 0 1380 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_6
timestamp 1621523292
transform 1 0 1656 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_18
timestamp 1621523292
transform 1 0 2760 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_30
timestamp 1621523292
transform 1 0 3864 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_42
timestamp 1621523292
transform 1 0 4968 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1621523292
transform 1 0 6348 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_54
timestamp 1621523292
transform 1 0 6072 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_58
timestamp 1621523292
transform 1 0 6440 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_70
timestamp 1621523292
transform 1 0 7544 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_82
timestamp 1621523292
transform 1 0 8648 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_94
timestamp 1621523292
transform 1 0 9752 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_106
timestamp 1621523292
transform 1 0 10856 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1621523292
transform 1 0 11592 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_115
timestamp 1621523292
transform 1 0 11684 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_127
timestamp 1621523292
transform 1 0 12788 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_139
timestamp 1621523292
transform 1 0 13892 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_151
timestamp 1621523292
transform 1 0 14996 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1621523292
transform 1 0 16836 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_163
timestamp 1621523292
transform 1 0 16100 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_172
timestamp 1621523292
transform 1 0 16928 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_184
timestamp 1621523292
transform 1 0 18032 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_196
timestamp 1621523292
transform 1 0 19136 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_208
timestamp 1621523292
transform 1 0 20240 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1812_
timestamp 1621523292
transform 1 0 22540 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1813_
timestamp 1621523292
transform 1 0 23184 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1621523292
transform 1 0 22080 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_220
timestamp 1621523292
transform 1 0 21344 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_229
timestamp 1621523292
transform 1 0 22172 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_236
timestamp 1621523292
transform 1 0 22816 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1815_
timestamp 1621523292
transform 1 0 23828 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1816_
timestamp 1621523292
transform 1 0 24472 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1883_
timestamp 1621523292
transform 1 0 25116 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_243
timestamp 1621523292
transform 1 0 23460 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_250
timestamp 1621523292
transform 1 0 24104 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_257
timestamp 1621523292
transform 1 0 24748 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1886_
timestamp 1621523292
transform 1 0 25760 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1888_
timestamp 1621523292
transform 1 0 26404 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_264
timestamp 1621523292
transform 1 0 25392 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_271
timestamp 1621523292
transform 1 0 26036 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_281
timestamp 1621523292
transform 1 0 26956 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1887_
timestamp 1621523292
transform 1 0 27784 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1893_
timestamp 1621523292
transform 1 0 28980 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1621523292
transform 1 0 27324 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_286
timestamp 1621523292
transform 1 0 27416 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_293
timestamp 1621523292
transform 1 0 28060 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_301
timestamp 1621523292
transform 1 0 28796 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1621523292
transform 1 0 30360 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_95_311
timestamp 1621523292
transform 1 0 29716 0 1 53856
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_317
timestamp 1621523292
transform 1 0 30268 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_326
timestamp 1621523292
transform 1 0 31096 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1488_
timestamp 1621523292
transform 1 0 33028 0 1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1621523292
transform 1 0 32568 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1621523292
transform 1 0 31464 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_338
timestamp 1621523292
transform 1 0 32200 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_343
timestamp 1621523292
transform 1 0 32660 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _2098_
timestamp 1621523292
transform 1 0 35236 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_356
timestamp 1621523292
transform 1 0 33856 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_368
timestamp 1621523292
transform 1 0 34960 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2095_
timestamp 1621523292
transform 1 0 36340 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_379
timestamp 1621523292
transform 1 0 35972 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_386
timestamp 1621523292
transform 1 0 36616 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1621523292
transform 1 0 37812 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_398
timestamp 1621523292
transform 1 0 37720 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_400
timestamp 1621523292
transform 1 0 37904 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_412
timestamp 1621523292
transform 1 0 39008 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_424
timestamp 1621523292
transform 1 0 40112 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_436
timestamp 1621523292
transform 1 0 41216 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1621523292
transform 1 0 43056 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_448
timestamp 1621523292
transform 1 0 42320 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_457
timestamp 1621523292
transform 1 0 43148 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_469
timestamp 1621523292
transform 1 0 44252 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_481
timestamp 1621523292
transform 1 0 45356 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_493
timestamp 1621523292
transform 1 0 46460 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1621523292
transform 1 0 48300 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_505
timestamp 1621523292
transform 1 0 47564 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_514
timestamp 1621523292
transform 1 0 48392 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_526
timestamp 1621523292
transform 1 0 49496 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_538
timestamp 1621523292
transform 1 0 50600 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_550
timestamp 1621523292
transform 1 0 51704 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_562
timestamp 1621523292
transform 1 0 52808 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1621523292
transform 1 0 53544 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_571
timestamp 1621523292
transform 1 0 53636 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_583
timestamp 1621523292
transform 1 0 54740 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1588_
timestamp 1621523292
transform 1 0 57224 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2179_
timestamp 1621523292
transform 1 0 56580 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1621523292
transform 1 0 55568 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_95_591
timestamp 1621523292
transform 1 0 55476 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_595
timestamp 1621523292
transform 1 0 55844 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_606
timestamp 1621523292
transform 1 0 56856 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1621523292
transform -1 0 58880 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output204
timestamp 1621523292
transform 1 0 57868 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_613
timestamp 1621523292
transform 1 0 57500 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1621523292
transform 1 0 58236 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1621523292
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1621523292
transform 1 0 1380 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_6
timestamp 1621523292
transform 1 0 1656 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_18
timestamp 1621523292
transform 1 0 2760 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1621523292
transform 1 0 3772 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_26
timestamp 1621523292
transform 1 0 3496 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_30
timestamp 1621523292
transform 1 0 3864 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_42
timestamp 1621523292
transform 1 0 4968 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_54
timestamp 1621523292
transform 1 0 6072 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1621523292
transform 1 0 9016 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_66
timestamp 1621523292
transform 1 0 7176 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_78
timestamp 1621523292
transform 1 0 8280 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_87
timestamp 1621523292
transform 1 0 9108 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_99
timestamp 1621523292
transform 1 0 10212 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_111
timestamp 1621523292
transform 1 0 11316 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_123
timestamp 1621523292
transform 1 0 12420 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1621523292
transform 1 0 14260 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_135
timestamp 1621523292
transform 1 0 13524 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_144
timestamp 1621523292
transform 1 0 14352 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_156
timestamp 1621523292
transform 1 0 15456 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_168
timestamp 1621523292
transform 1 0 16560 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_180
timestamp 1621523292
transform 1 0 17664 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_192
timestamp 1621523292
transform 1 0 18768 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1621523292
transform 1 0 19504 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_201
timestamp 1621523292
transform 1 0 19596 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_213
timestamp 1621523292
transform 1 0 20700 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2351_
timestamp 1621523292
transform 1 0 21988 0 -1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_96_225
timestamp 1621523292
transform 1 0 21804 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _1817_
timestamp 1621523292
transform 1 0 23828 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1621523292
transform 1 0 24748 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_243
timestamp 1621523292
transform 1 0 23460 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_253
timestamp 1621523292
transform 1 0 24380 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_258
timestamp 1621523292
transform 1 0 24840 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _2355_
timestamp 1621523292
transform 1 0 26036 0 -1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_96_270
timestamp 1621523292
transform 1 0 25944 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1827_
timestamp 1621523292
transform 1 0 27876 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1891_
timestamp 1621523292
transform 1 0 28520 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_287
timestamp 1621523292
transform 1 0 27508 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_294
timestamp 1621523292
transform 1 0 28152 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_96_304
timestamp 1621523292
transform 1 0 29072 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _2484_
timestamp 1621523292
transform 1 0 30728 0 -1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1621523292
transform 1 0 29992 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_96_312
timestamp 1621523292
transform 1 0 29808 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_315
timestamp 1621523292
transform 1 0 30084 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_321
timestamp 1621523292
transform 1 0 30636 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1490_
timestamp 1621523292
transform 1 0 32568 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_96_338
timestamp 1621523292
transform 1 0 32200 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2186_
timestamp 1621523292
transform 1 0 33764 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1621523292
transform 1 0 35236 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_351
timestamp 1621523292
transform 1 0 33396 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_364
timestamp 1621523292
transform 1 0 34592 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_370
timestamp 1621523292
transform 1 0 35144 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _2097_
timestamp 1621523292
transform 1 0 36800 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1621523292
transform 1 0 35696 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_96_372
timestamp 1621523292
transform 1 0 35328 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_384
timestamp 1621523292
transform 1 0 36432 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_391
timestamp 1621523292
transform 1 0 37076 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_403
timestamp 1621523292
transform 1 0 38180 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1621523292
transform 1 0 40480 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_415
timestamp 1621523292
transform 1 0 39284 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_427
timestamp 1621523292
transform 1 0 40388 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_429
timestamp 1621523292
transform 1 0 40572 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_441
timestamp 1621523292
transform 1 0 41676 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_453
timestamp 1621523292
transform 1 0 42780 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_465
timestamp 1621523292
transform 1 0 43884 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_477
timestamp 1621523292
transform 1 0 44988 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1621523292
transform 1 0 45724 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_486
timestamp 1621523292
transform 1 0 45816 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_498
timestamp 1621523292
transform 1 0 46920 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_510
timestamp 1621523292
transform 1 0 48024 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_522
timestamp 1621523292
transform 1 0 49128 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1621523292
transform 1 0 50968 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_534
timestamp 1621523292
transform 1 0 50232 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_96_543
timestamp 1621523292
transform 1 0 51060 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_555
timestamp 1621523292
transform 1 0 52164 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_567
timestamp 1621523292
transform 1 0 53268 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1621523292
transform 1 0 54924 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1621523292
transform 1 0 54280 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_96_575
timestamp 1621523292
transform 1 0 54004 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_581
timestamp 1621523292
transform 1 0 54556 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_96_588
timestamp 1621523292
transform 1 0 55200 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2144_
timestamp 1621523292
transform 1 0 56856 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1621523292
transform 1 0 56212 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1621523292
transform 1 0 55568 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_595
timestamp 1621523292
transform 1 0 55844 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_96_600
timestamp 1621523292
transform 1 0 56304 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_96_609
timestamp 1621523292
transform 1 0 57132 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2293_
timestamp 1621523292
transform 1 0 57500 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1621523292
transform -1 0 58880 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_621
timestamp 1621523292
transform 1 0 58236 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1621523292
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1621523292
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1621523292
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1621523292
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1621523292
transform 1 0 4692 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1621523292
transform 1 0 6348 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_97_51
timestamp 1621523292
transform 1 0 5796 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_97_58
timestamp 1621523292
transform 1 0 6440 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_70
timestamp 1621523292
transform 1 0 7544 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_82
timestamp 1621523292
transform 1 0 8648 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_94
timestamp 1621523292
transform 1 0 9752 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_106
timestamp 1621523292
transform 1 0 10856 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1621523292
transform 1 0 11592 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_115
timestamp 1621523292
transform 1 0 11684 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_127
timestamp 1621523292
transform 1 0 12788 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_139
timestamp 1621523292
transform 1 0 13892 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_151
timestamp 1621523292
transform 1 0 14996 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1621523292
transform 1 0 16836 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_163
timestamp 1621523292
transform 1 0 16100 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_172
timestamp 1621523292
transform 1 0 16928 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_184
timestamp 1621523292
transform 1 0 18032 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_196
timestamp 1621523292
transform 1 0 19136 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_208
timestamp 1621523292
transform 1 0 20240 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1814_
timestamp 1621523292
transform 1 0 22540 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1621523292
transform 1 0 22080 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_220
timestamp 1621523292
transform 1 0 21344 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_97_229
timestamp 1621523292
transform 1 0 22172 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_97_239
timestamp 1621523292
transform 1 0 23092 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2352_
timestamp 1621523292
transform 1 0 23736 0 1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_97_245
timestamp 1621523292
transform 1 0 23644 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_262
timestamp 1621523292
transform 1 0 25208 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1824_
timestamp 1621523292
transform 1 0 26404 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1621523292
transform 1 0 25576 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_269
timestamp 1621523292
transform 1 0 25852 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_97_278
timestamp 1621523292
transform 1 0 26680 0 1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1825_
timestamp 1621523292
transform 1 0 27784 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2382_
timestamp 1621523292
transform 1 0 28980 0 1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1621523292
transform 1 0 27324 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_284
timestamp 1621523292
transform 1 0 27232 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_286
timestamp 1621523292
transform 1 0 27416 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_97_293
timestamp 1621523292
transform 1 0 28060 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_301
timestamp 1621523292
transform 1 0 28796 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_319
timestamp 1621523292
transform 1 0 30452 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_327
timestamp 1621523292
transform 1 0 31188 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__o221a_1  _1492_
timestamp 1621523292
transform 1 0 33120 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2188_
timestamp 1621523292
transform 1 0 31372 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1621523292
transform 1 0 32568 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_338
timestamp 1621523292
transform 1 0 32200 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_343
timestamp 1621523292
transform 1 0 32660 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_347
timestamp 1621523292
transform 1 0 33028 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _2342_
timestamp 1621523292
transform 1 0 34776 0 1 54944
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_97_357
timestamp 1621523292
transform 1 0 33948 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_97_365
timestamp 1621523292
transform 1 0 34684 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_382
timestamp 1621523292
transform 1 0 36248 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1621523292
transform 1 0 37812 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_394
timestamp 1621523292
transform 1 0 37352 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_398
timestamp 1621523292
transform 1 0 37720 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_400
timestamp 1621523292
transform 1 0 37904 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_412
timestamp 1621523292
transform 1 0 39008 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_424
timestamp 1621523292
transform 1 0 40112 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_436
timestamp 1621523292
transform 1 0 41216 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1621523292
transform 1 0 43056 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_448
timestamp 1621523292
transform 1 0 42320 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_457
timestamp 1621523292
transform 1 0 43148 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_469
timestamp 1621523292
transform 1 0 44252 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_481
timestamp 1621523292
transform 1 0 45356 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_493
timestamp 1621523292
transform 1 0 46460 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1621523292
transform 1 0 48300 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_505
timestamp 1621523292
transform 1 0 47564 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_514
timestamp 1621523292
transform 1 0 48392 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_526
timestamp 1621523292
transform 1 0 49496 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_538
timestamp 1621523292
transform 1 0 50600 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_550
timestamp 1621523292
transform 1 0 51704 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_562
timestamp 1621523292
transform 1 0 52808 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1621523292
transform 1 0 53544 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1621523292
transform 1 0 55200 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input156
timestamp 1621523292
transform 1 0 54556 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_571
timestamp 1621523292
transform 1 0 53636 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_579
timestamp 1621523292
transform 1 0 54372 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_584
timestamp 1621523292
transform 1 0 54832 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1544_
timestamp 1621523292
transform 1 0 56488 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2180_
timestamp 1621523292
transform 1 0 55844 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output243
timestamp 1621523292
transform 1 0 57132 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_591
timestamp 1621523292
transform 1 0 55476 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_598
timestamp 1621523292
transform 1 0 56120 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_605
timestamp 1621523292
transform 1 0 56764 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1621523292
transform -1 0 58880 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output205
timestamp 1621523292
transform 1 0 57868 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_613
timestamp 1621523292
transform 1 0 57500 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1621523292
transform 1 0 58236 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1621523292
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1621523292
transform 1 0 1380 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input175
timestamp 1621523292
transform 1 0 2024 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_6
timestamp 1621523292
transform 1 0 1656 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_13
timestamp 1621523292
transform 1 0 2300 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1621523292
transform 1 0 3772 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1621523292
transform 1 0 4232 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_25
timestamp 1621523292
transform 1 0 3404 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_30
timestamp 1621523292
transform 1 0 3864 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_37
timestamp 1621523292
transform 1 0 4508 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_49
timestamp 1621523292
transform 1 0 5612 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_61
timestamp 1621523292
transform 1 0 6716 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1244
timestamp 1621523292
transform 1 0 9016 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_73
timestamp 1621523292
transform 1 0 7820 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_85
timestamp 1621523292
transform 1 0 8924 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_87
timestamp 1621523292
transform 1 0 9108 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_99
timestamp 1621523292
transform 1 0 10212 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_111
timestamp 1621523292
transform 1 0 11316 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_123
timestamp 1621523292
transform 1 0 12420 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1245
timestamp 1621523292
transform 1 0 14260 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_135
timestamp 1621523292
transform 1 0 13524 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_144
timestamp 1621523292
transform 1 0 14352 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_156
timestamp 1621523292
transform 1 0 15456 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_168
timestamp 1621523292
transform 1 0 16560 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_180
timestamp 1621523292
transform 1 0 17664 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_192
timestamp 1621523292
transform 1 0 18768 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1246
timestamp 1621523292
transform 1 0 19504 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_201
timestamp 1621523292
transform 1 0 19596 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_213
timestamp 1621523292
transform 1 0 20700 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_225
timestamp 1621523292
transform 1 0 21804 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_237
timestamp 1621523292
transform 1 0 22908 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1818_
timestamp 1621523292
transform 1 0 25208 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1819_
timestamp 1621523292
transform 1 0 24104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1247
timestamp 1621523292
transform 1 0 24748 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_249
timestamp 1621523292
transform 1 0 24012 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_253
timestamp 1621523292
transform 1 0 24380 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_258
timestamp 1621523292
transform 1 0 24840 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1821_
timestamp 1621523292
transform 1 0 25852 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1826_
timestamp 1621523292
transform 1 0 26496 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_265
timestamp 1621523292
transform 1 0 25484 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_272
timestamp 1621523292
transform 1 0 26128 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_282
timestamp 1621523292
transform 1 0 27048 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1828_
timestamp 1621523292
transform 1 0 28796 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1829_
timestamp 1621523292
transform 1 0 27876 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_290
timestamp 1621523292
transform 1 0 27784 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_297
timestamp 1621523292
transform 1 0 28428 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_304
timestamp 1621523292
transform 1 0 29072 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1832_
timestamp 1621523292
transform 1 0 30452 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1248
timestamp 1621523292
transform 1 0 29992 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_98_312
timestamp 1621523292
transform 1 0 29808 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_315
timestamp 1621523292
transform 1 0 30084 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_325
timestamp 1621523292
transform 1 0 31004 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1831_
timestamp 1621523292
transform 1 0 31372 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2187_
timestamp 1621523292
transform 1 0 32200 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_98_332
timestamp 1621523292
transform 1 0 31648 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_347
timestamp 1621523292
transform 1 0 33028 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2482_
timestamp 1621523292
transform 1 0 33396 0 -1 56032
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1249
timestamp 1621523292
transform 1 0 35236 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_367
timestamp 1621523292
transform 1 0 34868 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1621523292
transform 1 0 35696 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_372
timestamp 1621523292
transform 1 0 35328 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_379
timestamp 1621523292
transform 1 0 35972 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_391
timestamp 1621523292
transform 1 0 37076 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_403
timestamp 1621523292
transform 1 0 38180 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1250
timestamp 1621523292
transform 1 0 40480 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_415
timestamp 1621523292
transform 1 0 39284 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_427
timestamp 1621523292
transform 1 0 40388 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_429
timestamp 1621523292
transform 1 0 40572 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_441
timestamp 1621523292
transform 1 0 41676 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_453
timestamp 1621523292
transform 1 0 42780 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_465
timestamp 1621523292
transform 1 0 43884 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_477
timestamp 1621523292
transform 1 0 44988 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1251
timestamp 1621523292
transform 1 0 45724 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_486
timestamp 1621523292
transform 1 0 45816 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_498
timestamp 1621523292
transform 1 0 46920 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_510
timestamp 1621523292
transform 1 0 48024 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_522
timestamp 1621523292
transform 1 0 49128 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1252
timestamp 1621523292
transform 1 0 50968 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_534
timestamp 1621523292
transform 1 0 50232 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_98_543
timestamp 1621523292
transform 1 0 51060 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input154
timestamp 1621523292
transform 1 0 53176 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1621523292
transform 1 0 52532 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_555
timestamp 1621523292
transform 1 0 52164 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_562
timestamp 1621523292
transform 1 0 52808 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _2183_
timestamp 1621523292
transform 1 0 54464 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input155
timestamp 1621523292
transform 1 0 53820 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_569
timestamp 1621523292
transform 1 0 53452 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_576
timestamp 1621523292
transform 1 0 54096 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_583
timestamp 1621523292
transform 1 0 54740 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1621523292
transform 1 0 56764 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _2181_
timestamp 1621523292
transform 1 0 55568 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1253
timestamp 1621523292
transform 1 0 56212 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_591
timestamp 1621523292
transform 1 0 55476 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_595
timestamp 1621523292
transform 1 0 55844 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_600
timestamp 1621523292
transform 1 0 56304 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_604
timestamp 1621523292
transform 1 0 56672 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_608
timestamp 1621523292
transform 1 0 57040 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2329_
timestamp 1621523292
transform 1 0 57500 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1621523292
transform -1 0 58880 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_98_612
timestamp 1621523292
transform 1 0 57408 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_621
timestamp 1621523292
transform 1 0 58236 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_6
timestamp 1621523292
transform 1 0 1656 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_6
timestamp 1621523292
transform 1 0 1656 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1621523292
transform 1 0 1380 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1621523292
transform 1 0 1380 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1621523292
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1621523292
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_14
timestamp 1621523292
transform 1 0 2392 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_10
timestamp 1621523292
transform 1 0 2024 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_13
timestamp 1621523292
transform 1 0 2300 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input138
timestamp 1621523292
transform 1 0 2668 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 1621523292
transform 1 0 2024 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1621523292
transform 1 0 2116 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_20
timestamp 1621523292
transform 1 0 2944 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_30
timestamp 1621523292
transform 1 0 3864 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_25
timestamp 1621523292
transform 1 0 3404 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1264
timestamp 1621523292
transform 1 0 3772 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1621523292
transform 1 0 3128 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_99_39
timestamp 1621523292
transform 1 0 4692 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_35
timestamp 1621523292
transform 1 0 4324 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 4232 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1621523292
transform 1 0 4784 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_42
timestamp 1621523292
transform 1 0 4968 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_43
timestamp 1621523292
transform 1 0 5060 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__or4b_4  _1359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 3312 0 1 56032
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1254
timestamp 1621523292
transform 1 0 6348 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_99_55
timestamp 1621523292
transform 1 0 6164 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_58
timestamp 1621523292
transform 1 0 6440 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_54
timestamp 1621523292
transform 1 0 6072 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1265
timestamp 1621523292
transform 1 0 9016 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input174
timestamp 1621523292
transform 1 0 8188 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_70
timestamp 1621523292
transform 1 0 7544 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_82
timestamp 1621523292
transform 1 0 8648 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_66
timestamp 1621523292
transform 1 0 7176 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_74
timestamp 1621523292
transform 1 0 7912 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_80
timestamp 1621523292
transform 1 0 8464 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_87
timestamp 1621523292
transform 1 0 9108 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1621523292
transform 1 0 10580 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_94
timestamp 1621523292
transform 1 0 9752 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_106
timestamp 1621523292
transform 1 0 10856 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1621523292
transform 1 0 10212 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_106
timestamp 1621523292
transform 1 0 10856 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _1361_
timestamp 1621523292
transform 1 0 11684 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _1469_
timestamp 1621523292
transform 1 0 12052 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1255
timestamp 1621523292
transform 1 0 11592 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input133
timestamp 1621523292
transform 1 0 12972 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_115
timestamp 1621523292
transform 1 0 11684 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_128
timestamp 1621523292
transform 1 0 12880 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_114
timestamp 1621523292
transform 1 0 11592 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_124
timestamp 1621523292
transform 1 0 12512 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_128
timestamp 1621523292
transform 1 0 12880 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1353_
timestamp 1621523292
transform 1 0 14720 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1266
timestamp 1621523292
transform 1 0 14260 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_140
timestamp 1621523292
transform 1 0 13984 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_152
timestamp 1621523292
transform 1 0 15088 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_133
timestamp 1621523292
transform 1 0 13340 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_141
timestamp 1621523292
transform 1 0 14076 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_144
timestamp 1621523292
transform 1 0 14352 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1256
timestamp 1621523292
transform 1 0 16836 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1621523292
transform 1 0 16100 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_99_164
timestamp 1621523292
transform 1 0 16192 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_170
timestamp 1621523292
transform 1 0 16744 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_172
timestamp 1621523292
transform 1 0 16928 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_157
timestamp 1621523292
transform 1 0 15548 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_166
timestamp 1621523292
transform 1 0 16376 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _1352_
timestamp 1621523292
transform 1 0 17572 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_99_184
timestamp 1621523292
transform 1 0 18032 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_196
timestamp 1621523292
transform 1 0 19136 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_178
timestamp 1621523292
transform 1 0 17480 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_188
timestamp 1621523292
transform 1 0 18400 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _1355_
timestamp 1621523292
transform 1 0 19964 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1356_
timestamp 1621523292
transform 1 0 21160 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1267
timestamp 1621523292
transform 1 0 19504 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_208
timestamp 1621523292
transform 1 0 20240 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_201
timestamp 1621523292
transform 1 0 19596 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_214
timestamp 1621523292
transform 1 0 20792 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_227
timestamp 1621523292
transform 1 0 21988 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_220
timestamp 1621523292
transform 1 0 21344 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1257
timestamp 1621523292
transform 1 0 22080 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_234
timestamp 1621523292
transform 1 0 22632 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_235
timestamp 1621523292
transform 1 0 22724 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_229
timestamp 1621523292
transform 1 0 22172 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1621523292
transform 1 0 22816 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1621523292
transform 1 0 22356 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1354_
timestamp 1621523292
transform 1 0 23000 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_99_239
timestamp 1621523292
transform 1 0 23092 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2353_
timestamp 1621523292
transform 1 0 23460 0 1 56032
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1268
timestamp 1621523292
transform 1 0 24748 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_259
timestamp 1621523292
transform 1 0 24932 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_247
timestamp 1621523292
transform 1 0 23828 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_255
timestamp 1621523292
transform 1 0 24564 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_100_258
timestamp 1621523292
transform 1 0 24840 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1350_
timestamp 1621523292
transform 1 0 26680 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1823_
timestamp 1621523292
transform 1 0 25576 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _2354_
timestamp 1621523292
transform 1 0 25300 0 1 56032
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_99_279
timestamp 1621523292
transform 1 0 26772 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_100_272
timestamp 1621523292
transform 1 0 26128 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _1349_
timestamp 1621523292
transform 1 0 28612 0 -1 57120
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1830_
timestamp 1621523292
transform 1 0 27968 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _2356_
timestamp 1621523292
transform 1 0 27784 0 1 56032
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1258
timestamp 1621523292
transform 1 0 27324 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_286
timestamp 1621523292
transform 1 0 27416 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_287
timestamp 1621523292
transform 1 0 27508 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_291
timestamp 1621523292
transform 1 0 27876 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_295
timestamp 1621523292
transform 1 0 28244 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _2357_
timestamp 1621523292
transform 1 0 29624 0 1 56032
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2358_
timestamp 1621523292
transform 1 0 31004 0 -1 57120
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1269
timestamp 1621523292
transform 1 0 29992 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_306
timestamp 1621523292
transform 1 0 29256 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_326
timestamp 1621523292
transform 1 0 31096 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_310
timestamp 1621523292
transform 1 0 29624 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_315
timestamp 1621523292
transform 1 0 30084 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_323
timestamp 1621523292
transform 1 0 30820 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1351_
timestamp 1621523292
transform 1 0 33028 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1834_
timestamp 1621523292
transform 1 0 31464 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1259
timestamp 1621523292
transform 1 0 32568 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_338
timestamp 1621523292
transform 1 0 32200 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_343
timestamp 1621523292
transform 1 0 32660 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_341
timestamp 1621523292
transform 1 0 32476 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_349
timestamp 1621523292
transform 1 0 33212 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__o221a_1  _1491_
timestamp 1621523292
transform 1 0 34224 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _2483_
timestamp 1621523292
transform 1 0 33304 0 -1 57120
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1270
timestamp 1621523292
transform 1 0 35236 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_356
timestamp 1621523292
transform 1 0 33856 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_369
timestamp 1621523292
transform 1 0 35052 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_366
timestamp 1621523292
transform 1 0 34776 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_370
timestamp 1621523292
transform 1 0 35144 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_379
timestamp 1621523292
transform 1 0 35972 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_372
timestamp 1621523292
transform 1 0 35328 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_376
timestamp 1621523292
transform 1 0 35696 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1621523292
transform 1 0 36064 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1621523292
transform 1 0 35420 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1621523292
transform 1 0 35696 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_393
timestamp 1621523292
transform 1 0 37260 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_386
timestamp 1621523292
transform 1 0 36616 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1621523292
transform 1 0 36984 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1621523292
transform 1 0 36340 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_383
timestamp 1621523292
transform 1 0 36340 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1260
timestamp 1621523292
transform 1 0 37812 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1621523292
transform 1 0 37628 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_395
timestamp 1621523292
transform 1 0 37444 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_400
timestamp 1621523292
transform 1 0 37904 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_412
timestamp 1621523292
transform 1 0 39008 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_400
timestamp 1621523292
transform 1 0 37904 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_412
timestamp 1621523292
transform 1 0 39008 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1271
timestamp 1621523292
transform 1 0 40480 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1621523292
transform 1 0 39744 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_424
timestamp 1621523292
transform 1 0 40112 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_436
timestamp 1621523292
transform 1 0 41216 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_423
timestamp 1621523292
transform 1 0 40020 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_427
timestamp 1621523292
transform 1 0 40388 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_429
timestamp 1621523292
transform 1 0 40572 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1261
timestamp 1621523292
transform 1 0 43056 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input170
timestamp 1621523292
transform 1 0 42136 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_448
timestamp 1621523292
transform 1 0 42320 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_457
timestamp 1621523292
transform 1 0 43148 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_441
timestamp 1621523292
transform 1 0 41676 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_445
timestamp 1621523292
transform 1 0 42044 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_449
timestamp 1621523292
transform 1 0 42412 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_469
timestamp 1621523292
transform 1 0 44252 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_461
timestamp 1621523292
transform 1 0 43516 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_473
timestamp 1621523292
transform 1 0 44620 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1272
timestamp 1621523292
transform 1 0 45724 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_481
timestamp 1621523292
transform 1 0 45356 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_493
timestamp 1621523292
transform 1 0 46460 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_486
timestamp 1621523292
transform 1 0 45816 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_498
timestamp 1621523292
transform 1 0 46920 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1262
timestamp 1621523292
transform 1 0 48300 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_505
timestamp 1621523292
transform 1 0 47564 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_514
timestamp 1621523292
transform 1 0 48392 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_510
timestamp 1621523292
transform 1 0 48024 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_522
timestamp 1621523292
transform 1 0 49128 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1273
timestamp 1621523292
transform 1 0 50968 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_526
timestamp 1621523292
transform 1 0 49496 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_538
timestamp 1621523292
transform 1 0 50600 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_534
timestamp 1621523292
transform 1 0 50232 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_100_543
timestamp 1621523292
transform 1 0 51060 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_550
timestamp 1621523292
transform 1 0 51704 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_554
timestamp 1621523292
transform 1 0 52072 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_550
timestamp 1621523292
transform 1 0 51704 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1621523292
transform 1 0 51796 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1621523292
transform 1 0 52072 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1621523292
transform 1 0 51428 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_557
timestamp 1621523292
transform 1 0 52348 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_99_561
timestamp 1621523292
transform 1 0 52716 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input153
timestamp 1621523292
transform 1 0 52440 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_565
timestamp 1621523292
transform 1 0 53084 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _2185_
timestamp 1621523292
transform 1 0 53268 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_570
timestamp 1621523292
transform 1 0 53544 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_571
timestamp 1621523292
transform 1 0 53636 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_569
timestamp 1621523292
transform 1 0 53452 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1263
timestamp 1621523292
transform 1 0 53544 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _2182_
timestamp 1621523292
transform 1 0 53912 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_577
timestamp 1621523292
transform 1 0 54188 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_580
timestamp 1621523292
transform 1 0 54464 0 1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  _2332_
timestamp 1621523292
transform 1 0 54556 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1711_
timestamp 1621523292
transform 1 0 54188 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_100_589
timestamp 1621523292
transform 1 0 55292 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_586
timestamp 1621523292
transform 1 0 55016 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _1543_
timestamp 1621523292
transform 1 0 55108 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _2334_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 55752 0 1 56032
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1274
timestamp 1621523292
transform 1 0 56212 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output244
timestamp 1621523292
transform 1 0 56764 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_590
timestamp 1621523292
transform 1 0 55384 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_100_597
timestamp 1621523292
transform 1 0 56028 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_600
timestamp 1621523292
transform 1 0 56304 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_604
timestamp 1621523292
transform 1 0 56672 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_609
timestamp 1621523292
transform 1 0 57132 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_1  _2330_
timestamp 1621523292
transform 1 0 57500 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1621523292
transform -1 0 58880 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1621523292
transform -1 0 58880 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_615
timestamp 1621523292
transform 1 0 57684 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1621523292
transform 1 0 58420 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1621523292
transform 1 0 58236 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1621523292
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output255
timestamp 1621523292
transform 1 0 1748 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output288
timestamp 1621523292
transform 1 0 3036 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_3
timestamp 1621523292
transform 1 0 1380 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_11
timestamp 1621523292
transform 1 0 2116 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_19
timestamp 1621523292
transform 1 0 2852 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__ebufn_1  _2191_
timestamp 1621523292
transform 1 0 4232 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1275
timestamp 1621523292
transform 1 0 3772 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_25
timestamp 1621523292
transform 1 0 3404 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_30
timestamp 1621523292
transform 1 0 3864 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_42
timestamp 1621523292
transform 1 0 4968 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1276
timestamp 1621523292
transform 1 0 6440 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1621523292
transform 1 0 5336 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1621523292
transform 1 0 6900 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_50
timestamp 1621523292
transform 1 0 5704 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_59
timestamp 1621523292
transform 1 0 6532 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1277
timestamp 1621523292
transform 1 0 9108 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1621523292
transform 1 0 7544 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input173
timestamp 1621523292
transform 1 0 8188 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_66
timestamp 1621523292
transform 1 0 7176 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_73
timestamp 1621523292
transform 1 0 7820 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_80
timestamp 1621523292
transform 1 0 8464 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_86
timestamp 1621523292
transform 1 0 9016 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1621523292
transform 1 0 9568 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1621523292
transform 1 0 10212 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input131
timestamp 1621523292
transform 1 0 11040 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_88
timestamp 1621523292
transform 1 0 9200 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_95
timestamp 1621523292
transform 1 0 9844 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_102
timestamp 1621523292
transform 1 0 10488 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _1366_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1621523292
transform 1 0 12236 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1278
timestamp 1621523292
transform 1 0 11776 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_112
timestamp 1621523292
transform 1 0 11408 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_117
timestamp 1621523292
transform 1 0 11868 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_130
timestamp 1621523292
transform 1 0 13064 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1279
timestamp 1621523292
transform 1 0 14444 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  input132
timestamp 1621523292
transform 1 0 13432 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1621523292
transform 1 0 14904 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_138
timestamp 1621523292
transform 1 0 13800 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_144
timestamp 1621523292
transform 1 0 14352 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_146
timestamp 1621523292
transform 1 0 14536 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1280
timestamp 1621523292
transform 1 0 17112 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1621523292
transform 1 0 15548 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1621523292
transform 1 0 16192 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_153
timestamp 1621523292
transform 1 0 15180 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_160
timestamp 1621523292
transform 1 0 15824 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_167
timestamp 1621523292
transform 1 0 16468 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_173
timestamp 1621523292
transform 1 0 17020 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1621523292
transform 1 0 17572 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1621523292
transform 1 0 18216 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1621523292
transform 1 0 18860 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_175
timestamp 1621523292
transform 1 0 17204 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_182
timestamp 1621523292
transform 1 0 17848 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_189
timestamp 1621523292
transform 1 0 18492 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_196
timestamp 1621523292
transform 1 0 19136 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1281
timestamp 1621523292
transform 1 0 19780 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1621523292
transform 1 0 20240 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1621523292
transform 1 0 20884 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_202
timestamp 1621523292
transform 1 0 19688 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_204
timestamp 1621523292
transform 1 0 19872 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_211
timestamp 1621523292
transform 1 0 20516 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_218
timestamp 1621523292
transform 1 0 21160 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1282
timestamp 1621523292
transform 1 0 22448 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1621523292
transform 1 0 21528 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1621523292
transform 1 0 22908 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_225
timestamp 1621523292
transform 1 0 21804 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_231
timestamp 1621523292
transform 1 0 22356 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_233
timestamp 1621523292
transform 1 0 22540 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_240
timestamp 1621523292
transform 1 0 23184 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1820_
timestamp 1621523292
transform 1 0 24104 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1283
timestamp 1621523292
transform 1 0 25116 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_248
timestamp 1621523292
transform 1 0 23920 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_256
timestamp 1621523292
transform 1 0 24656 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_260
timestamp 1621523292
transform 1 0 25024 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_262
timestamp 1621523292
transform 1 0 25208 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _1357_
timestamp 1621523292
transform 1 0 26588 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1822_
timestamp 1621523292
transform 1 0 25944 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_273
timestamp 1621523292
transform 1 0 26220 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1621523292
transform 1 0 29072 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1284
timestamp 1621523292
transform 1 0 27784 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1621523292
transform 1 0 28244 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_286
timestamp 1621523292
transform 1 0 27416 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_291
timestamp 1621523292
transform 1 0 27876 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_298
timestamp 1621523292
transform 1 0 28520 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1285
timestamp 1621523292
transform 1 0 30452 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1621523292
transform 1 0 29716 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_307
timestamp 1621523292
transform 1 0 29348 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_314
timestamp 1621523292
transform 1 0 29992 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_318
timestamp 1621523292
transform 1 0 30360 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_320
timestamp 1621523292
transform 1 0 30544 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1833_
timestamp 1621523292
transform 1 0 31464 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1286
timestamp 1621523292
transform 1 0 33120 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1621523292
transform 1 0 32108 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_328
timestamp 1621523292
transform 1 0 31280 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_333
timestamp 1621523292
transform 1 0 31740 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_340
timestamp 1621523292
transform 1 0 32384 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_349
timestamp 1621523292
transform 1 0 33212 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1621523292
transform 1 0 33580 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1621523292
transform 1 0 34224 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input139
timestamp 1621523292
transform 1 0 35052 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_356
timestamp 1621523292
transform 1 0 33856 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_363
timestamp 1621523292
transform 1 0 34500 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1287
timestamp 1621523292
transform 1 0 35788 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1621523292
transform 1 0 36248 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1621523292
transform 1 0 36892 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_373
timestamp 1621523292
transform 1 0 35420 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_378
timestamp 1621523292
transform 1 0 35880 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_385
timestamp 1621523292
transform 1 0 36524 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_392
timestamp 1621523292
transform 1 0 37168 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1288
timestamp 1621523292
transform 1 0 38456 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1621523292
transform 1 0 37536 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1621523292
transform 1 0 38916 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_399
timestamp 1621523292
transform 1 0 37812 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_405
timestamp 1621523292
transform 1 0 38364 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_407
timestamp 1621523292
transform 1 0 38548 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_414
timestamp 1621523292
transform 1 0 39192 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1289
timestamp 1621523292
transform 1 0 41124 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1621523292
transform 1 0 39560 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1621523292
transform 1 0 40204 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_421
timestamp 1621523292
transform 1 0 39836 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_428
timestamp 1621523292
transform 1 0 40480 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_434
timestamp 1621523292
transform 1 0 41032 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_436
timestamp 1621523292
transform 1 0 41216 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input140
timestamp 1621523292
transform 1 0 42964 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1621523292
transform 1 0 41584 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1621523292
transform 1 0 42228 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_443
timestamp 1621523292
transform 1 0 41860 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_450
timestamp 1621523292
transform 1 0 42504 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_454
timestamp 1621523292
transform 1 0 42872 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_458
timestamp 1621523292
transform 1 0 43240 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1290
timestamp 1621523292
transform 1 0 43792 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1621523292
transform 1 0 44252 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1621523292
transform 1 0 44896 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_465
timestamp 1621523292
transform 1 0 43884 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_472
timestamp 1621523292
transform 1 0 44528 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_479
timestamp 1621523292
transform 1 0 45172 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1291
timestamp 1621523292
transform 1 0 46460 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1621523292
transform 1 0 45540 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1621523292
transform 1 0 46920 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_486
timestamp 1621523292
transform 1 0 45816 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_492
timestamp 1621523292
transform 1 0 46368 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_494
timestamp 1621523292
transform 1 0 46552 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_501
timestamp 1621523292
transform 1 0 47196 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1292
timestamp 1621523292
transform 1 0 49128 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1621523292
transform 1 0 47564 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input146
timestamp 1621523292
transform 1 0 48208 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_508
timestamp 1621523292
transform 1 0 47840 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_515
timestamp 1621523292
transform 1 0 48484 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_521
timestamp 1621523292
transform 1 0 49036 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_523
timestamp 1621523292
transform 1 0 49220 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1621523292
transform 1 0 49588 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1621523292
transform 1 0 50232 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1621523292
transform 1 0 50876 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_530
timestamp 1621523292
transform 1 0 49864 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_537
timestamp 1621523292
transform 1 0 50508 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_544
timestamp 1621523292
transform 1 0 51152 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1293
timestamp 1621523292
transform 1 0 51796 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1621523292
transform 1 0 52348 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output253
timestamp 1621523292
transform 1 0 52992 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_550
timestamp 1621523292
transform 1 0 51704 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_552
timestamp 1621523292
transform 1 0 51888 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_556
timestamp 1621523292
transform 1 0 52256 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_560
timestamp 1621523292
transform 1 0 52624 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1294
timestamp 1621523292
transform 1 0 54464 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output207
timestamp 1621523292
transform 1 0 55292 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output245
timestamp 1621523292
transform 1 0 53728 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_568
timestamp 1621523292
transform 1 0 53360 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_576
timestamp 1621523292
transform 1 0 54096 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_581
timestamp 1621523292
transform 1 0 54556 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__ebufn_1  _2331_
timestamp 1621523292
transform 1 0 56028 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1295
timestamp 1621523292
transform 1 0 57132 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_593
timestamp 1621523292
transform 1 0 55660 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_605
timestamp 1621523292
transform 1 0 56764 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_610
timestamp 1621523292
transform 1 0 57224 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1621523292
transform -1 0 58880 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output206
timestamp 1621523292
transform 1 0 57868 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_616
timestamp 1621523292
transform 1 0 57776 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1621523292
transform 1 0 58236 0 1 57120
box -38 -48 406 592
<< labels >>
rlabel metal2 s 5078 59200 5134 60000 6 active
port 0 nsew signal input
rlabel metal3 s 59200 144 60000 264 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 59200 15784 60000 15904 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 59200 17280 60000 17400 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 59200 18912 60000 19032 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 59200 22040 60000 22160 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 59200 23536 60000 23656 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 59200 25168 60000 25288 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 59200 26664 60000 26784 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 59200 28296 60000 28416 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 59200 29792 60000 29912 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 59200 1640 60000 1760 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 59200 31424 60000 31544 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 59200 32920 60000 33040 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 59200 34552 60000 34672 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 59200 36048 60000 36168 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 59200 37680 60000 37800 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 59200 39176 60000 39296 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 59200 40808 60000 40928 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 59200 42304 60000 42424 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 59200 43936 60000 44056 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 59200 45432 60000 45552 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 59200 3272 60000 3392 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 59200 47064 60000 47184 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 59200 48560 60000 48680 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 59200 50192 60000 50312 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 59200 51688 60000 51808 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 59200 53320 60000 53440 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 59200 54816 60000 54936 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 59200 56448 60000 56568 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59200 57944 60000 58064 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 59200 4768 60000 4888 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 59200 6400 60000 6520 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 59200 7896 60000 8016 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 59200 9528 60000 9648 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 59200 11024 60000 11144 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 59200 12656 60000 12776 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 59200 14152 60000 14272 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 59200 1096 60000 1216 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 59200 16736 60000 16856 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 59200 18368 60000 18488 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 59200 19864 60000 19984 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 59200 21496 60000 21616 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 59200 22992 60000 23112 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal3 s 59200 24624 60000 24744 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 59200 26120 60000 26240 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal3 s 59200 27752 60000 27872 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal3 s 59200 29248 60000 29368 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal3 s 59200 30880 60000 31000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal3 s 59200 2728 60000 2848 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 59200 32376 60000 32496 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 59200 34008 60000 34128 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal3 s 59200 35504 60000 35624 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal3 s 59200 37136 60000 37256 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal3 s 59200 38632 60000 38752 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 59200 40264 60000 40384 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 59200 41760 60000 41880 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal3 s 59200 43392 60000 43512 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal3 s 59200 44888 60000 45008 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 59200 46520 60000 46640 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal3 s 59200 4224 60000 4344 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 59200 48016 60000 48136 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 59200 49648 60000 49768 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 59200 51144 60000 51264 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 59200 52776 60000 52896 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 59200 54272 60000 54392 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 59200 55904 60000 56024 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 59200 57400 60000 57520 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 59200 59032 60000 59152 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal3 s 59200 5856 60000 5976 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 59200 7352 60000 7472 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 59200 8984 60000 9104 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 59200 10480 60000 10600 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal3 s 59200 12112 60000 12232 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal3 s 59200 13608 60000 13728 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal3 s 59200 15240 60000 15360 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 59200 552 60000 672 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 59200 16192 60000 16312 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 59200 17824 60000 17944 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 59200 19320 60000 19440 6 io_out[12]
port 80 nsew signal tristate
rlabel metal3 s 59200 20952 60000 21072 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 59200 22448 60000 22568 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 59200 24080 60000 24200 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 59200 25576 60000 25696 6 io_out[16]
port 84 nsew signal tristate
rlabel metal3 s 59200 27208 60000 27328 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 59200 28704 60000 28824 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 59200 30336 60000 30456 6 io_out[19]
port 87 nsew signal tristate
rlabel metal3 s 59200 2184 60000 2304 6 io_out[1]
port 88 nsew signal tristate
rlabel metal3 s 59200 31832 60000 31952 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 59200 33464 60000 33584 6 io_out[21]
port 90 nsew signal tristate
rlabel metal3 s 59200 34960 60000 35080 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 59200 36592 60000 36712 6 io_out[23]
port 92 nsew signal tristate
rlabel metal3 s 59200 38088 60000 38208 6 io_out[24]
port 93 nsew signal tristate
rlabel metal3 s 59200 39720 60000 39840 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 59200 41216 60000 41336 6 io_out[26]
port 95 nsew signal tristate
rlabel metal3 s 59200 42848 60000 42968 6 io_out[27]
port 96 nsew signal tristate
rlabel metal3 s 59200 44344 60000 44464 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 59200 45976 60000 46096 6 io_out[29]
port 98 nsew signal tristate
rlabel metal3 s 59200 3680 60000 3800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 59200 47472 60000 47592 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 59200 49104 60000 49224 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 59200 50600 60000 50720 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 59200 52232 60000 52352 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 59200 53728 60000 53848 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 59200 55360 60000 55480 6 io_out[35]
port 105 nsew signal tristate
rlabel metal3 s 59200 56856 60000 56976 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 59200 58488 60000 58608 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 59200 5312 60000 5432 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 59200 6808 60000 6928 6 io_out[4]
port 109 nsew signal tristate
rlabel metal3 s 59200 8440 60000 8560 6 io_out[5]
port 110 nsew signal tristate
rlabel metal3 s 59200 9936 60000 10056 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 59200 11568 60000 11688 6 io_out[7]
port 112 nsew signal tristate
rlabel metal3 s 59200 13064 60000 13184 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 59200 14696 60000 14816 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 59200 59576 60000 59696 6 irq[0]
port 115 nsew signal tristate
rlabel metal2 s 59450 0 59506 800 6 irq[1]
port 116 nsew signal tristate
rlabel metal3 s 0 59440 800 59560 6 irq[2]
port 117 nsew signal tristate
rlabel metal2 s 478 0 534 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 la_data_in[11]
port 120 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_data_in[12]
port 121 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 la_data_in[13]
port 122 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 la_data_in[14]
port 123 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_data_in[16]
port 125 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_data_in[17]
port 126 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_data_in[18]
port 127 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_data_in[20]
port 130 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[22]
port 132 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[24]
port 134 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[26]
port 136 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[27]
port 137 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[28]
port 138 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[29]
port 139 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_data_in[30]
port 141 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 la_data_in[3]
port 143 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la_data_in[4]
port 144 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 la_data_in[5]
port 145 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 la_data_in[6]
port 146 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 la_data_in[7]
port 147 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 la_data_in[8]
port 148 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 la_data_in[9]
port 149 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_out[0]
port 150 nsew signal tristate
rlabel metal2 s 39210 0 39266 800 6 la_data_out[10]
port 151 nsew signal tristate
rlabel metal2 s 40130 0 40186 800 6 la_data_out[11]
port 152 nsew signal tristate
rlabel metal2 s 41050 0 41106 800 6 la_data_out[12]
port 153 nsew signal tristate
rlabel metal2 s 41970 0 42026 800 6 la_data_out[13]
port 154 nsew signal tristate
rlabel metal2 s 42890 0 42946 800 6 la_data_out[14]
port 155 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 la_data_out[15]
port 156 nsew signal tristate
rlabel metal2 s 44730 0 44786 800 6 la_data_out[16]
port 157 nsew signal tristate
rlabel metal2 s 45650 0 45706 800 6 la_data_out[17]
port 158 nsew signal tristate
rlabel metal2 s 46570 0 46626 800 6 la_data_out[18]
port 159 nsew signal tristate
rlabel metal2 s 47490 0 47546 800 6 la_data_out[19]
port 160 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 la_data_out[1]
port 161 nsew signal tristate
rlabel metal2 s 48410 0 48466 800 6 la_data_out[20]
port 162 nsew signal tristate
rlabel metal2 s 49330 0 49386 800 6 la_data_out[21]
port 163 nsew signal tristate
rlabel metal2 s 50250 0 50306 800 6 la_data_out[22]
port 164 nsew signal tristate
rlabel metal2 s 51170 0 51226 800 6 la_data_out[23]
port 165 nsew signal tristate
rlabel metal2 s 52090 0 52146 800 6 la_data_out[24]
port 166 nsew signal tristate
rlabel metal2 s 53010 0 53066 800 6 la_data_out[25]
port 167 nsew signal tristate
rlabel metal2 s 53930 0 53986 800 6 la_data_out[26]
port 168 nsew signal tristate
rlabel metal2 s 54850 0 54906 800 6 la_data_out[27]
port 169 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 la_data_out[28]
port 170 nsew signal tristate
rlabel metal2 s 56690 0 56746 800 6 la_data_out[29]
port 171 nsew signal tristate
rlabel metal2 s 31850 0 31906 800 6 la_data_out[2]
port 172 nsew signal tristate
rlabel metal2 s 57610 0 57666 800 6 la_data_out[30]
port 173 nsew signal tristate
rlabel metal2 s 58530 0 58586 800 6 la_data_out[31]
port 174 nsew signal tristate
rlabel metal2 s 32770 0 32826 800 6 la_data_out[3]
port 175 nsew signal tristate
rlabel metal2 s 33690 0 33746 800 6 la_data_out[4]
port 176 nsew signal tristate
rlabel metal2 s 34610 0 34666 800 6 la_data_out[5]
port 177 nsew signal tristate
rlabel metal2 s 35530 0 35586 800 6 la_data_out[6]
port 178 nsew signal tristate
rlabel metal2 s 36450 0 36506 800 6 la_data_out[7]
port 179 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 la_data_out[8]
port 180 nsew signal tristate
rlabel metal2 s 38290 0 38346 800 6 la_data_out[9]
port 181 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 la_oenb[0]
port 182 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 la_oenb[10]
port 183 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 la_oenb[11]
port 184 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 la_oenb[12]
port 185 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 la_oenb[13]
port 186 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[14]
port 187 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 la_oenb[15]
port 188 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 la_oenb[16]
port 189 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[17]
port 190 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la_oenb[18]
port 191 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 la_oenb[19]
port 192 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 la_oenb[1]
port 193 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_oenb[20]
port 194 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 la_oenb[21]
port 195 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 la_oenb[22]
port 196 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 la_oenb[23]
port 197 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 la_oenb[24]
port 198 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 la_oenb[25]
port 199 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 la_oenb[26]
port 200 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 la_oenb[27]
port 201 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 la_oenb[28]
port 202 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la_oenb[29]
port 203 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 la_oenb[2]
port 204 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 la_oenb[30]
port 205 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 la_oenb[31]
port 206 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_oenb[3]
port 207 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 la_oenb[4]
port 208 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 la_oenb[5]
port 209 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_oenb[6]
port 210 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la_oenb[7]
port 211 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 la_oenb[8]
port 212 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 la_oenb[9]
port 213 nsew signal input
rlabel metal2 s 386 59200 442 60000 6 wb_clk_i
port 214 nsew signal input
rlabel metal2 s 1122 59200 1178 60000 6 wb_rst_i
port 215 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 wbs_ack_o
port 216 nsew signal tristate
rlabel metal2 s 9034 59200 9090 60000 6 wbs_adr_i[0]
port 217 nsew signal input
rlabel metal2 s 16946 59200 17002 60000 6 wbs_adr_i[10]
port 218 nsew signal input
rlabel metal2 s 17682 59200 17738 60000 6 wbs_adr_i[11]
port 219 nsew signal input
rlabel metal2 s 18510 59200 18566 60000 6 wbs_adr_i[12]
port 220 nsew signal input
rlabel metal2 s 19246 59200 19302 60000 6 wbs_adr_i[13]
port 221 nsew signal input
rlabel metal2 s 20074 59200 20130 60000 6 wbs_adr_i[14]
port 222 nsew signal input
rlabel metal2 s 20902 59200 20958 60000 6 wbs_adr_i[15]
port 223 nsew signal input
rlabel metal2 s 21638 59200 21694 60000 6 wbs_adr_i[16]
port 224 nsew signal input
rlabel metal2 s 22466 59200 22522 60000 6 wbs_adr_i[17]
port 225 nsew signal input
rlabel metal2 s 23202 59200 23258 60000 6 wbs_adr_i[18]
port 226 nsew signal input
rlabel metal2 s 24030 59200 24086 60000 6 wbs_adr_i[19]
port 227 nsew signal input
rlabel metal2 s 9770 59200 9826 60000 6 wbs_adr_i[1]
port 228 nsew signal input
rlabel metal2 s 24766 59200 24822 60000 6 wbs_adr_i[20]
port 229 nsew signal input
rlabel metal2 s 25594 59200 25650 60000 6 wbs_adr_i[21]
port 230 nsew signal input
rlabel metal2 s 26422 59200 26478 60000 6 wbs_adr_i[22]
port 231 nsew signal input
rlabel metal2 s 27158 59200 27214 60000 6 wbs_adr_i[23]
port 232 nsew signal input
rlabel metal2 s 27986 59200 28042 60000 6 wbs_adr_i[24]
port 233 nsew signal input
rlabel metal2 s 28722 59200 28778 60000 6 wbs_adr_i[25]
port 234 nsew signal input
rlabel metal2 s 29550 59200 29606 60000 6 wbs_adr_i[26]
port 235 nsew signal input
rlabel metal2 s 30378 59200 30434 60000 6 wbs_adr_i[27]
port 236 nsew signal input
rlabel metal2 s 31114 59200 31170 60000 6 wbs_adr_i[28]
port 237 nsew signal input
rlabel metal2 s 31942 59200 31998 60000 6 wbs_adr_i[29]
port 238 nsew signal input
rlabel metal2 s 10598 59200 10654 60000 6 wbs_adr_i[2]
port 239 nsew signal input
rlabel metal2 s 32678 59200 32734 60000 6 wbs_adr_i[30]
port 240 nsew signal input
rlabel metal2 s 33506 59200 33562 60000 6 wbs_adr_i[31]
port 241 nsew signal input
rlabel metal2 s 34242 59200 34298 60000 6 wbs_adr_i[32]
port 242 nsew signal input
rlabel metal2 s 11426 59200 11482 60000 6 wbs_adr_i[3]
port 243 nsew signal input
rlabel metal2 s 12162 59200 12218 60000 6 wbs_adr_i[4]
port 244 nsew signal input
rlabel metal2 s 12990 59200 13046 60000 6 wbs_adr_i[5]
port 245 nsew signal input
rlabel metal2 s 13726 59200 13782 60000 6 wbs_adr_i[6]
port 246 nsew signal input
rlabel metal2 s 14554 59200 14610 60000 6 wbs_adr_i[7]
port 247 nsew signal input
rlabel metal2 s 15382 59200 15438 60000 6 wbs_adr_i[8]
port 248 nsew signal input
rlabel metal2 s 16118 59200 16174 60000 6 wbs_adr_i[9]
port 249 nsew signal input
rlabel metal2 s 2686 59200 2742 60000 6 wbs_cyc_i
port 250 nsew signal input
rlabel metal2 s 35070 59200 35126 60000 6 wbs_dat_i[0]
port 251 nsew signal input
rlabel metal2 s 42982 59200 43038 60000 6 wbs_dat_i[10]
port 252 nsew signal input
rlabel metal2 s 43718 59200 43774 60000 6 wbs_dat_i[11]
port 253 nsew signal input
rlabel metal2 s 44546 59200 44602 60000 6 wbs_dat_i[12]
port 254 nsew signal input
rlabel metal2 s 45374 59200 45430 60000 6 wbs_dat_i[13]
port 255 nsew signal input
rlabel metal2 s 46110 59200 46166 60000 6 wbs_dat_i[14]
port 256 nsew signal input
rlabel metal2 s 46938 59200 46994 60000 6 wbs_dat_i[15]
port 257 nsew signal input
rlabel metal2 s 47674 59200 47730 60000 6 wbs_dat_i[16]
port 258 nsew signal input
rlabel metal2 s 48502 59200 48558 60000 6 wbs_dat_i[17]
port 259 nsew signal input
rlabel metal2 s 49238 59200 49294 60000 6 wbs_dat_i[18]
port 260 nsew signal input
rlabel metal2 s 50066 59200 50122 60000 6 wbs_dat_i[19]
port 261 nsew signal input
rlabel metal2 s 35898 59200 35954 60000 6 wbs_dat_i[1]
port 262 nsew signal input
rlabel metal2 s 50894 59200 50950 60000 6 wbs_dat_i[20]
port 263 nsew signal input
rlabel metal2 s 51630 59200 51686 60000 6 wbs_dat_i[21]
port 264 nsew signal input
rlabel metal2 s 52458 59200 52514 60000 6 wbs_dat_i[22]
port 265 nsew signal input
rlabel metal2 s 53194 59200 53250 60000 6 wbs_dat_i[23]
port 266 nsew signal input
rlabel metal2 s 54022 59200 54078 60000 6 wbs_dat_i[24]
port 267 nsew signal input
rlabel metal2 s 54758 59200 54814 60000 6 wbs_dat_i[25]
port 268 nsew signal input
rlabel metal2 s 55586 59200 55642 60000 6 wbs_dat_i[26]
port 269 nsew signal input
rlabel metal2 s 56414 59200 56470 60000 6 wbs_dat_i[27]
port 270 nsew signal input
rlabel metal2 s 57150 59200 57206 60000 6 wbs_dat_i[28]
port 271 nsew signal input
rlabel metal2 s 57978 59200 58034 60000 6 wbs_dat_i[29]
port 272 nsew signal input
rlabel metal2 s 36634 59200 36690 60000 6 wbs_dat_i[2]
port 273 nsew signal input
rlabel metal2 s 58714 59200 58770 60000 6 wbs_dat_i[30]
port 274 nsew signal input
rlabel metal2 s 59542 59200 59598 60000 6 wbs_dat_i[31]
port 275 nsew signal input
rlabel metal2 s 37462 59200 37518 60000 6 wbs_dat_i[3]
port 276 nsew signal input
rlabel metal2 s 38198 59200 38254 60000 6 wbs_dat_i[4]
port 277 nsew signal input
rlabel metal2 s 39026 59200 39082 60000 6 wbs_dat_i[5]
port 278 nsew signal input
rlabel metal2 s 39762 59200 39818 60000 6 wbs_dat_i[6]
port 279 nsew signal input
rlabel metal2 s 40590 59200 40646 60000 6 wbs_dat_i[7]
port 280 nsew signal input
rlabel metal2 s 41418 59200 41474 60000 6 wbs_dat_i[8]
port 281 nsew signal input
rlabel metal2 s 42154 59200 42210 60000 6 wbs_dat_i[9]
port 282 nsew signal input
rlabel metal3 s 0 416 800 536 6 wbs_dat_o[0]
port 283 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 wbs_dat_o[10]
port 284 nsew signal tristate
rlabel metal3 s 0 10480 800 10600 6 wbs_dat_o[11]
port 285 nsew signal tristate
rlabel metal3 s 0 11432 800 11552 6 wbs_dat_o[12]
port 286 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 wbs_dat_o[13]
port 287 nsew signal tristate
rlabel metal3 s 0 13200 800 13320 6 wbs_dat_o[14]
port 288 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 wbs_dat_o[15]
port 289 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 wbs_dat_o[16]
port 290 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 wbs_dat_o[17]
port 291 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 wbs_dat_o[18]
port 292 nsew signal tristate
rlabel metal3 s 0 17824 800 17944 6 wbs_dat_o[19]
port 293 nsew signal tristate
rlabel metal3 s 0 1232 800 1352 6 wbs_dat_o[1]
port 294 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 wbs_dat_o[20]
port 295 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[21]
port 296 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 wbs_dat_o[22]
port 297 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 wbs_dat_o[23]
port 298 nsew signal tristate
rlabel metal3 s 0 22448 800 22568 6 wbs_dat_o[24]
port 299 nsew signal tristate
rlabel metal3 s 0 23400 800 23520 6 wbs_dat_o[25]
port 300 nsew signal tristate
rlabel metal3 s 0 24352 800 24472 6 wbs_dat_o[26]
port 301 nsew signal tristate
rlabel metal3 s 0 25304 800 25424 6 wbs_dat_o[27]
port 302 nsew signal tristate
rlabel metal3 s 0 26120 800 26240 6 wbs_dat_o[28]
port 303 nsew signal tristate
rlabel metal3 s 0 27072 800 27192 6 wbs_dat_o[29]
port 304 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 wbs_dat_o[2]
port 305 nsew signal tristate
rlabel metal3 s 0 28024 800 28144 6 wbs_dat_o[30]
port 306 nsew signal tristate
rlabel metal3 s 0 28976 800 29096 6 wbs_dat_o[31]
port 307 nsew signal tristate
rlabel metal3 s 0 3136 800 3256 6 wbs_dat_o[3]
port 308 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[4]
port 309 nsew signal tristate
rlabel metal3 s 0 4904 800 5024 6 wbs_dat_o[5]
port 310 nsew signal tristate
rlabel metal3 s 0 5856 800 5976 6 wbs_dat_o[6]
port 311 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 wbs_dat_o[7]
port 312 nsew signal tristate
rlabel metal3 s 0 7760 800 7880 6 wbs_dat_o[8]
port 313 nsew signal tristate
rlabel metal3 s 0 8712 800 8832 6 wbs_dat_o[9]
port 314 nsew signal tristate
rlabel metal2 s 5906 59200 5962 60000 6 wbs_sel_i[0]
port 315 nsew signal input
rlabel metal2 s 6642 59200 6698 60000 6 wbs_sel_i[1]
port 316 nsew signal input
rlabel metal2 s 7470 59200 7526 60000 6 wbs_sel_i[2]
port 317 nsew signal input
rlabel metal2 s 8206 59200 8262 60000 6 wbs_sel_i[3]
port 318 nsew signal input
rlabel metal2 s 1950 59200 2006 60000 6 wbs_stb_i
port 319 nsew signal input
rlabel metal2 s 3514 59200 3570 60000 6 wbs_we_i
port 320 nsew signal input
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 321 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 322 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 323 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 324 nsew ground bidirectional
rlabel metal4 s 35588 2176 35908 57664 6 vccd2
port 325 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 57664 6 vccd2
port 326 nsew power bidirectional
rlabel metal4 s 50948 2176 51268 57664 6 vssd2
port 327 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 57664 6 vssd2
port 328 nsew ground bidirectional
rlabel metal4 s 36248 2176 36568 57664 6 vdda1
port 329 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 57664 6 vdda1
port 330 nsew power bidirectional
rlabel metal4 s 51608 2176 51928 57664 6 vssa1
port 331 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 57664 6 vssa1
port 332 nsew ground bidirectional
rlabel metal4 s 36908 2176 37228 57664 6 vdda2
port 333 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 57664 6 vdda2
port 334 nsew power bidirectional
rlabel metal4 s 52268 2176 52588 57664 6 vssa2
port 335 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 57664 6 vssa2
port 336 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
